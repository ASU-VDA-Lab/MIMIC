module fake_ibex_356_n_3238 (n_151, n_85, n_599, n_778, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_738, n_475, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_785, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_772, n_768, n_338, n_173, n_696, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_762, n_410, n_308, n_675, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_744, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_217, n_324, n_391, n_537, n_728, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_232, n_380, n_749, n_281, n_559, n_425, n_3238);

input n_151;
input n_85;
input n_599;
input n_778;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_738;
input n_475;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_785;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_772;
input n_768;
input n_338;
input n_173;
input n_696;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_744;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_3238;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_2720;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_2955;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_850;
wire n_3175;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_1307;
wire n_875;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_1937;
wire n_2311;
wire n_893;
wire n_1654;
wire n_2995;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_787;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_1427;
wire n_852;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_1637;
wire n_841;
wire n_2900;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_2767;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_3023;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_1296;
wire n_3060;
wire n_971;
wire n_1326;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_1702;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3203;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_2256;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3117;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3091;
wire n_3006;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_1217;
wire n_2866;
wire n_3153;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3218;
wire n_2821;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3055;
wire n_1633;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_1236;
wire n_832;
wire n_2297;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_1179;
wire n_907;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_2361;
wire n_1566;
wire n_1464;
wire n_944;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_2954;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2991;
wire n_2234;
wire n_847;
wire n_2699;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_1345;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3072;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1395;
wire n_1115;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2823;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_2418;
wire n_2184;
wire n_1087;
wire n_1400;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2612;
wire n_3034;
wire n_2193;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_2304;
wire n_1746;
wire n_1439;
wire n_2263;
wire n_2352;
wire n_2212;
wire n_2716;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3167;
wire n_997;
wire n_2308;
wire n_2986;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_2903;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2463;
wire n_2654;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_2997;
wire n_1349;
wire n_991;
wire n_1331;
wire n_1223;
wire n_961;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_2862;
wire n_3100;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_2647;
wire n_1626;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3220;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2698;
wire n_2274;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_1673;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2320;
wire n_2268;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_2758;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_826;
wire n_2154;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_839;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_2818;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_975;
wire n_934;
wire n_950;
wire n_2700;
wire n_3139;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_1114;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_2608;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2675;
wire n_2348;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_3085;
wire n_3059;
wire n_2567;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_885;
wire n_1530;
wire n_3215;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2803;
wire n_2816;
wire n_2433;
wire n_1256;
wire n_2798;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3109;
wire n_1961;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2864;
wire n_1632;
wire n_2406;
wire n_3104;
wire n_1542;
wire n_946;
wire n_1547;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_3014;
wire n_1812;
wire n_2703;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_2126;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_3102;
wire n_2872;
wire n_2653;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_2993;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_2843;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_2394;
wire n_3051;
wire n_1572;
wire n_1635;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2929;
wire n_2701;
wire n_3163;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_1986;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_1168;
wire n_865;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_3230;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3223;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3207;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3160;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_2492;
wire n_3081;
wire n_910;
wire n_2291;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2357;
wire n_2618;
wire n_2303;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3114;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_2136;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_3052;
wire n_2443;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_1158;
wire n_1974;
wire n_2988;
wire n_1882;
wire n_2770;
wire n_2961;
wire n_2996;
wire n_2704;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_1736;
wire n_2907;
wire n_1160;
wire n_1442;
wire n_2168;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_1383;
wire n_990;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_3193;
wire n_866;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_1335;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_2040;
wire n_1900;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_3195;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_867;
wire n_983;
wire n_1417;
wire n_2282;
wire n_970;
wire n_2673;
wire n_2430;
wire n_921;
wire n_2676;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

BUFx10_ASAP7_75t_L g787 ( 
.A(n_420),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_761),
.Y(n_788)
);

CKINVDCx14_ASAP7_75t_R g789 ( 
.A(n_354),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_571),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_85),
.Y(n_791)
);

BUFx8_ASAP7_75t_SL g792 ( 
.A(n_742),
.Y(n_792)
);

CKINVDCx14_ASAP7_75t_R g793 ( 
.A(n_268),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_758),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_755),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_422),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_555),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_175),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_313),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_539),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_616),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_760),
.Y(n_802)
);

CKINVDCx14_ASAP7_75t_R g803 ( 
.A(n_743),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_24),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_281),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_168),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_441),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_481),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_587),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_775),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_157),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_489),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_636),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_640),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_753),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_395),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_744),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_669),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_284),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_368),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_332),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_515),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_538),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_621),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_468),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_729),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_702),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_641),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_514),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_733),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_687),
.Y(n_831)
);

CKINVDCx14_ASAP7_75t_R g832 ( 
.A(n_374),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_179),
.Y(n_833)
);

INVx1_ASAP7_75t_SL g834 ( 
.A(n_41),
.Y(n_834)
);

BUFx10_ASAP7_75t_L g835 ( 
.A(n_659),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_408),
.Y(n_836)
);

BUFx10_ASAP7_75t_L g837 ( 
.A(n_541),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_732),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_551),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_782),
.Y(n_840)
);

BUFx2_ASAP7_75t_L g841 ( 
.A(n_783),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_724),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_446),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_754),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_528),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_762),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_632),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_706),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_204),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_784),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_662),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_676),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_431),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_78),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_321),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_395),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_500),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_423),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_690),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_518),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_714),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_688),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_770),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_563),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_477),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_667),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_774),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_130),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_785),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_447),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_187),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_570),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_163),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_296),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_52),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_451),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_734),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_721),
.Y(n_878)
);

BUFx10_ASAP7_75t_L g879 ( 
.A(n_474),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_422),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_452),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_646),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_35),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_498),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_654),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_726),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_427),
.Y(n_887)
);

CKINVDCx14_ASAP7_75t_R g888 ( 
.A(n_124),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_649),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_409),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_106),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_726),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_184),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_138),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_131),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_346),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_403),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_312),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_40),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_705),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_27),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_757),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_587),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_403),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_514),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_375),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_708),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_280),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_21),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_766),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_255),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_681),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_189),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_756),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_748),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_25),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_514),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_232),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_208),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_275),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_642),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_363),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_516),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_769),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_24),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_610),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_457),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_178),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_401),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_752),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_263),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_653),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_744),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_728),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_589),
.Y(n_935)
);

CKINVDCx14_ASAP7_75t_R g936 ( 
.A(n_480),
.Y(n_936)
);

BUFx5_ASAP7_75t_L g937 ( 
.A(n_92),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_581),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_712),
.Y(n_939)
);

INVx1_ASAP7_75t_SL g940 ( 
.A(n_367),
.Y(n_940)
);

BUFx8_ASAP7_75t_SL g941 ( 
.A(n_731),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_235),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_772),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_229),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_429),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_428),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_310),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_780),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_720),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_741),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_631),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_776),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_479),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_596),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_118),
.Y(n_955)
);

CKINVDCx20_ASAP7_75t_R g956 ( 
.A(n_368),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_564),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_311),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_578),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_649),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_764),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_424),
.Y(n_962)
);

CKINVDCx11_ASAP7_75t_R g963 ( 
.A(n_711),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_716),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_528),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_98),
.Y(n_966)
);

CKINVDCx14_ASAP7_75t_R g967 ( 
.A(n_350),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_46),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_504),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_680),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_388),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_781),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_418),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_586),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_681),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_736),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_449),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_170),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_767),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_578),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_268),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_240),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_368),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_730),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_740),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_322),
.Y(n_986)
);

BUFx5_ASAP7_75t_L g987 ( 
.A(n_739),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_164),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_714),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_374),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_338),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_708),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_606),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_299),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_12),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_510),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_310),
.Y(n_997)
);

CKINVDCx16_ASAP7_75t_R g998 ( 
.A(n_91),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_540),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_12),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_508),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_773),
.Y(n_1002)
);

INVx1_ASAP7_75t_SL g1003 ( 
.A(n_123),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_779),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_728),
.Y(n_1005)
);

BUFx5_ASAP7_75t_L g1006 ( 
.A(n_153),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_163),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_149),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_746),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_524),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_696),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_315),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_777),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_612),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_622),
.Y(n_1015)
);

BUFx8_ASAP7_75t_SL g1016 ( 
.A(n_704),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_558),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_710),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_403),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_709),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_655),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_432),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_452),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_22),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_483),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_701),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_439),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_270),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_277),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_313),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_595),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_763),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_759),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_747),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_360),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_321),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_697),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_79),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_348),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_151),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_382),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_499),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_707),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_510),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_672),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_378),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_335),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_737),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_41),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_373),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_107),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_216),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_444),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_417),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_673),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_703),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_298),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_768),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_727),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_548),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_72),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_786),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_718),
.Y(n_1063)
);

CKINVDCx20_ASAP7_75t_R g1064 ( 
.A(n_773),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_723),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_713),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_751),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_628),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_763),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_270),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_55),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_725),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_246),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_600),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_39),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_392),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_86),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_709),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_100),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_771),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_443),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_738),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_388),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_104),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_722),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_717),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_563),
.Y(n_1087)
);

BUFx5_ASAP7_75t_L g1088 ( 
.A(n_460),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_332),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_10),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_391),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_719),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_571),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_259),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_32),
.Y(n_1095)
);

CKINVDCx16_ASAP7_75t_R g1096 ( 
.A(n_82),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_87),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_597),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_227),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_537),
.Y(n_1100)
);

CKINVDCx16_ASAP7_75t_R g1101 ( 
.A(n_59),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_630),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_778),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_645),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_529),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_453),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_42),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_614),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_688),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_715),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_18),
.Y(n_1111)
);

CKINVDCx16_ASAP7_75t_R g1112 ( 
.A(n_430),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_745),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_629),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_75),
.Y(n_1115)
);

BUFx10_ASAP7_75t_L g1116 ( 
.A(n_82),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_105),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_436),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_501),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_750),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_774),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_274),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_402),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_295),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_563),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_630),
.Y(n_1126)
);

INVxp67_ASAP7_75t_L g1127 ( 
.A(n_507),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_613),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_406),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_36),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_460),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_765),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_500),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_427),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_337),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_766),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_51),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_79),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_133),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_267),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_4),
.Y(n_1141)
);

CKINVDCx20_ASAP7_75t_R g1142 ( 
.A(n_257),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_423),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_367),
.Y(n_1144)
);

CKINVDCx20_ASAP7_75t_R g1145 ( 
.A(n_108),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_551),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_354),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_10),
.Y(n_1148)
);

BUFx10_ASAP7_75t_L g1149 ( 
.A(n_621),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_361),
.Y(n_1150)
);

INVx2_ASAP7_75t_SL g1151 ( 
.A(n_748),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_574),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_88),
.Y(n_1153)
);

BUFx10_ASAP7_75t_L g1154 ( 
.A(n_412),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_228),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_283),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_761),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_568),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_365),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_749),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_525),
.Y(n_1161)
);

CKINVDCx20_ASAP7_75t_R g1162 ( 
.A(n_238),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_507),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_353),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_463),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_735),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_684),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_648),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_789),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_789),
.Y(n_1170)
);

CKINVDCx20_ASAP7_75t_R g1171 ( 
.A(n_793),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_832),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_832),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_888),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_812),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1040),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_936),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_973),
.B(n_0),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1105),
.B(n_0),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_987),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_967),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_953),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_803),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_803),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_998),
.B(n_1),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1156),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_953),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_792),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_941),
.Y(n_1189)
);

CKINVDCx14_ASAP7_75t_R g1190 ( 
.A(n_787),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_987),
.Y(n_1191)
);

INVxp67_ASAP7_75t_L g1192 ( 
.A(n_977),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_956),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1016),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_841),
.B(n_2),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1133),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_828),
.B(n_2),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_886),
.B(n_3),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_799),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_963),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1096),
.Y(n_1201)
);

INVxp33_ASAP7_75t_SL g1202 ( 
.A(n_838),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_807),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_956),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1101),
.B(n_3),
.Y(n_1205)
);

INVxp67_ASAP7_75t_SL g1206 ( 
.A(n_805),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_971),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_825),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_1019),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_833),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1112),
.Y(n_1211)
);

INVxp67_ASAP7_75t_SL g1212 ( 
.A(n_805),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_843),
.Y(n_1213)
);

NOR2xp67_ASAP7_75t_L g1214 ( 
.A(n_914),
.B(n_4),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_845),
.Y(n_1215)
);

INVxp67_ASAP7_75t_L g1216 ( 
.A(n_885),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1019),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_857),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_791),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_796),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_797),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_800),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_870),
.Y(n_1223)
);

CKINVDCx14_ASAP7_75t_R g1224 ( 
.A(n_787),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_806),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_872),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_1091),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_1091),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_881),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_808),
.Y(n_1230)
);

INVxp67_ASAP7_75t_SL g1231 ( 
.A(n_966),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_1162),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_804),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_873),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_906),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_988),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_811),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_893),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1151),
.B(n_5),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_921),
.B(n_5),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_904),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_1035),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_989),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_905),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_1036),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_1070),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_816),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_819),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_SL g1249 ( 
.A(n_837),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_1111),
.Y(n_1250)
);

INVxp33_ASAP7_75t_SL g1251 ( 
.A(n_1128),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_922),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_1182),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1190),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1186),
.B(n_1062),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1206),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1212),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1231),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1191),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1224),
.B(n_820),
.Y(n_1260)
);

INVxp67_ASAP7_75t_L g1261 ( 
.A(n_1196),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1192),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1176),
.B(n_821),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1199),
.Y(n_1264)
);

BUFx8_ASAP7_75t_L g1265 ( 
.A(n_1249),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1249),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_1187),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_1193),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1243),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1204),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1203),
.Y(n_1271)
);

XNOR2xp5_ASAP7_75t_L g1272 ( 
.A(n_1169),
.B(n_1129),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1208),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1219),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1210),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1220),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1213),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1221),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1216),
.B(n_794),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1222),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1215),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1218),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1170),
.B(n_844),
.Y(n_1283)
);

NAND2xp33_ASAP7_75t_L g1284 ( 
.A(n_1172),
.B(n_937),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1225),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1223),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1230),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1226),
.A2(n_798),
.B(n_790),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1174),
.B(n_837),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1177),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1181),
.B(n_844),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_1237),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1229),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1247),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1248),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1201),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1238),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1207),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1241),
.B(n_822),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1188),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1244),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_1209),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_SL g1303 ( 
.A1(n_1217),
.A2(n_1145),
.B1(n_1152),
.B2(n_1142),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1171),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1252),
.B(n_823),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_1227),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1183),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1184),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1197),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1197),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1198),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1211),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1198),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1239),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1239),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1189),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1173),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1214),
.Y(n_1318)
);

INVxp67_ASAP7_75t_L g1319 ( 
.A(n_1185),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1178),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1202),
.Y(n_1321)
);

INVxp67_ASAP7_75t_L g1322 ( 
.A(n_1205),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1179),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1179),
.Y(n_1324)
);

OA21x2_ASAP7_75t_L g1325 ( 
.A1(n_1240),
.A2(n_798),
.B(n_790),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1240),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1251),
.B(n_1043),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1195),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1194),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1200),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1228),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1233),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1232),
.Y(n_1333)
);

CKINVDCx20_ASAP7_75t_R g1334 ( 
.A(n_1234),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1235),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1236),
.B(n_1004),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1242),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1245),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1246),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1250),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1219),
.Y(n_1341)
);

INVxp67_ASAP7_75t_L g1342 ( 
.A(n_1196),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1206),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1180),
.Y(n_1344)
);

CKINVDCx16_ASAP7_75t_R g1345 ( 
.A(n_1190),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1206),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1180),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1190),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1190),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1206),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1190),
.B(n_829),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1190),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1180),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1206),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1206),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1190),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1206),
.Y(n_1357)
);

OR2x6_ASAP7_75t_L g1358 ( 
.A(n_1196),
.B(n_1127),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1180),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1206),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1249),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1206),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1192),
.B(n_879),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1190),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1180),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1206),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1190),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1180),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1190),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1190),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1190),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1186),
.B(n_1004),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1190),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1182),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_1182),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1206),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1190),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1190),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1190),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1206),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1190),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1180),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1190),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1192),
.B(n_879),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1186),
.B(n_1065),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1175),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1206),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1180),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1206),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1175),
.B(n_849),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1249),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1206),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1175),
.B(n_853),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1190),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1190),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1288),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1282),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1310),
.B(n_854),
.Y(n_1398)
);

INVx1_ASAP7_75t_SL g1399 ( 
.A(n_1262),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1319),
.B(n_937),
.Y(n_1400)
);

INVx1_ASAP7_75t_SL g1401 ( 
.A(n_1341),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1265),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1322),
.A2(n_1384),
.B1(n_1363),
.B2(n_1342),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1293),
.B(n_937),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1358),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1352),
.B(n_801),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1321),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1261),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1386),
.Y(n_1409)
);

OR2x6_ASAP7_75t_L g1410 ( 
.A(n_1378),
.B(n_801),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1299),
.B(n_937),
.Y(n_1411)
);

INVx5_ASAP7_75t_L g1412 ( 
.A(n_1273),
.Y(n_1412)
);

XOR2xp5_ASAP7_75t_L g1413 ( 
.A(n_1334),
.B(n_1272),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1265),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1288),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1311),
.B(n_1116),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1311),
.B(n_1116),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1280),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1269),
.B(n_1154),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1313),
.B(n_856),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1315),
.B(n_858),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1294),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1281),
.Y(n_1423)
);

AND2x6_ASAP7_75t_L g1424 ( 
.A(n_1266),
.B(n_1017),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1361),
.Y(n_1425)
);

INVx4_ASAP7_75t_SL g1426 ( 
.A(n_1307),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1281),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1324),
.A2(n_1089),
.B1(n_945),
.B2(n_947),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1332),
.Y(n_1429)
);

INVx4_ASAP7_75t_L g1430 ( 
.A(n_1254),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1379),
.Y(n_1431)
);

INVx4_ASAP7_75t_SL g1432 ( 
.A(n_1336),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1337),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1289),
.B(n_1154),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1314),
.B(n_868),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_1253),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1260),
.B(n_1351),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1255),
.A2(n_874),
.B1(n_875),
.B2(n_871),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1259),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1320),
.B(n_876),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1259),
.Y(n_1441)
);

XOR2xp5_ASAP7_75t_L g1442 ( 
.A(n_1267),
.B(n_1034),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_SL g1443 ( 
.A(n_1328),
.B(n_839),
.Y(n_1443)
);

OR2x6_ASAP7_75t_L g1444 ( 
.A(n_1304),
.B(n_1034),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1256),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1305),
.B(n_1006),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1257),
.B(n_1006),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1391),
.B(n_1064),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1258),
.Y(n_1449)
);

BUFx10_ASAP7_75t_L g1450 ( 
.A(n_1348),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1292),
.B(n_835),
.Y(n_1451)
);

AOI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1326),
.A2(n_883),
.B1(n_884),
.B2(n_880),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1295),
.B(n_835),
.Y(n_1453)
);

OAI22xp33_ASAP7_75t_SL g1454 ( 
.A1(n_1274),
.A2(n_890),
.B1(n_894),
.B2(n_887),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1372),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1343),
.A2(n_957),
.B1(n_958),
.B2(n_946),
.Y(n_1456)
);

BUFx8_ASAP7_75t_SL g1457 ( 
.A(n_1268),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1346),
.B(n_895),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1325),
.Y(n_1459)
);

NAND2xp33_ASAP7_75t_L g1460 ( 
.A(n_1349),
.B(n_1006),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1350),
.B(n_897),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1356),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1336),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1364),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1325),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1318),
.B(n_855),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1275),
.Y(n_1467)
);

NAND3xp33_ASAP7_75t_L g1468 ( 
.A(n_1327),
.B(n_899),
.C(n_898),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1354),
.A2(n_962),
.B1(n_965),
.B2(n_959),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1367),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_1395),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1355),
.B(n_1006),
.Y(n_1472)
);

INVx4_ASAP7_75t_L g1473 ( 
.A(n_1369),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1276),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1357),
.B(n_901),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1360),
.Y(n_1476)
);

INVx4_ASAP7_75t_L g1477 ( 
.A(n_1370),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1362),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1296),
.Y(n_1479)
);

INVx1_ASAP7_75t_SL g1480 ( 
.A(n_1278),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1264),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1371),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1366),
.B(n_908),
.Y(n_1483)
);

INVx4_ASAP7_75t_L g1484 ( 
.A(n_1373),
.Y(n_1484)
);

AND3x2_ASAP7_75t_L g1485 ( 
.A(n_1317),
.B(n_1098),
.C(n_842),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1312),
.B(n_834),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1376),
.B(n_911),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1377),
.B(n_1149),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1381),
.Y(n_1489)
);

NAND2xp33_ASAP7_75t_SL g1490 ( 
.A(n_1383),
.B(n_913),
.Y(n_1490)
);

AND2x6_ASAP7_75t_L g1491 ( 
.A(n_1380),
.B(n_860),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1372),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1394),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1290),
.B(n_1098),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1387),
.B(n_916),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1389),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1392),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1283),
.B(n_891),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1291),
.B(n_891),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1291),
.Y(n_1500)
);

BUFx8_ASAP7_75t_SL g1501 ( 
.A(n_1270),
.Y(n_1501)
);

BUFx10_ASAP7_75t_L g1502 ( 
.A(n_1330),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1279),
.A2(n_918),
.B1(n_919),
.B2(n_917),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1271),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1285),
.Y(n_1505)
);

INVx6_ASAP7_75t_L g1506 ( 
.A(n_1385),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_1298),
.Y(n_1507)
);

AND2x6_ASAP7_75t_L g1508 ( 
.A(n_1308),
.B(n_896),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1287),
.B(n_920),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1263),
.B(n_923),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1385),
.B(n_925),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1277),
.B(n_896),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1286),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1300),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1302),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1297),
.B(n_1088),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1301),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1390),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1344),
.Y(n_1519)
);

NAND2xp33_ASAP7_75t_L g1520 ( 
.A(n_1347),
.B(n_1088),
.Y(n_1520)
);

INVx5_ASAP7_75t_L g1521 ( 
.A(n_1353),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1393),
.B(n_927),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1359),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1284),
.B(n_1088),
.Y(n_1524)
);

AND2x6_ASAP7_75t_L g1525 ( 
.A(n_1365),
.B(n_909),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1339),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1316),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1368),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1388),
.B(n_929),
.C(n_928),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1338),
.B(n_931),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1333),
.B(n_942),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_SL g1532 ( 
.A(n_1340),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1382),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1306),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1374),
.Y(n_1535)
);

AO22x2_ASAP7_75t_L g1536 ( 
.A1(n_1331),
.A2(n_1335),
.B1(n_1303),
.B2(n_865),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1340),
.B(n_1329),
.Y(n_1537)
);

OR2x6_ASAP7_75t_L g1538 ( 
.A(n_1340),
.B(n_831),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1375),
.A2(n_1007),
.B1(n_1012),
.B2(n_1008),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1319),
.B(n_944),
.Y(n_1540)
);

INVx5_ASAP7_75t_L g1541 ( 
.A(n_1273),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1288),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1282),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1261),
.B(n_836),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1323),
.A2(n_1025),
.B1(n_1030),
.B2(n_1027),
.Y(n_1545)
);

INVx5_ASAP7_75t_L g1546 ( 
.A(n_1273),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1265),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1310),
.B(n_955),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1282),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1262),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1358),
.Y(n_1551)
);

CKINVDCx6p67_ASAP7_75t_R g1552 ( 
.A(n_1345),
.Y(n_1552)
);

INVxp67_ASAP7_75t_SL g1553 ( 
.A(n_1261),
.Y(n_1553)
);

XNOR2xp5_ASAP7_75t_L g1554 ( 
.A(n_1272),
.B(n_802),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1319),
.B(n_968),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_1334),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1319),
.B(n_969),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1282),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1288),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1282),
.Y(n_1560)
);

INVx6_ASAP7_75t_L g1561 ( 
.A(n_1265),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1310),
.B(n_978),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1265),
.Y(n_1563)
);

INVx4_ASAP7_75t_L g1564 ( 
.A(n_1358),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1386),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1282),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1261),
.B(n_981),
.Y(n_1567)
);

OAI22xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1358),
.A2(n_983),
.B1(n_990),
.B2(n_982),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1310),
.B(n_991),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1319),
.A2(n_995),
.B1(n_996),
.B2(n_994),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1386),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1309),
.B(n_1001),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1282),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1288),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1319),
.B(n_1158),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1310),
.B(n_997),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1319),
.B(n_1163),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1265),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1358),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1310),
.B(n_999),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1319),
.B(n_1164),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1310),
.B(n_1000),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1261),
.B(n_1165),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1309),
.B(n_1049),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1288),
.Y(n_1585)
);

BUFx6f_ASAP7_75t_L g1586 ( 
.A(n_1288),
.Y(n_1586)
);

NOR3xp33_ASAP7_75t_L g1587 ( 
.A(n_1303),
.B(n_980),
.C(n_940),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1540),
.B(n_1010),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1399),
.B(n_847),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1445),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1401),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1449),
.Y(n_1592)
);

NOR2xp67_ASAP7_75t_L g1593 ( 
.A(n_1564),
.B(n_5),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1542),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1408),
.B(n_1553),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1426),
.B(n_813),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1459),
.Y(n_1597)
);

NAND2x1_ASAP7_75t_L g1598 ( 
.A(n_1396),
.B(n_864),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1422),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1465),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1403),
.B(n_1023),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1415),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1555),
.B(n_1024),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1574),
.Y(n_1604)
);

AND2x2_ASAP7_75t_SL g1605 ( 
.A(n_1405),
.B(n_932),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1557),
.B(n_1028),
.Y(n_1606)
);

INVxp67_ASAP7_75t_L g1607 ( 
.A(n_1544),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1476),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1585),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1575),
.B(n_1038),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1414),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1577),
.B(n_1039),
.Y(n_1612)
);

OAI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1539),
.A2(n_1029),
.B1(n_1041),
.B2(n_1022),
.C(n_1003),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1419),
.B(n_1042),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1542),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1478),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1491),
.A2(n_1132),
.B1(n_1104),
.B2(n_1046),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1567),
.B(n_1052),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1581),
.B(n_1044),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1435),
.B(n_1047),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1559),
.Y(n_1621)
);

OAI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1438),
.A2(n_1452),
.B1(n_1570),
.B2(n_1545),
.C(n_1503),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1583),
.B(n_1020),
.Y(n_1623)
);

INVxp33_ASAP7_75t_L g1624 ( 
.A(n_1486),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1496),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1497),
.Y(n_1626)
);

NAND2xp33_ASAP7_75t_L g1627 ( 
.A(n_1424),
.B(n_1075),
.Y(n_1627)
);

OR2x6_ASAP7_75t_L g1628 ( 
.A(n_1561),
.B(n_848),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1551),
.B(n_1072),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1479),
.B(n_1050),
.Y(n_1630)
);

AO22x1_ASAP7_75t_L g1631 ( 
.A1(n_1480),
.A2(n_1053),
.B1(n_1054),
.B2(n_1051),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1409),
.B(n_1073),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1407),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1547),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1586),
.Y(n_1635)
);

AND2x6_ASAP7_75t_SL g1636 ( 
.A(n_1444),
.B(n_1410),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1420),
.B(n_1057),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1421),
.B(n_1060),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1548),
.B(n_1076),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1481),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1491),
.A2(n_1440),
.B1(n_1569),
.B2(n_1562),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1451),
.B(n_1079),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1521),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_R g1644 ( 
.A(n_1402),
.B(n_1078),
.Y(n_1644)
);

INVxp67_ASAP7_75t_SL g1645 ( 
.A(n_1579),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1576),
.B(n_1580),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1504),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1582),
.B(n_1155),
.Y(n_1648)
);

AOI221xp5_ASAP7_75t_L g1649 ( 
.A1(n_1568),
.A2(n_1084),
.B1(n_1087),
.B2(n_1083),
.C(n_1081),
.Y(n_1649)
);

OAI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1410),
.A2(n_1095),
.B1(n_1097),
.B2(n_1093),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1453),
.B(n_1099),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1509),
.B(n_1474),
.Y(n_1652)
);

INVx8_ASAP7_75t_L g1653 ( 
.A(n_1508),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1563),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1400),
.B(n_1115),
.Y(n_1655)
);

OAI22x1_ASAP7_75t_SL g1656 ( 
.A1(n_1556),
.A2(n_1118),
.B1(n_1119),
.B2(n_1117),
.Y(n_1656)
);

AO22x1_ASAP7_75t_L g1657 ( 
.A1(n_1505),
.A2(n_1474),
.B1(n_1433),
.B2(n_1429),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1518),
.B(n_1123),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1513),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_SL g1660 ( 
.A(n_1565),
.B(n_1144),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1571),
.B(n_1124),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1517),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1510),
.B(n_1125),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1458),
.B(n_1131),
.Y(n_1664)
);

BUFx5_ASAP7_75t_L g1665 ( 
.A(n_1427),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1467),
.Y(n_1666)
);

AND2x4_ASAP7_75t_SL g1667 ( 
.A(n_1502),
.B(n_878),
.Y(n_1667)
);

INVx8_ASAP7_75t_L g1668 ( 
.A(n_1508),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1437),
.B(n_1135),
.Y(n_1669)
);

AND2x6_ASAP7_75t_SL g1670 ( 
.A(n_1444),
.B(n_814),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1461),
.B(n_1139),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1457),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1411),
.A2(n_1146),
.B(n_1090),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1475),
.B(n_1483),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1487),
.B(n_1495),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1468),
.A2(n_1143),
.B1(n_1147),
.B2(n_1140),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1522),
.B(n_1148),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1428),
.B(n_1161),
.Y(n_1678)
);

NAND3xp33_ASAP7_75t_SL g1679 ( 
.A(n_1534),
.B(n_900),
.C(n_859),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1397),
.Y(n_1680)
);

INVx4_ASAP7_75t_L g1681 ( 
.A(n_1418),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1431),
.B(n_788),
.Y(n_1682)
);

BUFx3_ASAP7_75t_L g1683 ( 
.A(n_1578),
.Y(n_1683)
);

NOR2xp67_ASAP7_75t_L g1684 ( 
.A(n_1430),
.B(n_6),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_SL g1685 ( 
.A(n_1529),
.B(n_795),
.Y(n_1685)
);

NOR2xp67_ASAP7_75t_L g1686 ( 
.A(n_1473),
.B(n_6),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1456),
.B(n_1150),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1469),
.B(n_1153),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_SL g1689 ( 
.A(n_1543),
.B(n_809),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1511),
.A2(n_815),
.B1(n_826),
.B2(n_824),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1549),
.B(n_827),
.Y(n_1691)
);

NOR3xp33_ASAP7_75t_L g1692 ( 
.A(n_1454),
.B(n_1068),
.C(n_984),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1447),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1442),
.B(n_1535),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1406),
.B(n_1069),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1412),
.Y(n_1696)
);

NOR2x1p5_ASAP7_75t_L g1697 ( 
.A(n_1552),
.B(n_861),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1530),
.A2(n_850),
.B1(n_851),
.B2(n_830),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1463),
.B(n_1086),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1463),
.B(n_862),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1558),
.B(n_1061),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1560),
.B(n_1137),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1472),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1566),
.B(n_1138),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1434),
.B(n_863),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1573),
.B(n_1141),
.Y(n_1706)
);

INVx2_ASAP7_75t_SL g1707 ( 
.A(n_1538),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1443),
.B(n_1077),
.Y(n_1708)
);

AND2x4_ASAP7_75t_SL g1709 ( 
.A(n_1450),
.B(n_878),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1519),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1455),
.B(n_1134),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1531),
.A2(n_869),
.B1(n_877),
.B2(n_867),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1492),
.B(n_1094),
.Y(n_1713)
);

INVx4_ASAP7_75t_L g1714 ( 
.A(n_1426),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1506),
.B(n_892),
.Y(n_1715)
);

INVx8_ASAP7_75t_L g1716 ( 
.A(n_1532),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1500),
.B(n_889),
.Y(n_1717)
);

NAND3xp33_ASAP7_75t_L g1718 ( 
.A(n_1490),
.B(n_903),
.C(n_902),
.Y(n_1718)
);

BUFx6f_ASAP7_75t_L g1719 ( 
.A(n_1412),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1494),
.B(n_1432),
.Y(n_1720)
);

NOR2x1p5_ASAP7_75t_L g1721 ( 
.A(n_1514),
.B(n_907),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1416),
.B(n_1106),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1417),
.B(n_1107),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_SL g1724 ( 
.A(n_1493),
.Y(n_1724)
);

NOR2x2_ASAP7_75t_L g1725 ( 
.A(n_1554),
.B(n_930),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_SL g1726 ( 
.A(n_1412),
.B(n_1541),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1525),
.B(n_1130),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_1541),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1541),
.B(n_939),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1516),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1525),
.B(n_943),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1572),
.A2(n_1584),
.B1(n_1528),
.B2(n_1533),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1498),
.B(n_948),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1499),
.B(n_952),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1523),
.A2(n_938),
.B1(n_986),
.B2(n_864),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1512),
.B(n_961),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_SL g1737 ( 
.A(n_1477),
.B(n_964),
.Y(n_1737)
);

O2A1O1Ixp5_ASAP7_75t_L g1738 ( 
.A1(n_1446),
.A2(n_960),
.B(n_1033),
.C(n_934),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1404),
.A2(n_817),
.B1(n_840),
.B2(n_818),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1423),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1466),
.Y(n_1741)
);

NAND2xp33_ASAP7_75t_L g1742 ( 
.A(n_1524),
.B(n_987),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1488),
.B(n_976),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1526),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1546),
.B(n_979),
.Y(n_1745)
);

INVx2_ASAP7_75t_SL g1746 ( 
.A(n_1537),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1425),
.B(n_992),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1587),
.A2(n_938),
.B1(n_986),
.B2(n_864),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1448),
.B(n_993),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1460),
.B(n_1002),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_SL g1751 ( 
.A(n_1484),
.B(n_1005),
.Y(n_1751)
);

BUFx6f_ASAP7_75t_L g1752 ( 
.A(n_1439),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1527),
.B(n_1470),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1536),
.A2(n_938),
.B1(n_986),
.B2(n_864),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1515),
.B(n_1009),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1441),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1470),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_1501),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1520),
.B(n_1013),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1471),
.B(n_1018),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1471),
.B(n_1021),
.Y(n_1761)
);

NOR3x1_ASAP7_75t_L g1762 ( 
.A(n_1515),
.B(n_852),
.C(n_846),
.Y(n_1762)
);

OR2x6_ASAP7_75t_L g1763 ( 
.A(n_1482),
.B(n_934),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_SL g1764 ( 
.A(n_1462),
.B(n_1026),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1482),
.B(n_866),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1464),
.A2(n_882),
.B1(n_912),
.B2(n_910),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1489),
.B(n_1031),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1489),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1485),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1507),
.Y(n_1770)
);

AND2x6_ASAP7_75t_SL g1771 ( 
.A(n_1413),
.B(n_1436),
.Y(n_1771)
);

OR2x6_ASAP7_75t_L g1772 ( 
.A(n_1561),
.B(n_960),
.Y(n_1772)
);

A2O1A1Ixp33_ASAP7_75t_L g1773 ( 
.A1(n_1398),
.A2(n_915),
.B(n_926),
.C(n_924),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1491),
.A2(n_1100),
.B1(n_1122),
.B2(n_1071),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1540),
.B(n_1032),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1445),
.Y(n_1776)
);

BUFx6f_ASAP7_75t_SL g1777 ( 
.A(n_1414),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1399),
.Y(n_1778)
);

INVx8_ASAP7_75t_L g1779 ( 
.A(n_1508),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1426),
.B(n_933),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1399),
.B(n_1045),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1459),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_SL g1783 ( 
.A(n_1414),
.Y(n_1783)
);

O2A1O1Ixp33_ASAP7_75t_L g1784 ( 
.A1(n_1568),
.A2(n_949),
.B(n_950),
.C(n_935),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1445),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1550),
.B(n_1048),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1445),
.Y(n_1787)
);

AND2x6_ASAP7_75t_SL g1788 ( 
.A(n_1444),
.B(n_951),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1550),
.B(n_1055),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_SL g1790 ( 
.A(n_1564),
.B(n_1056),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1411),
.A2(n_970),
.B(n_954),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1399),
.A2(n_1063),
.B1(n_1066),
.B2(n_1058),
.Y(n_1792)
);

AOI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1399),
.A2(n_1074),
.B1(n_1082),
.B2(n_1067),
.Y(n_1793)
);

CKINVDCx20_ASAP7_75t_R g1794 ( 
.A(n_1457),
.Y(n_1794)
);

INVxp33_ASAP7_75t_L g1795 ( 
.A(n_1408),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1445),
.Y(n_1796)
);

AND2x6_ASAP7_75t_SL g1797 ( 
.A(n_1444),
.B(n_972),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1399),
.A2(n_1113),
.B1(n_1114),
.B2(n_1109),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1550),
.B(n_1120),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1491),
.A2(n_1100),
.B1(n_1122),
.B2(n_1071),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1399),
.B(n_1121),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1399),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1540),
.B(n_1160),
.Y(n_1803)
);

INVx2_ASAP7_75t_SL g1804 ( 
.A(n_1401),
.Y(n_1804)
);

INVx2_ASAP7_75t_SL g1805 ( 
.A(n_1401),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1491),
.A2(n_1159),
.B1(n_1122),
.B2(n_974),
.Y(n_1806)
);

OAI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1641),
.A2(n_1159),
.B1(n_975),
.B2(n_1011),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1607),
.B(n_1167),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1595),
.B(n_1168),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1624),
.B(n_985),
.Y(n_1810)
);

AOI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1646),
.A2(n_1015),
.B(n_1014),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1674),
.A2(n_1675),
.B(n_1742),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1778),
.B(n_1103),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1590),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1802),
.B(n_1126),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1693),
.A2(n_1059),
.B(n_1037),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1592),
.B(n_1136),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1602),
.A2(n_1085),
.B(n_1080),
.Y(n_1818)
);

INVxp67_ASAP7_75t_L g1819 ( 
.A(n_1591),
.Y(n_1819)
);

AOI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1604),
.A2(n_1609),
.B(n_1730),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1795),
.B(n_1092),
.Y(n_1821)
);

OAI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1703),
.A2(n_1102),
.B(n_1092),
.Y(n_1822)
);

NOR2x1_ASAP7_75t_L g1823 ( 
.A(n_1794),
.B(n_1102),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1804),
.B(n_810),
.Y(n_1824)
);

O2A1O1Ixp33_ASAP7_75t_L g1825 ( 
.A1(n_1773),
.A2(n_1166),
.B(n_1157),
.C(n_8),
.Y(n_1825)
);

BUFx6f_ASAP7_75t_L g1826 ( 
.A(n_1594),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1805),
.B(n_810),
.Y(n_1827)
);

A2O1A1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1791),
.A2(n_1110),
.B(n_1108),
.C(n_8),
.Y(n_1828)
);

BUFx3_ASAP7_75t_L g1829 ( 
.A(n_1716),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1623),
.B(n_7),
.Y(n_1830)
);

OAI321xp33_ASAP7_75t_L g1831 ( 
.A1(n_1650),
.A2(n_11),
.A3(n_13),
.B1(n_7),
.B2(n_9),
.C(n_12),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1608),
.B(n_9),
.Y(n_1832)
);

INVxp67_ASAP7_75t_L g1833 ( 
.A(n_1633),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1597),
.Y(n_1834)
);

O2A1O1Ixp33_ASAP7_75t_L g1835 ( 
.A1(n_1613),
.A2(n_1766),
.B(n_1784),
.C(n_1620),
.Y(n_1835)
);

O2A1O1Ixp33_ASAP7_75t_L g1836 ( 
.A1(n_1658),
.A2(n_1637),
.B(n_1639),
.C(n_1638),
.Y(n_1836)
);

OAI21xp33_ASAP7_75t_L g1837 ( 
.A1(n_1614),
.A2(n_11),
.B(n_14),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1616),
.B(n_14),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1625),
.B(n_14),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1589),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1600),
.Y(n_1841)
);

INVx3_ASAP7_75t_L g1842 ( 
.A(n_1719),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1601),
.B(n_15),
.Y(n_1843)
);

BUFx6f_ASAP7_75t_L g1844 ( 
.A(n_1594),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1626),
.B(n_1776),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1655),
.A2(n_16),
.B(n_17),
.Y(n_1846)
);

OAI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1782),
.A2(n_16),
.B(n_17),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1652),
.B(n_18),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1785),
.B(n_19),
.Y(n_1849)
);

OR2x6_ASAP7_75t_L g1850 ( 
.A(n_1653),
.B(n_19),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1787),
.B(n_20),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1796),
.B(n_22),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1629),
.B(n_22),
.Y(n_1853)
);

INVxp67_ASAP7_75t_L g1854 ( 
.A(n_1781),
.Y(n_1854)
);

NAND2xp33_ASAP7_75t_L g1855 ( 
.A(n_1653),
.B(n_24),
.Y(n_1855)
);

OAI21x1_ASAP7_75t_L g1856 ( 
.A1(n_1635),
.A2(n_583),
.B(n_582),
.Y(n_1856)
);

AOI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1588),
.A2(n_23),
.B(n_25),
.Y(n_1857)
);

AOI21xp33_ASAP7_75t_L g1858 ( 
.A1(n_1630),
.A2(n_23),
.B(n_25),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1737),
.B(n_26),
.Y(n_1859)
);

BUFx6f_ASAP7_75t_L g1860 ( 
.A(n_1594),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1603),
.A2(n_28),
.B(n_29),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1606),
.A2(n_28),
.B(n_30),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1640),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1687),
.B(n_30),
.Y(n_1864)
);

OAI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1610),
.A2(n_31),
.B(n_32),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1659),
.Y(n_1866)
);

AO22x1_ASAP7_75t_L g1867 ( 
.A1(n_1672),
.A2(n_33),
.B1(n_34),
.B2(n_32),
.Y(n_1867)
);

NAND2xp33_ASAP7_75t_L g1868 ( 
.A(n_1668),
.B(n_33),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_L g1869 ( 
.A(n_1770),
.B(n_31),
.Y(n_1869)
);

BUFx8_ASAP7_75t_SL g1870 ( 
.A(n_1758),
.Y(n_1870)
);

NOR2xp33_ASAP7_75t_L g1871 ( 
.A(n_1746),
.B(n_34),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1612),
.A2(n_34),
.B(n_35),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1642),
.B(n_36),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_SL g1874 ( 
.A(n_1605),
.B(n_36),
.Y(n_1874)
);

OAI22x1_ASAP7_75t_L g1875 ( 
.A1(n_1697),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1651),
.B(n_37),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1662),
.Y(n_1877)
);

OAI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1619),
.A2(n_37),
.B(n_38),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1647),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1879)
);

OAI21xp33_ASAP7_75t_L g1880 ( 
.A1(n_1648),
.A2(n_40),
.B(n_41),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1666),
.Y(n_1881)
);

AOI21x1_ASAP7_75t_L g1882 ( 
.A1(n_1727),
.A2(n_42),
.B(n_43),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1599),
.Y(n_1883)
);

AOI21xp5_ASAP7_75t_L g1884 ( 
.A1(n_1775),
.A2(n_42),
.B(n_43),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1692),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_SL g1886 ( 
.A(n_1790),
.B(n_1764),
.Y(n_1886)
);

OAI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1664),
.A2(n_46),
.B(n_47),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1688),
.B(n_47),
.Y(n_1888)
);

BUFx6f_ASAP7_75t_L g1889 ( 
.A(n_1615),
.Y(n_1889)
);

A2O1A1Ixp33_ASAP7_75t_L g1890 ( 
.A1(n_1663),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_1890)
);

OR2x6_ASAP7_75t_L g1891 ( 
.A(n_1668),
.B(n_48),
.Y(n_1891)
);

OAI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1677),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_1892)
);

OR2x6_ASAP7_75t_L g1893 ( 
.A(n_1779),
.B(n_51),
.Y(n_1893)
);

OAI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1671),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1894)
);

BUFx6f_ASAP7_75t_L g1895 ( 
.A(n_1615),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1678),
.B(n_56),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1695),
.B(n_57),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1699),
.B(n_58),
.Y(n_1898)
);

A2O1A1Ixp33_ASAP7_75t_L g1899 ( 
.A1(n_1669),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_1899)
);

OAI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1707),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1711),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1700),
.B(n_63),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1645),
.B(n_63),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1801),
.B(n_64),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1713),
.Y(n_1905)
);

AND2x4_ASAP7_75t_L g1906 ( 
.A(n_1714),
.B(n_64),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1803),
.A2(n_65),
.B(n_66),
.Y(n_1907)
);

OAI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1710),
.A2(n_65),
.B(n_66),
.Y(n_1908)
);

NOR3xp33_ASAP7_75t_L g1909 ( 
.A(n_1657),
.B(n_1679),
.C(n_1649),
.Y(n_1909)
);

BUFx3_ASAP7_75t_L g1910 ( 
.A(n_1716),
.Y(n_1910)
);

CKINVDCx8_ASAP7_75t_R g1911 ( 
.A(n_1636),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1644),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1617),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_1913)
);

AOI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1627),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_1914)
);

BUFx2_ASAP7_75t_SL g1915 ( 
.A(n_1777),
.Y(n_1915)
);

NAND3xp33_ASAP7_75t_L g1916 ( 
.A(n_1748),
.B(n_67),
.C(n_70),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1618),
.B(n_71),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1631),
.B(n_1701),
.Y(n_1918)
);

OAI321xp33_ASAP7_75t_L g1919 ( 
.A1(n_1806),
.A2(n_75),
.A3(n_77),
.B1(n_73),
.B2(n_74),
.C(n_76),
.Y(n_1919)
);

AOI21x1_ASAP7_75t_L g1920 ( 
.A1(n_1685),
.A2(n_73),
.B(n_75),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1702),
.B(n_1704),
.Y(n_1921)
);

NAND2xp33_ASAP7_75t_L g1922 ( 
.A(n_1719),
.B(n_78),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1706),
.Y(n_1923)
);

AOI21x1_ASAP7_75t_L g1924 ( 
.A1(n_1684),
.A2(n_1686),
.B(n_1593),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1680),
.Y(n_1925)
);

INVxp67_ASAP7_75t_SL g1926 ( 
.A(n_1719),
.Y(n_1926)
);

AO22x1_ASAP7_75t_L g1927 ( 
.A1(n_1762),
.A2(n_82),
.B1(n_83),
.B2(n_81),
.Y(n_1927)
);

NOR2x1_ASAP7_75t_L g1928 ( 
.A(n_1611),
.B(n_80),
.Y(n_1928)
);

OAI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1732),
.A2(n_84),
.B1(n_80),
.B2(n_81),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_1696),
.Y(n_1930)
);

AOI21x1_ASAP7_75t_L g1931 ( 
.A1(n_1740),
.A2(n_85),
.B(n_86),
.Y(n_1931)
);

BUFx4f_ASAP7_75t_L g1932 ( 
.A(n_1628),
.Y(n_1932)
);

BUFx6f_ASAP7_75t_L g1933 ( 
.A(n_1696),
.Y(n_1933)
);

AOI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1750),
.A2(n_87),
.B(n_88),
.Y(n_1934)
);

NAND2x1p5_ASAP7_75t_L g1935 ( 
.A(n_1714),
.B(n_87),
.Y(n_1935)
);

NAND3xp33_ASAP7_75t_L g1936 ( 
.A(n_1774),
.B(n_88),
.C(n_89),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1759),
.A2(n_89),
.B(n_90),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1722),
.B(n_90),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1723),
.B(n_91),
.Y(n_1939)
);

OAI321xp33_ASAP7_75t_L g1940 ( 
.A1(n_1763),
.A2(n_93),
.A3(n_95),
.B1(n_91),
.B2(n_92),
.C(n_94),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1743),
.A2(n_92),
.B(n_93),
.Y(n_1941)
);

OAI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1708),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_1942)
);

CKINVDCx10_ASAP7_75t_R g1943 ( 
.A(n_1777),
.Y(n_1943)
);

AO21x1_ASAP7_75t_L g1944 ( 
.A1(n_1731),
.A2(n_585),
.B(n_584),
.Y(n_1944)
);

AOI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1765),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_1945)
);

AND2x4_ASAP7_75t_L g1946 ( 
.A(n_1681),
.B(n_101),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1741),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1765),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_1948)
);

INVx3_ASAP7_75t_L g1949 ( 
.A(n_1728),
.Y(n_1949)
);

NAND2x1p5_ASAP7_75t_L g1950 ( 
.A(n_1753),
.B(n_104),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1596),
.Y(n_1951)
);

AOI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1769),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1676),
.B(n_106),
.Y(n_1953)
);

A2O1A1Ixp33_ASAP7_75t_L g1954 ( 
.A1(n_1705),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_1954)
);

OAI21xp5_ASAP7_75t_L g1955 ( 
.A1(n_1736),
.A2(n_109),
.B(n_110),
.Y(n_1955)
);

OAI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1643),
.A2(n_1800),
.B1(n_1772),
.B2(n_1786),
.Y(n_1956)
);

AOI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1689),
.A2(n_111),
.B(n_112),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1596),
.Y(n_1958)
);

AOI21xp5_ASAP7_75t_L g1959 ( 
.A1(n_1691),
.A2(n_111),
.B(n_112),
.Y(n_1959)
);

AOI21x1_ASAP7_75t_L g1960 ( 
.A1(n_1726),
.A2(n_113),
.B(n_114),
.Y(n_1960)
);

OAI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1643),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_1961)
);

O2A1O1Ixp33_ASAP7_75t_L g1962 ( 
.A1(n_1755),
.A2(n_1749),
.B(n_1682),
.C(n_1734),
.Y(n_1962)
);

AOI21x1_ASAP7_75t_L g1963 ( 
.A1(n_1729),
.A2(n_113),
.B(n_114),
.Y(n_1963)
);

OAI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1733),
.A2(n_1712),
.B(n_1698),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1789),
.B(n_115),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1694),
.B(n_115),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1799),
.B(n_116),
.Y(n_1967)
);

INVx3_ASAP7_75t_L g1968 ( 
.A(n_1728),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1792),
.B(n_116),
.Y(n_1969)
);

CKINVDCx20_ASAP7_75t_R g1970 ( 
.A(n_1634),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1690),
.A2(n_117),
.B(n_118),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1780),
.Y(n_1972)
);

OAI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1772),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_1973)
);

AND2x4_ASAP7_75t_L g1974 ( 
.A(n_1768),
.B(n_119),
.Y(n_1974)
);

INVx2_ASAP7_75t_SL g1975 ( 
.A(n_1654),
.Y(n_1975)
);

BUFx6f_ASAP7_75t_L g1976 ( 
.A(n_1752),
.Y(n_1976)
);

OAI21xp33_ASAP7_75t_L g1977 ( 
.A1(n_1793),
.A2(n_119),
.B(n_120),
.Y(n_1977)
);

OAI321xp33_ASAP7_75t_L g1978 ( 
.A1(n_1735),
.A2(n_122),
.A3(n_124),
.B1(n_120),
.B2(n_121),
.C(n_123),
.Y(n_1978)
);

A2O1A1Ixp33_ASAP7_75t_L g1979 ( 
.A1(n_1715),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1665),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1780),
.Y(n_1981)
);

AOI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1632),
.A2(n_122),
.B(n_124),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1720),
.B(n_125),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1798),
.B(n_125),
.Y(n_1984)
);

INVx3_ASAP7_75t_L g1985 ( 
.A(n_1744),
.Y(n_1985)
);

AOI21xp5_ASAP7_75t_L g1986 ( 
.A1(n_1660),
.A2(n_1661),
.B(n_1747),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1717),
.A2(n_126),
.B(n_127),
.Y(n_1987)
);

AOI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1721),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_1988)
);

A2O1A1Ixp33_ASAP7_75t_L g1989 ( 
.A1(n_1718),
.A2(n_130),
.B(n_128),
.C(n_129),
.Y(n_1989)
);

INVx1_ASAP7_75t_SL g1990 ( 
.A(n_1753),
.Y(n_1990)
);

AOI22xp5_ASAP7_75t_L g1991 ( 
.A1(n_1767),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1760),
.B(n_131),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1761),
.B(n_132),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1757),
.B(n_133),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1751),
.B(n_1667),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_SL g1996 ( 
.A(n_1783),
.B(n_132),
.Y(n_1996)
);

AOI21xp5_ASAP7_75t_L g1997 ( 
.A1(n_1752),
.A2(n_134),
.B(n_135),
.Y(n_1997)
);

OAI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1745),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1683),
.B(n_136),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1709),
.B(n_137),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1670),
.B(n_137),
.Y(n_2001)
);

AOI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1756),
.A2(n_139),
.B(n_140),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1756),
.Y(n_2003)
);

OAI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1656),
.A2(n_141),
.B(n_142),
.Y(n_2004)
);

BUFx6f_ASAP7_75t_L g2005 ( 
.A(n_1788),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1724),
.A2(n_141),
.B(n_142),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1724),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1725),
.B(n_142),
.Y(n_2008)
);

AND2x2_ASAP7_75t_SL g2009 ( 
.A(n_1797),
.B(n_143),
.Y(n_2009)
);

OR2x6_ASAP7_75t_L g2010 ( 
.A(n_1783),
.B(n_143),
.Y(n_2010)
);

AOI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_1771),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_2011)
);

OAI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_1738),
.A2(n_144),
.B(n_145),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1607),
.B(n_145),
.Y(n_2013)
);

AOI21x1_ASAP7_75t_L g2014 ( 
.A1(n_1598),
.A2(n_146),
.B(n_147),
.Y(n_2014)
);

OAI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_1738),
.A2(n_146),
.B(n_147),
.Y(n_2015)
);

A2O1A1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_1646),
.A2(n_149),
.B(n_147),
.C(n_148),
.Y(n_2016)
);

NOR2xp67_ASAP7_75t_L g2017 ( 
.A(n_1802),
.B(n_150),
.Y(n_2017)
);

OAI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1641),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1607),
.B(n_152),
.Y(n_2019)
);

AOI21xp33_ASAP7_75t_L g2020 ( 
.A1(n_1624),
.A2(n_154),
.B(n_155),
.Y(n_2020)
);

AND2x4_ASAP7_75t_L g2021 ( 
.A(n_1591),
.B(n_155),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1607),
.B(n_156),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1591),
.B(n_157),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1607),
.B(n_156),
.Y(n_2024)
);

BUFx6f_ASAP7_75t_L g2025 ( 
.A(n_1594),
.Y(n_2025)
);

AND2x4_ASAP7_75t_L g2026 ( 
.A(n_1591),
.B(n_158),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_SL g2027 ( 
.A(n_1591),
.B(n_159),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1597),
.Y(n_2028)
);

AOI21xp33_ASAP7_75t_L g2029 ( 
.A1(n_1624),
.A2(n_160),
.B(n_161),
.Y(n_2029)
);

OR2x4_ASAP7_75t_L g2030 ( 
.A(n_1694),
.B(n_160),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_SL g2031 ( 
.A(n_1802),
.B(n_162),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1597),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1607),
.B(n_165),
.Y(n_2033)
);

NOR2xp67_ASAP7_75t_L g2034 ( 
.A(n_1802),
.B(n_165),
.Y(n_2034)
);

NOR2x1_ASAP7_75t_R g2035 ( 
.A(n_1672),
.B(n_165),
.Y(n_2035)
);

AOI21xp33_ASAP7_75t_L g2036 ( 
.A1(n_1624),
.A2(n_166),
.B(n_167),
.Y(n_2036)
);

INVxp67_ASAP7_75t_SL g2037 ( 
.A(n_1778),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1607),
.B(n_168),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1607),
.B(n_169),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1607),
.B(n_171),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_L g2041 ( 
.A(n_1624),
.B(n_172),
.Y(n_2041)
);

AOI21xp5_ASAP7_75t_L g2042 ( 
.A1(n_1646),
.A2(n_173),
.B(n_174),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1778),
.B(n_173),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1591),
.B(n_177),
.Y(n_2044)
);

OAI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_1641),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_2045)
);

AO21x1_ASAP7_75t_L g2046 ( 
.A1(n_1673),
.A2(n_585),
.B(n_584),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1590),
.Y(n_2047)
);

CKINVDCx10_ASAP7_75t_R g2048 ( 
.A(n_1777),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1778),
.B(n_180),
.Y(n_2049)
);

INVx4_ASAP7_75t_L g2050 ( 
.A(n_1716),
.Y(n_2050)
);

OAI21x1_ASAP7_75t_L g2051 ( 
.A1(n_1621),
.A2(n_588),
.B(n_586),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_L g2052 ( 
.A(n_1624),
.B(n_181),
.Y(n_2052)
);

O2A1O1Ixp33_ASAP7_75t_L g2053 ( 
.A1(n_1646),
.A2(n_184),
.B(n_182),
.C(n_183),
.Y(n_2053)
);

O2A1O1Ixp33_ASAP7_75t_L g2054 ( 
.A1(n_1646),
.A2(n_186),
.B(n_184),
.C(n_185),
.Y(n_2054)
);

INVx11_ASAP7_75t_L g2055 ( 
.A(n_1777),
.Y(n_2055)
);

AO22x1_ASAP7_75t_L g2056 ( 
.A1(n_1672),
.A2(n_190),
.B1(n_191),
.B2(n_189),
.Y(n_2056)
);

BUFx2_ASAP7_75t_L g2057 ( 
.A(n_1778),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_1778),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1591),
.B(n_190),
.Y(n_2059)
);

AOI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_1646),
.A2(n_188),
.B(n_191),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1597),
.Y(n_2061)
);

O2A1O1Ixp5_ASAP7_75t_L g2062 ( 
.A1(n_1598),
.A2(n_194),
.B(n_192),
.C(n_193),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1778),
.B(n_192),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1590),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1607),
.B(n_195),
.Y(n_2065)
);

INVx1_ASAP7_75t_SL g2066 ( 
.A(n_1778),
.Y(n_2066)
);

NAND2xp33_ASAP7_75t_L g2067 ( 
.A(n_1653),
.B(n_197),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1607),
.B(n_196),
.Y(n_2068)
);

CKINVDCx10_ASAP7_75t_R g2069 ( 
.A(n_1777),
.Y(n_2069)
);

NOR3xp33_ASAP7_75t_SL g2070 ( 
.A(n_1672),
.B(n_198),
.C(n_199),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1590),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1590),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1597),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1607),
.B(n_198),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1607),
.B(n_199),
.Y(n_2075)
);

BUFx6f_ASAP7_75t_L g2076 ( 
.A(n_1594),
.Y(n_2076)
);

OA21x2_ASAP7_75t_L g2077 ( 
.A1(n_1738),
.A2(n_200),
.B(n_201),
.Y(n_2077)
);

BUFx6f_ASAP7_75t_L g2078 ( 
.A(n_1594),
.Y(n_2078)
);

INVx3_ASAP7_75t_L g2079 ( 
.A(n_1719),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1590),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_SL g2081 ( 
.A(n_1591),
.B(n_202),
.Y(n_2081)
);

AO21x1_ASAP7_75t_L g2082 ( 
.A1(n_1673),
.A2(n_590),
.B(n_588),
.Y(n_2082)
);

NOR2xp67_ASAP7_75t_L g2083 ( 
.A(n_1802),
.B(n_203),
.Y(n_2083)
);

A2O1A1Ixp33_ASAP7_75t_L g2084 ( 
.A1(n_1646),
.A2(n_205),
.B(n_203),
.C(n_204),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1607),
.B(n_205),
.Y(n_2085)
);

CKINVDCx10_ASAP7_75t_R g2086 ( 
.A(n_1777),
.Y(n_2086)
);

AO32x2_ASAP7_75t_L g2087 ( 
.A1(n_1739),
.A2(n_208),
.A3(n_206),
.B1(n_207),
.B2(n_209),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1778),
.B(n_207),
.Y(n_2088)
);

OAI321xp33_ASAP7_75t_L g2089 ( 
.A1(n_1754),
.A2(n_210),
.A3(n_212),
.B1(n_208),
.B2(n_209),
.C(n_211),
.Y(n_2089)
);

A2O1A1Ixp33_ASAP7_75t_L g2090 ( 
.A1(n_1646),
.A2(n_212),
.B(n_210),
.C(n_211),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_1778),
.Y(n_2091)
);

HB1xp67_ASAP7_75t_L g2092 ( 
.A(n_1778),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1590),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_SL g2094 ( 
.A(n_1591),
.B(n_214),
.Y(n_2094)
);

AO21x1_ASAP7_75t_L g2095 ( 
.A1(n_1673),
.A2(n_592),
.B(n_591),
.Y(n_2095)
);

NOR2xp67_ASAP7_75t_SL g2096 ( 
.A(n_1778),
.B(n_213),
.Y(n_2096)
);

A2O1A1Ixp33_ASAP7_75t_L g2097 ( 
.A1(n_1646),
.A2(n_216),
.B(n_214),
.C(n_215),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1607),
.B(n_215),
.Y(n_2098)
);

AND2x4_ASAP7_75t_L g2099 ( 
.A(n_1591),
.B(n_217),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1607),
.B(n_217),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_1778),
.B(n_218),
.Y(n_2101)
);

INVx1_ASAP7_75t_SL g2102 ( 
.A(n_1778),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1597),
.Y(n_2103)
);

OAI21xp5_ASAP7_75t_L g2104 ( 
.A1(n_1738),
.A2(n_218),
.B(n_219),
.Y(n_2104)
);

NAND3xp33_ASAP7_75t_L g2105 ( 
.A(n_1641),
.B(n_220),
.C(n_221),
.Y(n_2105)
);

NOR2xp67_ASAP7_75t_L g2106 ( 
.A(n_1802),
.B(n_221),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1607),
.B(n_222),
.Y(n_2107)
);

AOI21xp5_ASAP7_75t_L g2108 ( 
.A1(n_1646),
.A2(n_223),
.B(n_224),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1607),
.B(n_224),
.Y(n_2109)
);

AOI21xp5_ASAP7_75t_L g2110 ( 
.A1(n_1646),
.A2(n_225),
.B(n_226),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1607),
.B(n_225),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1597),
.Y(n_2112)
);

OR2x6_ASAP7_75t_L g2113 ( 
.A(n_1653),
.B(n_226),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1590),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_SL g2115 ( 
.A(n_1591),
.B(n_228),
.Y(n_2115)
);

AOI21xp5_ASAP7_75t_L g2116 ( 
.A1(n_1646),
.A2(n_227),
.B(n_229),
.Y(n_2116)
);

AOI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_1646),
.A2(n_230),
.B(n_231),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1607),
.B(n_230),
.Y(n_2118)
);

BUFx6f_ASAP7_75t_L g2119 ( 
.A(n_1594),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1591),
.B(n_234),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1607),
.B(n_233),
.Y(n_2121)
);

BUFx3_ASAP7_75t_L g2122 ( 
.A(n_1716),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1778),
.B(n_234),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_1591),
.B(n_236),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1607),
.B(n_237),
.Y(n_2125)
);

A2O1A1Ixp33_ASAP7_75t_L g2126 ( 
.A1(n_1646),
.A2(n_239),
.B(n_237),
.C(n_238),
.Y(n_2126)
);

BUFx6f_ASAP7_75t_L g2127 ( 
.A(n_1594),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1597),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1590),
.Y(n_2129)
);

BUFx6f_ASAP7_75t_L g2130 ( 
.A(n_1594),
.Y(n_2130)
);

OAI21xp5_ASAP7_75t_L g2131 ( 
.A1(n_1738),
.A2(n_240),
.B(n_241),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1590),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1607),
.B(n_241),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1607),
.B(n_242),
.Y(n_2134)
);

INVx11_ASAP7_75t_L g2135 ( 
.A(n_1777),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1597),
.Y(n_2136)
);

AOI21x1_ASAP7_75t_L g2137 ( 
.A1(n_1598),
.A2(n_242),
.B(n_243),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1607),
.B(n_244),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1590),
.Y(n_2139)
);

NOR3xp33_ASAP7_75t_L g2140 ( 
.A(n_1622),
.B(n_247),
.C(n_246),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1607),
.B(n_245),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1607),
.B(n_248),
.Y(n_2142)
);

AOI21xp5_ASAP7_75t_L g2143 ( 
.A1(n_1646),
.A2(n_249),
.B(n_250),
.Y(n_2143)
);

AOI21xp5_ASAP7_75t_L g2144 ( 
.A1(n_1646),
.A2(n_250),
.B(n_251),
.Y(n_2144)
);

AOI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_1646),
.A2(n_251),
.B(n_252),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1590),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_SL g2147 ( 
.A(n_1591),
.B(n_252),
.Y(n_2147)
);

NOR3xp33_ASAP7_75t_L g2148 ( 
.A(n_1622),
.B(n_254),
.C(n_253),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1607),
.B(n_253),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_1597),
.Y(n_2150)
);

AOI21x1_ASAP7_75t_L g2151 ( 
.A1(n_1598),
.A2(n_253),
.B(n_254),
.Y(n_2151)
);

AOI21x1_ASAP7_75t_L g2152 ( 
.A1(n_1598),
.A2(n_254),
.B(n_255),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1607),
.B(n_255),
.Y(n_2153)
);

OAI21xp5_ASAP7_75t_L g2154 ( 
.A1(n_1738),
.A2(n_256),
.B(n_258),
.Y(n_2154)
);

OAI21xp5_ASAP7_75t_L g2155 ( 
.A1(n_1738),
.A2(n_258),
.B(n_259),
.Y(n_2155)
);

AOI22xp33_ASAP7_75t_L g2156 ( 
.A1(n_1622),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_1778),
.B(n_260),
.Y(n_2157)
);

A2O1A1Ixp33_ASAP7_75t_L g2158 ( 
.A1(n_1646),
.A2(n_262),
.B(n_260),
.C(n_261),
.Y(n_2158)
);

AOI21xp5_ASAP7_75t_L g2159 ( 
.A1(n_1646),
.A2(n_261),
.B(n_262),
.Y(n_2159)
);

AOI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_1622),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.Y(n_2160)
);

A2O1A1Ixp33_ASAP7_75t_L g2161 ( 
.A1(n_1646),
.A2(n_266),
.B(n_264),
.C(n_265),
.Y(n_2161)
);

AOI21xp5_ASAP7_75t_L g2162 ( 
.A1(n_1646),
.A2(n_266),
.B(n_267),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1590),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_1624),
.B(n_269),
.Y(n_2164)
);

AOI21xp5_ASAP7_75t_L g2165 ( 
.A1(n_1646),
.A2(n_271),
.B(n_272),
.Y(n_2165)
);

AOI21xp5_ASAP7_75t_L g2166 ( 
.A1(n_1646),
.A2(n_272),
.B(n_273),
.Y(n_2166)
);

OAI21xp5_ASAP7_75t_L g2167 ( 
.A1(n_1738),
.A2(n_273),
.B(n_274),
.Y(n_2167)
);

INVxp67_ASAP7_75t_L g2168 ( 
.A(n_1778),
.Y(n_2168)
);

INVx1_ASAP7_75t_SL g2169 ( 
.A(n_1778),
.Y(n_2169)
);

BUFx6f_ASAP7_75t_L g2170 ( 
.A(n_1594),
.Y(n_2170)
);

NOR3xp33_ASAP7_75t_L g2171 ( 
.A(n_1622),
.B(n_275),
.C(n_274),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_1607),
.B(n_273),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_1591),
.B(n_278),
.Y(n_2173)
);

AOI21xp5_ASAP7_75t_L g2174 ( 
.A1(n_1646),
.A2(n_276),
.B(n_279),
.Y(n_2174)
);

AOI21xp5_ASAP7_75t_L g2175 ( 
.A1(n_1646),
.A2(n_279),
.B(n_280),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_1607),
.B(n_279),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_SL g2177 ( 
.A(n_1591),
.B(n_282),
.Y(n_2177)
);

INVx3_ASAP7_75t_L g2178 ( 
.A(n_1719),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1590),
.Y(n_2179)
);

INVx5_ASAP7_75t_L g2180 ( 
.A(n_2050),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_1923),
.B(n_280),
.Y(n_2181)
);

BUFx2_ASAP7_75t_L g2182 ( 
.A(n_1970),
.Y(n_2182)
);

OAI21xp5_ASAP7_75t_L g2183 ( 
.A1(n_1836),
.A2(n_283),
.B(n_284),
.Y(n_2183)
);

AOI21xp5_ASAP7_75t_L g2184 ( 
.A1(n_1812),
.A2(n_283),
.B(n_284),
.Y(n_2184)
);

BUFx2_ASAP7_75t_L g2185 ( 
.A(n_1932),
.Y(n_2185)
);

OR2x2_ASAP7_75t_L g2186 ( 
.A(n_2066),
.B(n_2102),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_SL g2187 ( 
.A(n_2050),
.B(n_285),
.Y(n_2187)
);

BUFx6f_ASAP7_75t_L g2188 ( 
.A(n_1826),
.Y(n_2188)
);

OAI21xp5_ASAP7_75t_L g2189 ( 
.A1(n_1921),
.A2(n_285),
.B(n_286),
.Y(n_2189)
);

OR2x2_ASAP7_75t_L g2190 ( 
.A(n_2169),
.B(n_287),
.Y(n_2190)
);

BUFx2_ASAP7_75t_L g2191 ( 
.A(n_2057),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1901),
.B(n_288),
.Y(n_2192)
);

AOI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_1820),
.A2(n_288),
.B(n_289),
.Y(n_2193)
);

AOI21xp33_ASAP7_75t_L g2194 ( 
.A1(n_1835),
.A2(n_289),
.B(n_290),
.Y(n_2194)
);

OAI21x1_ASAP7_75t_L g2195 ( 
.A1(n_1856),
.A2(n_289),
.B(n_290),
.Y(n_2195)
);

OAI21x1_ASAP7_75t_L g2196 ( 
.A1(n_2051),
.A2(n_290),
.B(n_291),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1814),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1834),
.Y(n_2198)
);

OAI21x1_ASAP7_75t_L g2199 ( 
.A1(n_2014),
.A2(n_292),
.B(n_293),
.Y(n_2199)
);

O2A1O1Ixp5_ASAP7_75t_L g2200 ( 
.A1(n_1924),
.A2(n_295),
.B(n_293),
.C(n_294),
.Y(n_2200)
);

INVx2_ASAP7_75t_SL g2201 ( 
.A(n_1829),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1905),
.B(n_294),
.Y(n_2202)
);

AOI21xp5_ASAP7_75t_L g2203 ( 
.A1(n_1986),
.A2(n_294),
.B(n_295),
.Y(n_2203)
);

AOI21xp5_ASAP7_75t_L g2204 ( 
.A1(n_1845),
.A2(n_296),
.B(n_297),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1841),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_1848),
.B(n_297),
.Y(n_2206)
);

AOI21xp5_ASAP7_75t_L g2207 ( 
.A1(n_2012),
.A2(n_297),
.B(n_298),
.Y(n_2207)
);

AOI21xp5_ASAP7_75t_L g2208 ( 
.A1(n_2015),
.A2(n_298),
.B(n_299),
.Y(n_2208)
);

AOI21x1_ASAP7_75t_SL g2209 ( 
.A1(n_1918),
.A2(n_299),
.B(n_300),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2037),
.B(n_300),
.Y(n_2210)
);

AOI21xp5_ASAP7_75t_L g2211 ( 
.A1(n_2104),
.A2(n_300),
.B(n_301),
.Y(n_2211)
);

AOI21x1_ASAP7_75t_L g2212 ( 
.A1(n_1931),
.A2(n_301),
.B(n_302),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2140),
.B(n_301),
.Y(n_2213)
);

INVx3_ASAP7_75t_L g2214 ( 
.A(n_1930),
.Y(n_2214)
);

AO31x2_ASAP7_75t_L g2215 ( 
.A1(n_2046),
.A2(n_304),
.A3(n_302),
.B(n_303),
.Y(n_2215)
);

AO31x2_ASAP7_75t_L g2216 ( 
.A1(n_2082),
.A2(n_305),
.A3(n_303),
.B(n_304),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2028),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_1840),
.B(n_305),
.Y(n_2218)
);

OAI22x1_ASAP7_75t_L g2219 ( 
.A1(n_2011),
.A2(n_307),
.B1(n_305),
.B2(n_306),
.Y(n_2219)
);

OAI21xp33_ASAP7_75t_L g2220 ( 
.A1(n_1874),
.A2(n_306),
.B(n_308),
.Y(n_2220)
);

AO31x2_ASAP7_75t_L g2221 ( 
.A1(n_2095),
.A2(n_311),
.A3(n_308),
.B(n_309),
.Y(n_2221)
);

OAI21xp5_ASAP7_75t_L g2222 ( 
.A1(n_2148),
.A2(n_308),
.B(n_313),
.Y(n_2222)
);

OR2x2_ASAP7_75t_L g2223 ( 
.A(n_2058),
.B(n_314),
.Y(n_2223)
);

AOI21xp5_ASAP7_75t_L g2224 ( 
.A1(n_2131),
.A2(n_314),
.B(n_315),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2171),
.B(n_1843),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2091),
.B(n_316),
.Y(n_2226)
);

BUFx3_ASAP7_75t_L g2227 ( 
.A(n_1910),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2092),
.B(n_316),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2032),
.Y(n_2229)
);

AOI21xp5_ASAP7_75t_L g2230 ( 
.A1(n_2154),
.A2(n_316),
.B(n_317),
.Y(n_2230)
);

AOI21xp5_ASAP7_75t_L g2231 ( 
.A1(n_2155),
.A2(n_318),
.B(n_319),
.Y(n_2231)
);

OAI21x1_ASAP7_75t_L g2232 ( 
.A1(n_2137),
.A2(n_318),
.B(n_319),
.Y(n_2232)
);

AOI21xp5_ASAP7_75t_L g2233 ( 
.A1(n_2167),
.A2(n_318),
.B(n_319),
.Y(n_2233)
);

XNOR2xp5_ASAP7_75t_L g2234 ( 
.A(n_2009),
.B(n_1912),
.Y(n_2234)
);

AOI21xp5_ASAP7_75t_SL g2235 ( 
.A1(n_1850),
.A2(n_320),
.B(n_322),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2047),
.B(n_2064),
.Y(n_2236)
);

NOR2xp67_ASAP7_75t_SL g2237 ( 
.A(n_1911),
.B(n_323),
.Y(n_2237)
);

BUFx8_ASAP7_75t_L g2238 ( 
.A(n_2122),
.Y(n_2238)
);

AOI221xp5_ASAP7_75t_L g2239 ( 
.A1(n_1830),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.C(n_326),
.Y(n_2239)
);

AOI21xp5_ASAP7_75t_L g2240 ( 
.A1(n_2170),
.A2(n_1844),
.B(n_1826),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2071),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2072),
.B(n_326),
.Y(n_2242)
);

OAI21xp5_ASAP7_75t_L g2243 ( 
.A1(n_1873),
.A2(n_327),
.B(n_328),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2061),
.Y(n_2244)
);

INVxp67_ASAP7_75t_L g2245 ( 
.A(n_2031),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_1854),
.B(n_329),
.Y(n_2246)
);

OAI21x1_ASAP7_75t_L g2247 ( 
.A1(n_2151),
.A2(n_329),
.B(n_330),
.Y(n_2247)
);

OAI21x1_ASAP7_75t_L g2248 ( 
.A1(n_2152),
.A2(n_330),
.B(n_331),
.Y(n_2248)
);

A2O1A1Ixp33_ASAP7_75t_L g2249 ( 
.A1(n_2160),
.A2(n_1876),
.B(n_1967),
.C(n_1825),
.Y(n_2249)
);

OAI22xp5_ASAP7_75t_L g2250 ( 
.A1(n_2160),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_2250)
);

BUFx6f_ASAP7_75t_L g2251 ( 
.A(n_1860),
.Y(n_2251)
);

OAI21x1_ASAP7_75t_L g2252 ( 
.A1(n_2003),
.A2(n_333),
.B(n_334),
.Y(n_2252)
);

AO21x1_ASAP7_75t_L g2253 ( 
.A1(n_1908),
.A2(n_594),
.B(n_593),
.Y(n_2253)
);

INVx4_ASAP7_75t_L g2254 ( 
.A(n_2055),
.Y(n_2254)
);

AO31x2_ASAP7_75t_L g2255 ( 
.A1(n_1944),
.A2(n_337),
.A3(n_335),
.B(n_336),
.Y(n_2255)
);

BUFx6f_ASAP7_75t_L g2256 ( 
.A(n_1889),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2073),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2080),
.Y(n_2258)
);

AO31x2_ASAP7_75t_L g2259 ( 
.A1(n_1828),
.A2(n_341),
.A3(n_339),
.B(n_340),
.Y(n_2259)
);

OAI21xp5_ASAP7_75t_L g2260 ( 
.A1(n_1811),
.A2(n_341),
.B(n_342),
.Y(n_2260)
);

AOI21x1_ASAP7_75t_L g2261 ( 
.A1(n_1882),
.A2(n_341),
.B(n_342),
.Y(n_2261)
);

AO31x2_ASAP7_75t_L g2262 ( 
.A1(n_1807),
.A2(n_345),
.A3(n_343),
.B(n_344),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2093),
.B(n_344),
.Y(n_2263)
);

OR2x2_ASAP7_75t_L g2264 ( 
.A(n_2168),
.B(n_344),
.Y(n_2264)
);

AOI21x1_ASAP7_75t_SL g2265 ( 
.A1(n_1965),
.A2(n_345),
.B(n_346),
.Y(n_2265)
);

AOI22xp5_ASAP7_75t_L g2266 ( 
.A1(n_1853),
.A2(n_347),
.B1(n_345),
.B2(n_346),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2114),
.Y(n_2267)
);

O2A1O1Ixp5_ASAP7_75t_L g2268 ( 
.A1(n_1824),
.A2(n_349),
.B(n_347),
.C(n_348),
.Y(n_2268)
);

INVx2_ASAP7_75t_SL g2269 ( 
.A(n_1943),
.Y(n_2269)
);

INVxp67_ASAP7_75t_SL g2270 ( 
.A(n_1833),
.Y(n_2270)
);

CKINVDCx8_ASAP7_75t_R g2271 ( 
.A(n_1943),
.Y(n_2271)
);

INVx1_ASAP7_75t_SL g2272 ( 
.A(n_1990),
.Y(n_2272)
);

OAI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_1816),
.A2(n_349),
.B(n_350),
.Y(n_2273)
);

O2A1O1Ixp5_ASAP7_75t_L g2274 ( 
.A1(n_1827),
.A2(n_352),
.B(n_350),
.C(n_351),
.Y(n_2274)
);

AO221x1_ASAP7_75t_L g2275 ( 
.A1(n_1875),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.C(n_355),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2129),
.B(n_353),
.Y(n_2276)
);

BUFx10_ASAP7_75t_L g2277 ( 
.A(n_2010),
.Y(n_2277)
);

OAI22x1_ASAP7_75t_L g2278 ( 
.A1(n_2011),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2043),
.B(n_357),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2049),
.B(n_357),
.Y(n_2280)
);

BUFx6f_ASAP7_75t_L g2281 ( 
.A(n_1895),
.Y(n_2281)
);

NAND3xp33_ASAP7_75t_L g2282 ( 
.A(n_1909),
.B(n_358),
.C(n_359),
.Y(n_2282)
);

HB1xp67_ASAP7_75t_L g2283 ( 
.A(n_1850),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2132),
.Y(n_2284)
);

AND2x4_ASAP7_75t_L g2285 ( 
.A(n_1891),
.B(n_358),
.Y(n_2285)
);

BUFx2_ASAP7_75t_L g2286 ( 
.A(n_1891),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2139),
.Y(n_2287)
);

AND2x4_ASAP7_75t_L g2288 ( 
.A(n_1891),
.B(n_360),
.Y(n_2288)
);

OA22x2_ASAP7_75t_L g2289 ( 
.A1(n_1893),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_2289)
);

INVx3_ASAP7_75t_L g2290 ( 
.A(n_1930),
.Y(n_2290)
);

AOI21xp5_ASAP7_75t_L g2291 ( 
.A1(n_1895),
.A2(n_2076),
.B(n_2025),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2103),
.Y(n_2292)
);

AOI21xp5_ASAP7_75t_L g2293 ( 
.A1(n_2025),
.A2(n_2078),
.B(n_2076),
.Y(n_2293)
);

A2O1A1Ixp33_ASAP7_75t_L g2294 ( 
.A1(n_1865),
.A2(n_364),
.B(n_362),
.C(n_363),
.Y(n_2294)
);

NAND2x1p5_ASAP7_75t_L g2295 ( 
.A(n_1886),
.B(n_363),
.Y(n_2295)
);

OAI21x1_ASAP7_75t_L g2296 ( 
.A1(n_1980),
.A2(n_366),
.B(n_367),
.Y(n_2296)
);

AO31x2_ASAP7_75t_L g2297 ( 
.A1(n_2018),
.A2(n_371),
.A3(n_369),
.B(n_370),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2146),
.B(n_369),
.Y(n_2298)
);

AOI21xp5_ASAP7_75t_SL g2299 ( 
.A1(n_1893),
.A2(n_369),
.B(n_370),
.Y(n_2299)
);

OAI21x1_ASAP7_75t_SL g2300 ( 
.A1(n_1847),
.A2(n_370),
.B(n_371),
.Y(n_2300)
);

A2O1A1Ixp33_ASAP7_75t_L g2301 ( 
.A1(n_1872),
.A2(n_374),
.B(n_372),
.C(n_373),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2163),
.B(n_372),
.Y(n_2302)
);

OAI21xp5_ASAP7_75t_L g2303 ( 
.A1(n_1822),
.A2(n_375),
.B(n_376),
.Y(n_2303)
);

BUFx2_ASAP7_75t_L g2304 ( 
.A(n_1893),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2179),
.Y(n_2305)
);

OAI21x1_ASAP7_75t_L g2306 ( 
.A1(n_1960),
.A2(n_377),
.B(n_378),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_1898),
.B(n_378),
.Y(n_2307)
);

INVx1_ASAP7_75t_SL g2308 ( 
.A(n_1883),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_1866),
.Y(n_2309)
);

OAI21xp5_ASAP7_75t_L g2310 ( 
.A1(n_2105),
.A2(n_379),
.B(n_380),
.Y(n_2310)
);

OAI21xp33_ASAP7_75t_L g2311 ( 
.A1(n_1837),
.A2(n_379),
.B(n_380),
.Y(n_2311)
);

INVxp67_ASAP7_75t_L g2312 ( 
.A(n_1996),
.Y(n_2312)
);

NAND2x1p5_ASAP7_75t_L g2313 ( 
.A(n_2096),
.B(n_1975),
.Y(n_2313)
);

AND3x4_ASAP7_75t_L g2314 ( 
.A(n_2070),
.B(n_381),
.C(n_383),
.Y(n_2314)
);

AOI21xp5_ASAP7_75t_L g2315 ( 
.A1(n_2119),
.A2(n_2130),
.B(n_2127),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1877),
.Y(n_2316)
);

CKINVDCx5p33_ASAP7_75t_R g2317 ( 
.A(n_2048),
.Y(n_2317)
);

OAI21x1_ASAP7_75t_L g2318 ( 
.A1(n_2112),
.A2(n_383),
.B(n_384),
.Y(n_2318)
);

OAI21xp5_ASAP7_75t_L g2319 ( 
.A1(n_1818),
.A2(n_384),
.B(n_385),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_1902),
.B(n_386),
.Y(n_2320)
);

AO31x2_ASAP7_75t_L g2321 ( 
.A1(n_2045),
.A2(n_389),
.A3(n_387),
.B(n_388),
.Y(n_2321)
);

OAI21xp5_ASAP7_75t_L g2322 ( 
.A1(n_2156),
.A2(n_387),
.B(n_389),
.Y(n_2322)
);

INVx5_ASAP7_75t_L g2323 ( 
.A(n_2113),
.Y(n_2323)
);

A2O1A1Ixp33_ASAP7_75t_L g2324 ( 
.A1(n_1878),
.A2(n_392),
.B(n_390),
.C(n_391),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2128),
.Y(n_2325)
);

OAI21x1_ASAP7_75t_L g2326 ( 
.A1(n_2136),
.A2(n_390),
.B(n_392),
.Y(n_2326)
);

AOI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_2130),
.A2(n_393),
.B(n_394),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_1832),
.Y(n_2328)
);

AND2x4_ASAP7_75t_L g2329 ( 
.A(n_2113),
.B(n_393),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_1809),
.B(n_394),
.Y(n_2330)
);

AND2x4_ASAP7_75t_L g2331 ( 
.A(n_2113),
.B(n_396),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2063),
.B(n_397),
.Y(n_2332)
);

OAI21x1_ASAP7_75t_L g2333 ( 
.A1(n_2150),
.A2(n_398),
.B(n_399),
.Y(n_2333)
);

OAI21x1_ASAP7_75t_L g2334 ( 
.A1(n_1920),
.A2(n_400),
.B(n_402),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2088),
.B(n_404),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1838),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_1925),
.Y(n_2337)
);

A2O1A1Ixp33_ASAP7_75t_L g2338 ( 
.A1(n_1971),
.A2(n_407),
.B(n_405),
.C(n_406),
.Y(n_2338)
);

BUFx10_ASAP7_75t_L g2339 ( 
.A(n_1999),
.Y(n_2339)
);

OAI21x1_ASAP7_75t_L g2340 ( 
.A1(n_1963),
.A2(n_405),
.B(n_406),
.Y(n_2340)
);

HB1xp67_ASAP7_75t_L g2341 ( 
.A(n_1819),
.Y(n_2341)
);

AOI21xp33_ASAP7_75t_L g2342 ( 
.A1(n_1962),
.A2(n_409),
.B(n_410),
.Y(n_2342)
);

OAI21x1_ASAP7_75t_L g2343 ( 
.A1(n_2077),
.A2(n_409),
.B(n_410),
.Y(n_2343)
);

A2O1A1Ixp33_ASAP7_75t_L g2344 ( 
.A1(n_1887),
.A2(n_412),
.B(n_410),
.C(n_411),
.Y(n_2344)
);

OAI21xp5_ASAP7_75t_L g2345 ( 
.A1(n_1964),
.A2(n_411),
.B(n_413),
.Y(n_2345)
);

INVx3_ASAP7_75t_L g2346 ( 
.A(n_1933),
.Y(n_2346)
);

OAI21xp5_ASAP7_75t_L g2347 ( 
.A1(n_1992),
.A2(n_1993),
.B(n_1888),
.Y(n_2347)
);

OAI21x1_ASAP7_75t_L g2348 ( 
.A1(n_2062),
.A2(n_413),
.B(n_414),
.Y(n_2348)
);

BUFx3_ASAP7_75t_L g2349 ( 
.A(n_1870),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_1839),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_1897),
.B(n_415),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2101),
.B(n_415),
.Y(n_2352)
);

NAND2x1p5_ASAP7_75t_L g2353 ( 
.A(n_1946),
.B(n_416),
.Y(n_2353)
);

OAI21xp5_ASAP7_75t_L g2354 ( 
.A1(n_1864),
.A2(n_417),
.B(n_418),
.Y(n_2354)
);

AOI21xp5_ASAP7_75t_L g2355 ( 
.A1(n_1896),
.A2(n_418),
.B(n_419),
.Y(n_2355)
);

BUFx3_ASAP7_75t_L g2356 ( 
.A(n_1999),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_1849),
.Y(n_2357)
);

INVx4_ASAP7_75t_L g2358 ( 
.A(n_2135),
.Y(n_2358)
);

INVx1_ASAP7_75t_SL g2359 ( 
.A(n_1946),
.Y(n_2359)
);

AOI21x1_ASAP7_75t_L g2360 ( 
.A1(n_1851),
.A2(n_421),
.B(n_422),
.Y(n_2360)
);

BUFx12f_ASAP7_75t_L g2361 ( 
.A(n_2005),
.Y(n_2361)
);

INVx3_ASAP7_75t_L g2362 ( 
.A(n_1933),
.Y(n_2362)
);

NAND2x1p5_ASAP7_75t_L g2363 ( 
.A(n_1906),
.B(n_424),
.Y(n_2363)
);

BUFx6f_ASAP7_75t_L g2364 ( 
.A(n_1976),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2013),
.B(n_425),
.Y(n_2365)
);

OAI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_1938),
.A2(n_426),
.B(n_427),
.Y(n_2366)
);

OAI21xp5_ASAP7_75t_L g2367 ( 
.A1(n_1939),
.A2(n_426),
.B(n_428),
.Y(n_2367)
);

OAI22xp5_ASAP7_75t_L g2368 ( 
.A1(n_1914),
.A2(n_429),
.B1(n_426),
.B2(n_428),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_1863),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2019),
.B(n_429),
.Y(n_2370)
);

AND2x4_ASAP7_75t_L g2371 ( 
.A(n_1949),
.B(n_430),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2022),
.B(n_430),
.Y(n_2372)
);

AOI221x1_ASAP7_75t_L g2373 ( 
.A1(n_1880),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.C(n_434),
.Y(n_2373)
);

AOI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_1966),
.A2(n_435),
.B1(n_433),
.B2(n_434),
.Y(n_2374)
);

OAI21x1_ASAP7_75t_L g2375 ( 
.A1(n_1842),
.A2(n_433),
.B(n_434),
.Y(n_2375)
);

INVxp67_ASAP7_75t_SL g2376 ( 
.A(n_1855),
.Y(n_2376)
);

BUFx10_ASAP7_75t_L g2377 ( 
.A(n_1906),
.Y(n_2377)
);

INVx6_ASAP7_75t_SL g2378 ( 
.A(n_2021),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2024),
.B(n_436),
.Y(n_2379)
);

OAI22x1_ASAP7_75t_L g2380 ( 
.A1(n_1988),
.A2(n_439),
.B1(n_437),
.B2(n_438),
.Y(n_2380)
);

NOR2x1_ASAP7_75t_L g2381 ( 
.A(n_1915),
.B(n_437),
.Y(n_2381)
);

CKINVDCx5p33_ASAP7_75t_R g2382 ( 
.A(n_2048),
.Y(n_2382)
);

NOR2xp33_ASAP7_75t_L g2383 ( 
.A(n_1951),
.B(n_437),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_1852),
.Y(n_2384)
);

OAI21x1_ASAP7_75t_L g2385 ( 
.A1(n_2079),
.A2(n_440),
.B(n_441),
.Y(n_2385)
);

CKINVDCx5p33_ASAP7_75t_R g2386 ( 
.A(n_2069),
.Y(n_2386)
);

OAI22xp5_ASAP7_75t_L g2387 ( 
.A1(n_1914),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.Y(n_2387)
);

OR2x2_ASAP7_75t_L g2388 ( 
.A(n_1904),
.B(n_442),
.Y(n_2388)
);

A2O1A1Ixp33_ASAP7_75t_L g2389 ( 
.A1(n_1857),
.A2(n_447),
.B(n_445),
.C(n_446),
.Y(n_2389)
);

A2O1A1Ixp33_ASAP7_75t_L g2390 ( 
.A1(n_1861),
.A2(n_448),
.B(n_445),
.C(n_447),
.Y(n_2390)
);

OAI22xp33_ASAP7_75t_L g2391 ( 
.A1(n_1945),
.A2(n_452),
.B1(n_450),
.B2(n_451),
.Y(n_2391)
);

AOI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_1956),
.A2(n_451),
.B(n_453),
.Y(n_2392)
);

BUFx2_ASAP7_75t_L g2393 ( 
.A(n_1926),
.Y(n_2393)
);

AO21x2_ASAP7_75t_L g2394 ( 
.A1(n_1955),
.A2(n_454),
.B(n_455),
.Y(n_2394)
);

AND2x4_ASAP7_75t_L g2395 ( 
.A(n_1949),
.B(n_455),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_1958),
.B(n_1972),
.Y(n_2396)
);

NOR2xp67_ASAP7_75t_L g2397 ( 
.A(n_2007),
.B(n_456),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2123),
.B(n_458),
.Y(n_2398)
);

CKINVDCx14_ASAP7_75t_R g2399 ( 
.A(n_2005),
.Y(n_2399)
);

OAI21x1_ASAP7_75t_L g2400 ( 
.A1(n_2178),
.A2(n_459),
.B(n_461),
.Y(n_2400)
);

INVx1_ASAP7_75t_SL g2401 ( 
.A(n_2157),
.Y(n_2401)
);

INVx4_ASAP7_75t_L g2402 ( 
.A(n_2178),
.Y(n_2402)
);

AOI21xp5_ASAP7_75t_L g2403 ( 
.A1(n_1881),
.A2(n_461),
.B(n_462),
.Y(n_2403)
);

OAI21x1_ASAP7_75t_L g2404 ( 
.A1(n_1997),
.A2(n_462),
.B(n_463),
.Y(n_2404)
);

NOR2xp67_ASAP7_75t_L g2405 ( 
.A(n_1995),
.B(n_462),
.Y(n_2405)
);

BUFx6f_ASAP7_75t_L g2406 ( 
.A(n_1976),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_SL g2407 ( 
.A(n_2017),
.B(n_2034),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2033),
.B(n_463),
.Y(n_2408)
);

OAI22xp5_ASAP7_75t_L g2409 ( 
.A1(n_1945),
.A2(n_466),
.B1(n_464),
.B2(n_465),
.Y(n_2409)
);

OAI21xp33_ASAP7_75t_L g2410 ( 
.A1(n_1977),
.A2(n_464),
.B(n_465),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2038),
.B(n_464),
.Y(n_2411)
);

AO31x2_ASAP7_75t_L g2412 ( 
.A1(n_2016),
.A2(n_467),
.A3(n_465),
.B(n_466),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2039),
.B(n_467),
.Y(n_2413)
);

OAI22xp5_ASAP7_75t_L g2414 ( 
.A1(n_1948),
.A2(n_1991),
.B1(n_1885),
.B2(n_1950),
.Y(n_2414)
);

AND2x6_ASAP7_75t_L g2415 ( 
.A(n_1974),
.B(n_468),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2040),
.B(n_468),
.Y(n_2416)
);

A2O1A1Ixp33_ASAP7_75t_L g2417 ( 
.A1(n_1862),
.A2(n_471),
.B(n_469),
.C(n_470),
.Y(n_2417)
);

CKINVDCx5p33_ASAP7_75t_R g2418 ( 
.A(n_2086),
.Y(n_2418)
);

AOI21x1_ASAP7_75t_L g2419 ( 
.A1(n_2083),
.A2(n_471),
.B(n_472),
.Y(n_2419)
);

OAI21xp33_ASAP7_75t_SL g2420 ( 
.A1(n_1948),
.A2(n_472),
.B(n_473),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_SL g2421 ( 
.A(n_2106),
.B(n_597),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2065),
.B(n_474),
.Y(n_2422)
);

OAI21x1_ASAP7_75t_L g2423 ( 
.A1(n_2002),
.A2(n_475),
.B(n_476),
.Y(n_2423)
);

NAND3xp33_ASAP7_75t_L g2424 ( 
.A(n_2053),
.B(n_475),
.C(n_476),
.Y(n_2424)
);

NOR2xp33_ASAP7_75t_L g2425 ( 
.A(n_1981),
.B(n_476),
.Y(n_2425)
);

OAI21x1_ASAP7_75t_L g2426 ( 
.A1(n_1985),
.A2(n_477),
.B(n_478),
.Y(n_2426)
);

OR2x2_ASAP7_75t_L g2427 ( 
.A(n_2068),
.B(n_477),
.Y(n_2427)
);

HB1xp67_ASAP7_75t_L g2428 ( 
.A(n_2026),
.Y(n_2428)
);

AO21x1_ASAP7_75t_L g2429 ( 
.A1(n_1868),
.A2(n_599),
.B(n_598),
.Y(n_2429)
);

OR2x2_ASAP7_75t_L g2430 ( 
.A(n_2074),
.B(n_479),
.Y(n_2430)
);

OA22x2_ASAP7_75t_L g2431 ( 
.A1(n_2004),
.A2(n_1991),
.B1(n_1952),
.B2(n_2026),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2075),
.B(n_480),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2085),
.B(n_481),
.Y(n_2433)
);

A2O1A1Ixp33_ASAP7_75t_L g2434 ( 
.A1(n_1846),
.A2(n_484),
.B(n_482),
.C(n_483),
.Y(n_2434)
);

AOI21xp5_ASAP7_75t_L g2435 ( 
.A1(n_1817),
.A2(n_482),
.B(n_483),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2098),
.B(n_484),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2100),
.B(n_485),
.Y(n_2437)
);

AND2x4_ASAP7_75t_L g2438 ( 
.A(n_1968),
.B(n_486),
.Y(n_2438)
);

AND2x2_ASAP7_75t_L g2439 ( 
.A(n_2008),
.B(n_486),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2107),
.B(n_487),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2109),
.B(n_487),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2111),
.B(n_488),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2118),
.B(n_488),
.Y(n_2443)
);

OAI21xp5_ASAP7_75t_SL g2444 ( 
.A1(n_1935),
.A2(n_490),
.B(n_491),
.Y(n_2444)
);

NOR2xp33_ASAP7_75t_R g2445 ( 
.A(n_2067),
.B(n_490),
.Y(n_2445)
);

BUFx3_ASAP7_75t_L g2446 ( 
.A(n_2099),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_1947),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_1969),
.B(n_492),
.Y(n_2448)
);

BUFx6f_ASAP7_75t_L g2449 ( 
.A(n_1976),
.Y(n_2449)
);

AOI221xp5_ASAP7_75t_SL g2450 ( 
.A1(n_1884),
.A2(n_494),
.B1(n_492),
.B2(n_493),
.C(n_495),
.Y(n_2450)
);

INVx4_ASAP7_75t_L g2451 ( 
.A(n_1974),
.Y(n_2451)
);

AOI21xp5_ASAP7_75t_L g2452 ( 
.A1(n_1922),
.A2(n_494),
.B(n_495),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2087),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2087),
.Y(n_2454)
);

AOI21xp33_ASAP7_75t_L g2455 ( 
.A1(n_2121),
.A2(n_496),
.B(n_497),
.Y(n_2455)
);

CKINVDCx20_ASAP7_75t_R g2456 ( 
.A(n_2030),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_1871),
.B(n_497),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2125),
.B(n_498),
.Y(n_2458)
);

INVx2_ASAP7_75t_SL g2459 ( 
.A(n_1928),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2087),
.Y(n_2460)
);

OAI22xp5_ASAP7_75t_L g2461 ( 
.A1(n_1952),
.A2(n_503),
.B1(n_501),
.B2(n_502),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2133),
.B(n_503),
.Y(n_2462)
);

AOI21xp33_ASAP7_75t_L g2463 ( 
.A1(n_2134),
.A2(n_2141),
.B(n_2138),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_1942),
.Y(n_2464)
);

OAI21xp5_ASAP7_75t_L g2465 ( 
.A1(n_1907),
.A2(n_1953),
.B(n_1941),
.Y(n_2465)
);

INVx1_ASAP7_75t_SL g2466 ( 
.A(n_2000),
.Y(n_2466)
);

NAND2x1_ASAP7_75t_L g2467 ( 
.A(n_1940),
.B(n_505),
.Y(n_2467)
);

AOI22xp5_ASAP7_75t_L g2468 ( 
.A1(n_1983),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.Y(n_2468)
);

AOI21xp33_ASAP7_75t_L g2469 ( 
.A1(n_2142),
.A2(n_506),
.B(n_508),
.Y(n_2469)
);

NAND2x1p5_ASAP7_75t_L g2470 ( 
.A(n_1823),
.B(n_509),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2149),
.B(n_511),
.Y(n_2471)
);

AOI21xp33_ASAP7_75t_L g2472 ( 
.A1(n_2153),
.A2(n_511),
.B(n_512),
.Y(n_2472)
);

A2O1A1Ixp33_ASAP7_75t_L g2473 ( 
.A1(n_2054),
.A2(n_516),
.B(n_513),
.C(n_515),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2172),
.B(n_2176),
.Y(n_2474)
);

OAI21xp33_ASAP7_75t_L g2475 ( 
.A1(n_1810),
.A2(n_517),
.B(n_518),
.Y(n_2475)
);

INVx4_ASAP7_75t_L g2476 ( 
.A(n_2035),
.Y(n_2476)
);

OAI21xp5_ASAP7_75t_L g2477 ( 
.A1(n_1916),
.A2(n_519),
.B(n_520),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_1903),
.B(n_520),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_1808),
.B(n_521),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_2001),
.Y(n_2480)
);

OA21x2_ASAP7_75t_L g2481 ( 
.A1(n_2042),
.A2(n_522),
.B(n_523),
.Y(n_2481)
);

NAND2x1p5_ASAP7_75t_L g2482 ( 
.A(n_1859),
.B(n_523),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_1961),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_1984),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2041),
.B(n_526),
.Y(n_2485)
);

OAI21xp5_ASAP7_75t_L g2486 ( 
.A1(n_1937),
.A2(n_527),
.B(n_530),
.Y(n_2486)
);

AND2x4_ASAP7_75t_L g2487 ( 
.A(n_1987),
.B(n_531),
.Y(n_2487)
);

BUFx12f_ASAP7_75t_L g2488 ( 
.A(n_1867),
.Y(n_2488)
);

A2O1A1Ixp33_ASAP7_75t_L g2489 ( 
.A1(n_2060),
.A2(n_533),
.B(n_531),
.C(n_532),
.Y(n_2489)
);

AND3x4_ASAP7_75t_L g2490 ( 
.A(n_1927),
.B(n_2056),
.C(n_1831),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_1917),
.B(n_532),
.Y(n_2491)
);

OAI21xp5_ASAP7_75t_L g2492 ( 
.A1(n_1934),
.A2(n_533),
.B(n_534),
.Y(n_2492)
);

BUFx12f_ASAP7_75t_L g2493 ( 
.A(n_1973),
.Y(n_2493)
);

AOI22xp33_ASAP7_75t_L g2494 ( 
.A1(n_2431),
.A2(n_1869),
.B1(n_2164),
.B2(n_2052),
.Y(n_2494)
);

INVx4_ASAP7_75t_L g2495 ( 
.A(n_2180),
.Y(n_2495)
);

BUFx2_ASAP7_75t_L g2496 ( 
.A(n_2378),
.Y(n_2496)
);

OR2x6_ASAP7_75t_L g2497 ( 
.A(n_2235),
.B(n_2006),
.Y(n_2497)
);

O2A1O1Ixp33_ASAP7_75t_L g2498 ( 
.A1(n_2225),
.A2(n_1979),
.B(n_1954),
.C(n_1899),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2337),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2197),
.Y(n_2500)
);

BUFx2_ASAP7_75t_L g2501 ( 
.A(n_2378),
.Y(n_2501)
);

CKINVDCx20_ASAP7_75t_R g2502 ( 
.A(n_2238),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_2317),
.Y(n_2503)
);

INVx3_ASAP7_75t_L g2504 ( 
.A(n_2238),
.Y(n_2504)
);

OAI22xp5_ASAP7_75t_L g2505 ( 
.A1(n_2414),
.A2(n_2084),
.B1(n_2097),
.B2(n_2090),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2198),
.Y(n_2506)
);

INVx3_ASAP7_75t_L g2507 ( 
.A(n_2227),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2401),
.B(n_1821),
.Y(n_2508)
);

INVxp67_ASAP7_75t_L g2509 ( 
.A(n_2186),
.Y(n_2509)
);

BUFx2_ASAP7_75t_L g2510 ( 
.A(n_2323),
.Y(n_2510)
);

OR2x6_ASAP7_75t_L g2511 ( 
.A(n_2299),
.B(n_1982),
.Y(n_2511)
);

OR2x2_ASAP7_75t_L g2512 ( 
.A(n_2191),
.B(n_1813),
.Y(n_2512)
);

O2A1O1Ixp33_ASAP7_75t_L g2513 ( 
.A1(n_2249),
.A2(n_1858),
.B(n_1890),
.C(n_2126),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2205),
.Y(n_2514)
);

INVx1_ASAP7_75t_SL g2515 ( 
.A(n_2182),
.Y(n_2515)
);

INVx3_ASAP7_75t_L g2516 ( 
.A(n_2377),
.Y(n_2516)
);

OAI22xp5_ASAP7_75t_L g2517 ( 
.A1(n_2323),
.A2(n_2161),
.B1(n_2158),
.B2(n_2027),
.Y(n_2517)
);

BUFx2_ASAP7_75t_L g2518 ( 
.A(n_2185),
.Y(n_2518)
);

AOI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2187),
.A2(n_2023),
.B1(n_2059),
.B2(n_2044),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2217),
.Y(n_2520)
);

AND2x2_ASAP7_75t_L g2521 ( 
.A(n_2448),
.B(n_2020),
.Y(n_2521)
);

BUFx6f_ASAP7_75t_L g2522 ( 
.A(n_2377),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2229),
.Y(n_2523)
);

AOI22xp5_ASAP7_75t_L g2524 ( 
.A1(n_2490),
.A2(n_2094),
.B1(n_2115),
.B2(n_2081),
.Y(n_2524)
);

BUFx6f_ASAP7_75t_L g2525 ( 
.A(n_2188),
.Y(n_2525)
);

AOI22xp5_ASAP7_75t_L g2526 ( 
.A1(n_2285),
.A2(n_2120),
.B1(n_2147),
.B2(n_2124),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2244),
.Y(n_2527)
);

AOI21xp5_ASAP7_75t_L g2528 ( 
.A1(n_2465),
.A2(n_2110),
.B(n_2108),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2218),
.B(n_2029),
.Y(n_2529)
);

CKINVDCx16_ASAP7_75t_R g2530 ( 
.A(n_2476),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2241),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2257),
.Y(n_2532)
);

AND2x4_ASAP7_75t_L g2533 ( 
.A(n_2254),
.B(n_1994),
.Y(n_2533)
);

INVx5_ASAP7_75t_L g2534 ( 
.A(n_2358),
.Y(n_2534)
);

OAI22xp5_ASAP7_75t_L g2535 ( 
.A1(n_2376),
.A2(n_2177),
.B1(n_2173),
.B2(n_1892),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2258),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2267),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2285),
.B(n_2288),
.Y(n_2538)
);

INVx3_ASAP7_75t_L g2539 ( 
.A(n_2358),
.Y(n_2539)
);

AND2x2_ASAP7_75t_SL g2540 ( 
.A(n_2288),
.B(n_1815),
.Y(n_2540)
);

OR2x6_ASAP7_75t_L g2541 ( 
.A(n_2476),
.B(n_2269),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2284),
.B(n_2159),
.Y(n_2542)
);

AOI21xp5_ASAP7_75t_L g2543 ( 
.A1(n_2347),
.A2(n_2117),
.B(n_2116),
.Y(n_2543)
);

AND2x2_ASAP7_75t_L g2544 ( 
.A(n_2329),
.B(n_2036),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2292),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2287),
.B(n_2165),
.Y(n_2546)
);

BUFx10_ASAP7_75t_L g2547 ( 
.A(n_2382),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2305),
.B(n_2166),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2309),
.Y(n_2549)
);

OAI22xp5_ASAP7_75t_L g2550 ( 
.A1(n_2353),
.A2(n_1894),
.B1(n_1913),
.B2(n_1989),
.Y(n_2550)
);

A2O1A1Ixp33_ASAP7_75t_SL g2551 ( 
.A1(n_2237),
.A2(n_1919),
.B(n_1978),
.C(n_2089),
.Y(n_2551)
);

BUFx2_ASAP7_75t_L g2552 ( 
.A(n_2356),
.Y(n_2552)
);

AND2x4_ASAP7_75t_L g2553 ( 
.A(n_2286),
.B(n_1957),
.Y(n_2553)
);

INVx3_ASAP7_75t_L g2554 ( 
.A(n_2339),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2316),
.Y(n_2555)
);

AOI22xp5_ASAP7_75t_L g2556 ( 
.A1(n_2331),
.A2(n_1998),
.B1(n_1900),
.B2(n_1929),
.Y(n_2556)
);

OR2x2_ASAP7_75t_SL g2557 ( 
.A(n_2283),
.B(n_1936),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2236),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2325),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_SL g2560 ( 
.A(n_2445),
.B(n_1879),
.Y(n_2560)
);

NOR2xp33_ASAP7_75t_L g2561 ( 
.A(n_2493),
.B(n_1959),
.Y(n_2561)
);

CKINVDCx5p33_ASAP7_75t_R g2562 ( 
.A(n_2386),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2369),
.Y(n_2563)
);

INVx3_ASAP7_75t_L g2564 ( 
.A(n_2339),
.Y(n_2564)
);

A2O1A1Ixp33_ASAP7_75t_SL g2565 ( 
.A1(n_2243),
.A2(n_2183),
.B(n_2367),
.C(n_2366),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2447),
.Y(n_2566)
);

AOI22xp5_ASAP7_75t_L g2567 ( 
.A1(n_2415),
.A2(n_2144),
.B1(n_2145),
.B2(n_2143),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2242),
.Y(n_2568)
);

AND2x2_ASAP7_75t_L g2569 ( 
.A(n_2279),
.B(n_534),
.Y(n_2569)
);

CKINVDCx11_ASAP7_75t_R g2570 ( 
.A(n_2271),
.Y(n_2570)
);

OR2x2_ASAP7_75t_L g2571 ( 
.A(n_2388),
.B(n_2162),
.Y(n_2571)
);

CKINVDCx5p33_ASAP7_75t_R g2572 ( 
.A(n_2418),
.Y(n_2572)
);

INVx1_ASAP7_75t_SL g2573 ( 
.A(n_2308),
.Y(n_2573)
);

INVxp67_ASAP7_75t_L g2574 ( 
.A(n_2270),
.Y(n_2574)
);

BUFx12f_ASAP7_75t_L g2575 ( 
.A(n_2361),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_SL g2576 ( 
.A(n_2245),
.B(n_2174),
.Y(n_2576)
);

AOI22xp33_ASAP7_75t_SL g2577 ( 
.A1(n_2488),
.A2(n_2175),
.B1(n_536),
.B2(n_534),
.Y(n_2577)
);

AND2x2_ASAP7_75t_L g2578 ( 
.A(n_2280),
.B(n_535),
.Y(n_2578)
);

BUFx12f_ASAP7_75t_L g2579 ( 
.A(n_2349),
.Y(n_2579)
);

OAI21xp33_ASAP7_75t_L g2580 ( 
.A1(n_2220),
.A2(n_538),
.B(n_539),
.Y(n_2580)
);

AOI22xp5_ASAP7_75t_L g2581 ( 
.A1(n_2415),
.A2(n_542),
.B1(n_539),
.B2(n_540),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2263),
.Y(n_2582)
);

AOI221x1_ASAP7_75t_L g2583 ( 
.A1(n_2380),
.A2(n_543),
.B1(n_540),
.B2(n_542),
.C(n_544),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2328),
.B(n_542),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2276),
.Y(n_2585)
);

AND2x4_ASAP7_75t_L g2586 ( 
.A(n_2304),
.B(n_543),
.Y(n_2586)
);

INVx4_ASAP7_75t_L g2587 ( 
.A(n_2277),
.Y(n_2587)
);

BUFx6f_ASAP7_75t_L g2588 ( 
.A(n_2188),
.Y(n_2588)
);

AND2x2_ASAP7_75t_L g2589 ( 
.A(n_2332),
.B(n_544),
.Y(n_2589)
);

AO21x1_ASAP7_75t_L g2590 ( 
.A1(n_2444),
.A2(n_544),
.B(n_545),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2426),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2298),
.Y(n_2592)
);

AND2x4_ASAP7_75t_L g2593 ( 
.A(n_2201),
.B(n_545),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2335),
.B(n_545),
.Y(n_2594)
);

BUFx4f_ASAP7_75t_SL g2595 ( 
.A(n_2277),
.Y(n_2595)
);

AOI21xp5_ASAP7_75t_L g2596 ( 
.A1(n_2240),
.A2(n_546),
.B(n_547),
.Y(n_2596)
);

AOI21xp5_ASAP7_75t_L g2597 ( 
.A1(n_2291),
.A2(n_546),
.B(n_547),
.Y(n_2597)
);

OR2x2_ASAP7_75t_L g2598 ( 
.A(n_2223),
.B(n_2359),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2352),
.B(n_546),
.Y(n_2599)
);

CKINVDCx20_ASAP7_75t_R g2600 ( 
.A(n_2399),
.Y(n_2600)
);

BUFx6f_ASAP7_75t_L g2601 ( 
.A(n_2188),
.Y(n_2601)
);

AOI21xp5_ASAP7_75t_L g2602 ( 
.A1(n_2293),
.A2(n_548),
.B(n_549),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2302),
.Y(n_2603)
);

INVxp67_ASAP7_75t_SL g2604 ( 
.A(n_2428),
.Y(n_2604)
);

INVx4_ASAP7_75t_L g2605 ( 
.A(n_2363),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2398),
.B(n_549),
.Y(n_2606)
);

CKINVDCx8_ASAP7_75t_R g2607 ( 
.A(n_2415),
.Y(n_2607)
);

AND2x4_ASAP7_75t_L g2608 ( 
.A(n_2446),
.B(n_550),
.Y(n_2608)
);

OR2x6_ASAP7_75t_L g2609 ( 
.A(n_2313),
.B(n_552),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2336),
.B(n_552),
.Y(n_2610)
);

AND2x4_ASAP7_75t_L g2611 ( 
.A(n_2451),
.B(n_552),
.Y(n_2611)
);

OAI21x1_ASAP7_75t_L g2612 ( 
.A1(n_2315),
.A2(n_553),
.B(n_554),
.Y(n_2612)
);

OR2x6_ASAP7_75t_L g2613 ( 
.A(n_2312),
.B(n_553),
.Y(n_2613)
);

AND2x4_ASAP7_75t_L g2614 ( 
.A(n_2451),
.B(n_553),
.Y(n_2614)
);

INVx5_ASAP7_75t_L g2615 ( 
.A(n_2251),
.Y(n_2615)
);

INVx4_ASAP7_75t_L g2616 ( 
.A(n_2371),
.Y(n_2616)
);

INVx2_ASAP7_75t_SL g2617 ( 
.A(n_2371),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2210),
.B(n_2226),
.Y(n_2618)
);

AOI22xp33_ASAP7_75t_SL g2619 ( 
.A1(n_2289),
.A2(n_558),
.B1(n_556),
.B2(n_557),
.Y(n_2619)
);

CKINVDCx5p33_ASAP7_75t_R g2620 ( 
.A(n_2456),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2228),
.B(n_557),
.Y(n_2621)
);

INVx2_ASAP7_75t_SL g2622 ( 
.A(n_2395),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2181),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2350),
.B(n_559),
.Y(n_2624)
);

BUFx2_ASAP7_75t_SL g2625 ( 
.A(n_2405),
.Y(n_2625)
);

BUFx4f_ASAP7_75t_L g2626 ( 
.A(n_2314),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2192),
.Y(n_2627)
);

BUFx2_ASAP7_75t_L g2628 ( 
.A(n_2393),
.Y(n_2628)
);

O2A1O1Ixp5_ASAP7_75t_L g2629 ( 
.A1(n_2407),
.A2(n_561),
.B(n_559),
.C(n_560),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2202),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2357),
.B(n_559),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2384),
.B(n_560),
.Y(n_2632)
);

INVx3_ASAP7_75t_L g2633 ( 
.A(n_2438),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2439),
.B(n_2457),
.Y(n_2634)
);

INVx4_ASAP7_75t_L g2635 ( 
.A(n_2438),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2246),
.B(n_562),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2330),
.B(n_565),
.Y(n_2637)
);

BUFx6f_ASAP7_75t_L g2638 ( 
.A(n_2251),
.Y(n_2638)
);

O2A1O1Ixp5_ASAP7_75t_L g2639 ( 
.A1(n_2194),
.A2(n_567),
.B(n_565),
.C(n_566),
.Y(n_2639)
);

AND2x4_ASAP7_75t_L g2640 ( 
.A(n_2341),
.B(n_566),
.Y(n_2640)
);

AOI21xp5_ASAP7_75t_L g2641 ( 
.A1(n_2463),
.A2(n_2208),
.B(n_2207),
.Y(n_2641)
);

AOI21xp5_ASAP7_75t_L g2642 ( 
.A1(n_2211),
.A2(n_566),
.B(n_567),
.Y(n_2642)
);

AOI21xp5_ASAP7_75t_L g2643 ( 
.A1(n_2224),
.A2(n_567),
.B(n_568),
.Y(n_2643)
);

BUFx4f_ASAP7_75t_L g2644 ( 
.A(n_2470),
.Y(n_2644)
);

OAI22xp5_ASAP7_75t_SL g2645 ( 
.A1(n_2234),
.A2(n_572),
.B1(n_569),
.B2(n_570),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2318),
.Y(n_2646)
);

CKINVDCx5p33_ASAP7_75t_R g2647 ( 
.A(n_2480),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2326),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2485),
.B(n_572),
.Y(n_2649)
);

AOI22xp5_ASAP7_75t_L g2650 ( 
.A1(n_2250),
.A2(n_575),
.B1(n_573),
.B2(n_574),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_2466),
.B(n_574),
.Y(n_2651)
);

INVx1_ASAP7_75t_SL g2652 ( 
.A(n_2190),
.Y(n_2652)
);

AOI21xp5_ASAP7_75t_L g2653 ( 
.A1(n_2230),
.A2(n_575),
.B(n_576),
.Y(n_2653)
);

INVx3_ASAP7_75t_L g2654 ( 
.A(n_2402),
.Y(n_2654)
);

AND2x4_ASAP7_75t_L g2655 ( 
.A(n_2459),
.B(n_576),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_SL g2656 ( 
.A(n_2345),
.B(n_576),
.Y(n_2656)
);

BUFx12f_ASAP7_75t_L g2657 ( 
.A(n_2264),
.Y(n_2657)
);

BUFx6f_ASAP7_75t_L g2658 ( 
.A(n_2256),
.Y(n_2658)
);

BUFx6f_ASAP7_75t_L g2659 ( 
.A(n_2256),
.Y(n_2659)
);

INVx2_ASAP7_75t_SL g2660 ( 
.A(n_2272),
.Y(n_2660)
);

AOI21xp5_ASAP7_75t_L g2661 ( 
.A1(n_2231),
.A2(n_577),
.B(n_578),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2360),
.Y(n_2662)
);

AOI21xp5_ASAP7_75t_L g2663 ( 
.A1(n_2233),
.A2(n_577),
.B(n_579),
.Y(n_2663)
);

O2A1O1Ixp33_ASAP7_75t_L g2664 ( 
.A1(n_2473),
.A2(n_581),
.B(n_579),
.C(n_580),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2307),
.Y(n_2665)
);

AND2x4_ASAP7_75t_L g2666 ( 
.A(n_2381),
.B(n_581),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2479),
.B(n_2484),
.Y(n_2667)
);

A2O1A1Ixp33_ASAP7_75t_L g2668 ( 
.A1(n_2273),
.A2(n_603),
.B(n_601),
.C(n_602),
.Y(n_2668)
);

OA21x2_ASAP7_75t_L g2669 ( 
.A1(n_2343),
.A2(n_603),
.B(n_604),
.Y(n_2669)
);

INVxp67_ASAP7_75t_SL g2670 ( 
.A(n_2281),
.Y(n_2670)
);

OAI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2468),
.A2(n_608),
.B1(n_605),
.B2(n_607),
.Y(n_2671)
);

INVx3_ASAP7_75t_L g2672 ( 
.A(n_2295),
.Y(n_2672)
);

CKINVDCx5p33_ASAP7_75t_R g2673 ( 
.A(n_2219),
.Y(n_2673)
);

NAND2x1_ASAP7_75t_L g2674 ( 
.A(n_2300),
.B(n_609),
.Y(n_2674)
);

AOI22xp5_ASAP7_75t_L g2675 ( 
.A1(n_2420),
.A2(n_611),
.B1(n_609),
.B2(n_610),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2333),
.Y(n_2676)
);

NOR2x1_ASAP7_75t_SL g2677 ( 
.A(n_2409),
.B(n_614),
.Y(n_2677)
);

BUFx2_ASAP7_75t_L g2678 ( 
.A(n_2214),
.Y(n_2678)
);

INVx3_ASAP7_75t_L g2679 ( 
.A(n_2214),
.Y(n_2679)
);

AOI22xp33_ASAP7_75t_L g2680 ( 
.A1(n_2222),
.A2(n_617),
.B1(n_615),
.B2(n_616),
.Y(n_2680)
);

O2A1O1Ixp33_ASAP7_75t_L g2681 ( 
.A1(n_2474),
.A2(n_618),
.B(n_615),
.C(n_617),
.Y(n_2681)
);

NAND2xp33_ASAP7_75t_L g2682 ( 
.A(n_2338),
.B(n_618),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2375),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2206),
.B(n_2483),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2481),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2464),
.B(n_619),
.Y(n_2686)
);

INVxp67_ASAP7_75t_L g2687 ( 
.A(n_2320),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2385),
.Y(n_2688)
);

NOR2xp33_ASAP7_75t_L g2689 ( 
.A(n_2478),
.B(n_620),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2481),
.Y(n_2690)
);

OR2x6_ASAP7_75t_L g2691 ( 
.A(n_2278),
.B(n_620),
.Y(n_2691)
);

INVx2_ASAP7_75t_SL g2692 ( 
.A(n_2290),
.Y(n_2692)
);

INVxp67_ASAP7_75t_SL g2693 ( 
.A(n_2281),
.Y(n_2693)
);

OR2x6_ASAP7_75t_L g2694 ( 
.A(n_2482),
.B(n_622),
.Y(n_2694)
);

O2A1O1Ixp33_ASAP7_75t_L g2695 ( 
.A1(n_2213),
.A2(n_625),
.B(n_623),
.C(n_624),
.Y(n_2695)
);

AND2x4_ASAP7_75t_L g2696 ( 
.A(n_2397),
.B(n_625),
.Y(n_2696)
);

INVx2_ASAP7_75t_L g2697 ( 
.A(n_2400),
.Y(n_2697)
);

A2O1A1Ixp33_ASAP7_75t_SL g2698 ( 
.A1(n_2354),
.A2(n_628),
.B(n_626),
.C(n_627),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2351),
.B(n_786),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2262),
.Y(n_2700)
);

O2A1O1Ixp33_ASAP7_75t_L g2701 ( 
.A1(n_2491),
.A2(n_632),
.B(n_627),
.C(n_629),
.Y(n_2701)
);

HB1xp67_ASAP7_75t_L g2702 ( 
.A(n_2487),
.Y(n_2702)
);

AND2x4_ASAP7_75t_L g2703 ( 
.A(n_2346),
.B(n_785),
.Y(n_2703)
);

A2O1A1Ixp33_ASAP7_75t_L g2704 ( 
.A1(n_2189),
.A2(n_635),
.B(n_633),
.C(n_634),
.Y(n_2704)
);

BUFx6f_ASAP7_75t_L g2705 ( 
.A(n_2364),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2500),
.Y(n_2706)
);

OAI22xp5_ASAP7_75t_L g2707 ( 
.A1(n_2607),
.A2(n_2391),
.B1(n_2461),
.B2(n_2368),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2499),
.Y(n_2708)
);

AND2x4_ASAP7_75t_L g2709 ( 
.A(n_2605),
.B(n_2346),
.Y(n_2709)
);

AOI22xp33_ASAP7_75t_L g2710 ( 
.A1(n_2626),
.A2(n_2275),
.B1(n_2387),
.B2(n_2475),
.Y(n_2710)
);

AOI21x1_ASAP7_75t_L g2711 ( 
.A1(n_2662),
.A2(n_2212),
.B(n_2261),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2506),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2634),
.B(n_2618),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2514),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2520),
.Y(n_2715)
);

AND2x2_ASAP7_75t_L g2716 ( 
.A(n_2569),
.B(n_2383),
.Y(n_2716)
);

NAND2x1p5_ASAP7_75t_L g2717 ( 
.A(n_2534),
.B(n_2467),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2523),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2531),
.Y(n_2719)
);

BUFx12f_ASAP7_75t_L g2720 ( 
.A(n_2570),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2558),
.B(n_2450),
.Y(n_2721)
);

AO21x1_ASAP7_75t_SL g2722 ( 
.A1(n_2702),
.A2(n_2303),
.B(n_2310),
.Y(n_2722)
);

INVx5_ASAP7_75t_L g2723 ( 
.A(n_2575),
.Y(n_2723)
);

INVx3_ASAP7_75t_L g2724 ( 
.A(n_2534),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2536),
.Y(n_2725)
);

BUFx2_ASAP7_75t_L g2726 ( 
.A(n_2628),
.Y(n_2726)
);

INVx3_ASAP7_75t_L g2727 ( 
.A(n_2495),
.Y(n_2727)
);

INVx6_ASAP7_75t_L g2728 ( 
.A(n_2579),
.Y(n_2728)
);

INVx3_ASAP7_75t_L g2729 ( 
.A(n_2539),
.Y(n_2729)
);

CKINVDCx20_ASAP7_75t_R g2730 ( 
.A(n_2502),
.Y(n_2730)
);

BUFx2_ASAP7_75t_L g2731 ( 
.A(n_2670),
.Y(n_2731)
);

CKINVDCx6p67_ASAP7_75t_R g2732 ( 
.A(n_2600),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2527),
.Y(n_2733)
);

AND2x2_ASAP7_75t_L g2734 ( 
.A(n_2578),
.B(n_2589),
.Y(n_2734)
);

INVx6_ASAP7_75t_L g2735 ( 
.A(n_2522),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2537),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2652),
.B(n_2425),
.Y(n_2737)
);

AOI22xp33_ASAP7_75t_L g2738 ( 
.A1(n_2560),
.A2(n_2429),
.B1(n_2322),
.B2(n_2239),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2549),
.Y(n_2739)
);

BUFx3_ASAP7_75t_L g2740 ( 
.A(n_2507),
.Y(n_2740)
);

OR2x6_ASAP7_75t_L g2741 ( 
.A(n_2541),
.B(n_2452),
.Y(n_2741)
);

AOI22xp33_ASAP7_75t_SL g2742 ( 
.A1(n_2540),
.A2(n_2394),
.B1(n_2260),
.B2(n_2282),
.Y(n_2742)
);

BUFx6f_ASAP7_75t_L g2743 ( 
.A(n_2522),
.Y(n_2743)
);

INVx2_ASAP7_75t_SL g2744 ( 
.A(n_2504),
.Y(n_2744)
);

CKINVDCx5p33_ASAP7_75t_R g2745 ( 
.A(n_2503),
.Y(n_2745)
);

BUFx2_ASAP7_75t_R g2746 ( 
.A(n_2562),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2532),
.Y(n_2747)
);

OAI22xp33_ASAP7_75t_L g2748 ( 
.A1(n_2694),
.A2(n_2266),
.B1(n_2374),
.B2(n_2319),
.Y(n_2748)
);

OA21x2_ASAP7_75t_L g2749 ( 
.A1(n_2685),
.A2(n_2454),
.B(n_2453),
.Y(n_2749)
);

CKINVDCx20_ASAP7_75t_R g2750 ( 
.A(n_2572),
.Y(n_2750)
);

OAI21x1_ASAP7_75t_SL g2751 ( 
.A1(n_2590),
.A2(n_2253),
.B(n_2392),
.Y(n_2751)
);

OAI21x1_ASAP7_75t_L g2752 ( 
.A1(n_2697),
.A2(n_2265),
.B(n_2209),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2555),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2566),
.Y(n_2754)
);

INVx1_ASAP7_75t_SL g2755 ( 
.A(n_2573),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2545),
.Y(n_2756)
);

INVx3_ASAP7_75t_L g2757 ( 
.A(n_2644),
.Y(n_2757)
);

OAI22xp5_ASAP7_75t_L g2758 ( 
.A1(n_2581),
.A2(n_2301),
.B1(n_2324),
.B2(n_2294),
.Y(n_2758)
);

BUFx12f_ASAP7_75t_L g2759 ( 
.A(n_2547),
.Y(n_2759)
);

INVxp33_ASAP7_75t_L g2760 ( 
.A(n_2538),
.Y(n_2760)
);

CKINVDCx5p33_ASAP7_75t_R g2761 ( 
.A(n_2541),
.Y(n_2761)
);

INVx1_ASAP7_75t_SL g2762 ( 
.A(n_2595),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2559),
.Y(n_2763)
);

INVx4_ASAP7_75t_L g2764 ( 
.A(n_2609),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2563),
.Y(n_2765)
);

INVx3_ASAP7_75t_L g2766 ( 
.A(n_2616),
.Y(n_2766)
);

BUFx3_ASAP7_75t_L g2767 ( 
.A(n_2552),
.Y(n_2767)
);

OAI21x1_ASAP7_75t_L g2768 ( 
.A1(n_2591),
.A2(n_2196),
.B(n_2195),
.Y(n_2768)
);

AOI22xp33_ASAP7_75t_L g2769 ( 
.A1(n_2497),
.A2(n_2424),
.B1(n_2342),
.B2(n_2421),
.Y(n_2769)
);

BUFx4f_ASAP7_75t_L g2770 ( 
.A(n_2609),
.Y(n_2770)
);

OA21x2_ASAP7_75t_L g2771 ( 
.A1(n_2690),
.A2(n_2460),
.B(n_2373),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2686),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2669),
.Y(n_2773)
);

OR2x6_ASAP7_75t_L g2774 ( 
.A(n_2694),
.B(n_2204),
.Y(n_2774)
);

AOI22xp33_ASAP7_75t_L g2775 ( 
.A1(n_2497),
.A2(n_2691),
.B1(n_2505),
.B2(n_2544),
.Y(n_2775)
);

AOI22xp33_ASAP7_75t_SL g2776 ( 
.A1(n_2673),
.A2(n_2477),
.B1(n_2492),
.B2(n_2486),
.Y(n_2776)
);

OAI21xp33_ASAP7_75t_L g2777 ( 
.A1(n_2494),
.A2(n_2410),
.B(n_2311),
.Y(n_2777)
);

AND2x2_ASAP7_75t_L g2778 ( 
.A(n_2594),
.B(n_2396),
.Y(n_2778)
);

BUFx2_ASAP7_75t_L g2779 ( 
.A(n_2693),
.Y(n_2779)
);

INVx1_ASAP7_75t_SL g2780 ( 
.A(n_2518),
.Y(n_2780)
);

BUFx2_ASAP7_75t_L g2781 ( 
.A(n_2635),
.Y(n_2781)
);

HB1xp67_ASAP7_75t_L g2782 ( 
.A(n_2574),
.Y(n_2782)
);

BUFx4f_ASAP7_75t_SL g2783 ( 
.A(n_2515),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2667),
.Y(n_2784)
);

NAND2x1p5_ASAP7_75t_L g2785 ( 
.A(n_2587),
.B(n_2362),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2665),
.Y(n_2786)
);

OAI22xp5_ASAP7_75t_L g2787 ( 
.A1(n_2619),
.A2(n_2344),
.B1(n_2489),
.B2(n_2390),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2509),
.B(n_2412),
.Y(n_2788)
);

BUFx4f_ASAP7_75t_L g2789 ( 
.A(n_2613),
.Y(n_2789)
);

AO21x2_ASAP7_75t_L g2790 ( 
.A1(n_2683),
.A2(n_2419),
.B(n_2296),
.Y(n_2790)
);

AOI22xp33_ASAP7_75t_L g2791 ( 
.A1(n_2561),
.A2(n_2469),
.B1(n_2472),
.B2(n_2455),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2584),
.Y(n_2792)
);

AND2x2_ASAP7_75t_L g2793 ( 
.A(n_2599),
.B(n_635),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2610),
.Y(n_2794)
);

INVx6_ASAP7_75t_L g2795 ( 
.A(n_2530),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2624),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2631),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2632),
.Y(n_2798)
);

AND2x2_ASAP7_75t_L g2799 ( 
.A(n_2606),
.B(n_636),
.Y(n_2799)
);

NAND2x1p5_ASAP7_75t_L g2800 ( 
.A(n_2510),
.B(n_2615),
.Y(n_2800)
);

INVx4_ASAP7_75t_L g2801 ( 
.A(n_2516),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2612),
.Y(n_2802)
);

CKINVDCx5p33_ASAP7_75t_R g2803 ( 
.A(n_2620),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2623),
.Y(n_2804)
);

OAI22xp5_ASAP7_75t_L g2805 ( 
.A1(n_2556),
.A2(n_2675),
.B1(n_2680),
.B2(n_2524),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2627),
.Y(n_2806)
);

OA21x2_ASAP7_75t_L g2807 ( 
.A1(n_2700),
.A2(n_2200),
.B(n_2199),
.Y(n_2807)
);

OAI21x1_ASAP7_75t_L g2808 ( 
.A1(n_2646),
.A2(n_2306),
.B(n_2334),
.Y(n_2808)
);

BUFx2_ASAP7_75t_L g2809 ( 
.A(n_2525),
.Y(n_2809)
);

BUFx2_ASAP7_75t_L g2810 ( 
.A(n_2525),
.Y(n_2810)
);

OAI22xp5_ASAP7_75t_L g2811 ( 
.A1(n_2577),
.A2(n_2417),
.B1(n_2434),
.B2(n_2389),
.Y(n_2811)
);

OAI21xp5_ASAP7_75t_SL g2812 ( 
.A1(n_2519),
.A2(n_2435),
.B(n_2355),
.Y(n_2812)
);

INVx3_ASAP7_75t_L g2813 ( 
.A(n_2654),
.Y(n_2813)
);

INVx3_ASAP7_75t_L g2814 ( 
.A(n_2554),
.Y(n_2814)
);

INVx3_ASAP7_75t_L g2815 ( 
.A(n_2564),
.Y(n_2815)
);

BUFx6f_ASAP7_75t_L g2816 ( 
.A(n_2588),
.Y(n_2816)
);

OR2x2_ASAP7_75t_L g2817 ( 
.A(n_2598),
.B(n_2427),
.Y(n_2817)
);

AOI22xp5_ASAP7_75t_L g2818 ( 
.A1(n_2645),
.A2(n_2370),
.B1(n_2372),
.B2(n_2365),
.Y(n_2818)
);

INVx3_ASAP7_75t_L g2819 ( 
.A(n_2611),
.Y(n_2819)
);

CKINVDCx11_ASAP7_75t_R g2820 ( 
.A(n_2657),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2630),
.Y(n_2821)
);

INVx2_ASAP7_75t_SL g2822 ( 
.A(n_2496),
.Y(n_2822)
);

BUFx6f_ASAP7_75t_L g2823 ( 
.A(n_2588),
.Y(n_2823)
);

HB1xp67_ASAP7_75t_L g2824 ( 
.A(n_2604),
.Y(n_2824)
);

INVx3_ASAP7_75t_L g2825 ( 
.A(n_2614),
.Y(n_2825)
);

CKINVDCx5p33_ASAP7_75t_R g2826 ( 
.A(n_2647),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2568),
.Y(n_2827)
);

OAI22xp5_ASAP7_75t_L g2828 ( 
.A1(n_2526),
.A2(n_2430),
.B1(n_2379),
.B2(n_2411),
.Y(n_2828)
);

OAI21x1_ASAP7_75t_L g2829 ( 
.A1(n_2648),
.A2(n_2340),
.B(n_2252),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2582),
.Y(n_2830)
);

INVx1_ASAP7_75t_SL g2831 ( 
.A(n_2501),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2585),
.Y(n_2832)
);

INVx5_ASAP7_75t_L g2833 ( 
.A(n_2601),
.Y(n_2833)
);

AOI21x1_ASAP7_75t_L g2834 ( 
.A1(n_2688),
.A2(n_2247),
.B(n_2232),
.Y(n_2834)
);

OAI22xp5_ASAP7_75t_L g2835 ( 
.A1(n_2650),
.A2(n_2408),
.B1(n_2416),
.B2(n_2413),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2592),
.Y(n_2836)
);

BUFx12f_ASAP7_75t_L g2837 ( 
.A(n_2660),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2603),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2542),
.Y(n_2839)
);

INVx4_ASAP7_75t_L g2840 ( 
.A(n_2633),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2638),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2638),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2546),
.Y(n_2843)
);

HB1xp67_ASAP7_75t_L g2844 ( 
.A(n_2617),
.Y(n_2844)
);

OAI21x1_ASAP7_75t_L g2845 ( 
.A1(n_2676),
.A2(n_2348),
.B(n_2248),
.Y(n_2845)
);

BUFx8_ASAP7_75t_L g2846 ( 
.A(n_2586),
.Y(n_2846)
);

HB1xp67_ASAP7_75t_L g2847 ( 
.A(n_2622),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2548),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2684),
.Y(n_2849)
);

NAND2x1p5_ASAP7_75t_L g2850 ( 
.A(n_2723),
.B(n_2593),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2708),
.Y(n_2851)
);

HB1xp67_ASAP7_75t_L g2852 ( 
.A(n_2824),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2749),
.Y(n_2853)
);

INVx5_ASAP7_75t_L g2854 ( 
.A(n_2795),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2749),
.Y(n_2855)
);

OR2x2_ASAP7_75t_L g2856 ( 
.A(n_2726),
.B(n_2512),
.Y(n_2856)
);

HB1xp67_ASAP7_75t_L g2857 ( 
.A(n_2726),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2712),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2714),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2715),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2718),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2839),
.Y(n_2862)
);

INVx3_ASAP7_75t_L g2863 ( 
.A(n_2731),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2843),
.Y(n_2864)
);

INVx2_ASAP7_75t_SL g2865 ( 
.A(n_2795),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2848),
.Y(n_2866)
);

HB1xp67_ASAP7_75t_L g2867 ( 
.A(n_2782),
.Y(n_2867)
);

AND2x2_ASAP7_75t_L g2868 ( 
.A(n_2734),
.B(n_2649),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2733),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2706),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2747),
.Y(n_2871)
);

OA21x2_ASAP7_75t_L g2872 ( 
.A1(n_2752),
.A2(n_2641),
.B(n_2528),
.Y(n_2872)
);

AO21x2_ASAP7_75t_L g2873 ( 
.A1(n_2711),
.A2(n_2698),
.B(n_2576),
.Y(n_2873)
);

HB1xp67_ASAP7_75t_L g2874 ( 
.A(n_2779),
.Y(n_2874)
);

AND2x2_ASAP7_75t_L g2875 ( 
.A(n_2713),
.B(n_2621),
.Y(n_2875)
);

CKINVDCx5p33_ASAP7_75t_R g2876 ( 
.A(n_2730),
.Y(n_2876)
);

BUFx2_ASAP7_75t_L g2877 ( 
.A(n_2781),
.Y(n_2877)
);

BUFx3_ASAP7_75t_L g2878 ( 
.A(n_2723),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2719),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2725),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2784),
.B(n_2849),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2736),
.Y(n_2882)
);

BUFx3_ASAP7_75t_L g2883 ( 
.A(n_2723),
.Y(n_2883)
);

INVxp67_ASAP7_75t_L g2884 ( 
.A(n_2767),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2739),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2753),
.Y(n_2886)
);

INVx1_ASAP7_75t_SL g2887 ( 
.A(n_2783),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2754),
.Y(n_2888)
);

AND2x2_ASAP7_75t_L g2889 ( 
.A(n_2760),
.B(n_2778),
.Y(n_2889)
);

INVx2_ASAP7_75t_L g2890 ( 
.A(n_2756),
.Y(n_2890)
);

INVx2_ASAP7_75t_SL g2891 ( 
.A(n_2735),
.Y(n_2891)
);

CKINVDCx20_ASAP7_75t_R g2892 ( 
.A(n_2750),
.Y(n_2892)
);

AND2x4_ASAP7_75t_L g2893 ( 
.A(n_2781),
.B(n_2553),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2763),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2765),
.Y(n_2895)
);

AOI21x1_ASAP7_75t_L g2896 ( 
.A1(n_2834),
.A2(n_2674),
.B(n_2583),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2771),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2830),
.Y(n_2898)
);

CKINVDCx5p33_ASAP7_75t_R g2899 ( 
.A(n_2732),
.Y(n_2899)
);

INVx3_ASAP7_75t_L g2900 ( 
.A(n_2727),
.Y(n_2900)
);

NOR2x1p5_ASAP7_75t_L g2901 ( 
.A(n_2764),
.B(n_2666),
.Y(n_2901)
);

HB1xp67_ASAP7_75t_L g2902 ( 
.A(n_2780),
.Y(n_2902)
);

NAND2x1p5_ASAP7_75t_L g2903 ( 
.A(n_2770),
.B(n_2608),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2804),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2806),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2821),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2827),
.B(n_2687),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2832),
.B(n_2836),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2788),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2773),
.Y(n_2910)
);

BUFx3_ASAP7_75t_L g2911 ( 
.A(n_2740),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2802),
.Y(n_2912)
);

INVx3_ASAP7_75t_L g2913 ( 
.A(n_2813),
.Y(n_2913)
);

INVx3_ASAP7_75t_L g2914 ( 
.A(n_2800),
.Y(n_2914)
);

AND2x2_ASAP7_75t_L g2915 ( 
.A(n_2786),
.B(n_2655),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2838),
.Y(n_2916)
);

AND2x2_ASAP7_75t_L g2917 ( 
.A(n_2793),
.B(n_2529),
.Y(n_2917)
);

AND2x2_ASAP7_75t_L g2918 ( 
.A(n_2799),
.B(n_2521),
.Y(n_2918)
);

INVx1_ASAP7_75t_SL g2919 ( 
.A(n_2761),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2768),
.Y(n_2920)
);

OR2x2_ASAP7_75t_L g2921 ( 
.A(n_2755),
.B(n_2508),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2807),
.Y(n_2922)
);

AOI21xp5_ASAP7_75t_L g2923 ( 
.A1(n_2777),
.A2(n_2565),
.B(n_2656),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2841),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2842),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2809),
.Y(n_2926)
);

HB1xp67_ASAP7_75t_L g2927 ( 
.A(n_2844),
.Y(n_2927)
);

HB1xp67_ASAP7_75t_L g2928 ( 
.A(n_2847),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2716),
.B(n_2640),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_2792),
.B(n_2651),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2808),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2809),
.Y(n_2932)
);

BUFx2_ASAP7_75t_L g2933 ( 
.A(n_2743),
.Y(n_2933)
);

INVx3_ASAP7_75t_L g2934 ( 
.A(n_2801),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2829),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2845),
.Y(n_2936)
);

AO21x2_ASAP7_75t_L g2937 ( 
.A1(n_2751),
.A2(n_2580),
.B(n_2543),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2790),
.Y(n_2938)
);

INVx3_ASAP7_75t_L g2939 ( 
.A(n_2724),
.Y(n_2939)
);

HB1xp67_ASAP7_75t_L g2940 ( 
.A(n_2810),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2721),
.Y(n_2941)
);

OR2x6_ASAP7_75t_L g2942 ( 
.A(n_2774),
.B(n_2625),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2794),
.B(n_2796),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2797),
.B(n_2571),
.Y(n_2944)
);

BUFx6f_ASAP7_75t_L g2945 ( 
.A(n_2743),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2772),
.Y(n_2946)
);

OAI211xp5_ASAP7_75t_L g2947 ( 
.A1(n_2877),
.A2(n_2775),
.B(n_2776),
.C(n_2710),
.Y(n_2947)
);

BUFx2_ASAP7_75t_L g2948 ( 
.A(n_2934),
.Y(n_2948)
);

INVx2_ASAP7_75t_SL g2949 ( 
.A(n_2911),
.Y(n_2949)
);

AND2x4_ASAP7_75t_SL g2950 ( 
.A(n_2934),
.B(n_2766),
.Y(n_2950)
);

INVx3_ASAP7_75t_L g2951 ( 
.A(n_2863),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2916),
.Y(n_2952)
);

AND2x2_ASAP7_75t_L g2953 ( 
.A(n_2889),
.B(n_2819),
.Y(n_2953)
);

OAI221xp5_ASAP7_75t_L g2954 ( 
.A1(n_2942),
.A2(n_2789),
.B1(n_2774),
.B2(n_2791),
.C(n_2742),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2909),
.B(n_2798),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2863),
.Y(n_2956)
);

AND2x2_ASAP7_75t_L g2957 ( 
.A(n_2918),
.B(n_2825),
.Y(n_2957)
);

INVxp67_ASAP7_75t_L g2958 ( 
.A(n_2874),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2916),
.Y(n_2959)
);

AND2x2_ASAP7_75t_L g2960 ( 
.A(n_2917),
.B(n_2817),
.Y(n_2960)
);

AOI22xp33_ASAP7_75t_L g2961 ( 
.A1(n_2942),
.A2(n_2805),
.B1(n_2707),
.B2(n_2748),
.Y(n_2961)
);

HB1xp67_ASAP7_75t_L g2962 ( 
.A(n_2852),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2941),
.B(n_2215),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2851),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2941),
.B(n_2862),
.Y(n_2965)
);

AND2x2_ASAP7_75t_L g2966 ( 
.A(n_2875),
.B(n_2822),
.Y(n_2966)
);

AND2x2_ASAP7_75t_L g2967 ( 
.A(n_2868),
.B(n_2831),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2946),
.Y(n_2968)
);

OR2x2_ASAP7_75t_L g2969 ( 
.A(n_2867),
.B(n_2856),
.Y(n_2969)
);

AOI221x1_ASAP7_75t_L g2970 ( 
.A1(n_2923),
.A2(n_2814),
.B1(n_2815),
.B2(n_2737),
.C(n_2729),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2946),
.Y(n_2971)
);

INVx3_ASAP7_75t_L g2972 ( 
.A(n_2893),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2862),
.B(n_2215),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2864),
.B(n_2215),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2858),
.Y(n_2975)
);

HB1xp67_ASAP7_75t_L g2976 ( 
.A(n_2857),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2864),
.B(n_2216),
.Y(n_2977)
);

INVx2_ASAP7_75t_SL g2978 ( 
.A(n_2878),
.Y(n_2978)
);

BUFx3_ASAP7_75t_L g2979 ( 
.A(n_2883),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2866),
.B(n_2216),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2870),
.Y(n_2981)
);

NOR4xp25_ASAP7_75t_SL g2982 ( 
.A(n_2899),
.B(n_2812),
.C(n_2803),
.D(n_2745),
.Y(n_2982)
);

CKINVDCx5p33_ASAP7_75t_R g2983 ( 
.A(n_2876),
.Y(n_2983)
);

HB1xp67_ASAP7_75t_L g2984 ( 
.A(n_2927),
.Y(n_2984)
);

HB1xp67_ASAP7_75t_L g2985 ( 
.A(n_2928),
.Y(n_2985)
);

BUFx2_ASAP7_75t_L g2986 ( 
.A(n_2900),
.Y(n_2986)
);

AND2x2_ASAP7_75t_L g2987 ( 
.A(n_2929),
.B(n_2902),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2859),
.Y(n_2988)
);

AOI22xp33_ASAP7_75t_L g2989 ( 
.A1(n_2901),
.A2(n_2511),
.B1(n_2722),
.B2(n_2811),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_2940),
.B(n_2744),
.Y(n_2990)
);

AOI221xp5_ASAP7_75t_L g2991 ( 
.A1(n_2930),
.A2(n_2828),
.B1(n_2835),
.B2(n_2689),
.C(n_2787),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2860),
.Y(n_2992)
);

OR2x2_ASAP7_75t_L g2993 ( 
.A(n_2921),
.B(n_2840),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2879),
.Y(n_2994)
);

OR2x2_ASAP7_75t_L g2995 ( 
.A(n_2904),
.B(n_2741),
.Y(n_2995)
);

BUFx2_ASAP7_75t_SL g2996 ( 
.A(n_2854),
.Y(n_2996)
);

AND2x2_ASAP7_75t_L g2997 ( 
.A(n_2908),
.B(n_2837),
.Y(n_2997)
);

AND2x4_ASAP7_75t_L g2998 ( 
.A(n_2926),
.B(n_2741),
.Y(n_2998)
);

AND2x2_ASAP7_75t_L g2999 ( 
.A(n_2907),
.B(n_2932),
.Y(n_2999)
);

AOI21xp5_ASAP7_75t_SL g3000 ( 
.A1(n_2884),
.A2(n_2717),
.B(n_2696),
.Y(n_3000)
);

OR2x2_ASAP7_75t_L g3001 ( 
.A(n_2905),
.B(n_2906),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2861),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2880),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2869),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2871),
.Y(n_3005)
);

AND2x2_ASAP7_75t_L g3006 ( 
.A(n_2882),
.B(n_2678),
.Y(n_3006)
);

CKINVDCx5p33_ASAP7_75t_R g3007 ( 
.A(n_2892),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2885),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_SL g3009 ( 
.A(n_2948),
.B(n_2979),
.Y(n_3009)
);

NOR3xp33_ASAP7_75t_SL g3010 ( 
.A(n_2954),
.B(n_2826),
.C(n_2758),
.Y(n_3010)
);

NAND3xp33_ASAP7_75t_L g3011 ( 
.A(n_2961),
.B(n_2947),
.C(n_2991),
.Y(n_3011)
);

AND2x2_ASAP7_75t_L g3012 ( 
.A(n_2999),
.B(n_2865),
.Y(n_3012)
);

NOR2xp33_ASAP7_75t_L g3013 ( 
.A(n_2949),
.B(n_2887),
.Y(n_3013)
);

AND2x2_ASAP7_75t_SL g3014 ( 
.A(n_2950),
.B(n_2900),
.Y(n_3014)
);

OAI21xp33_ASAP7_75t_L g3015 ( 
.A1(n_2947),
.A2(n_2943),
.B(n_2881),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2962),
.B(n_2898),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_SL g3017 ( 
.A(n_2978),
.B(n_2854),
.Y(n_3017)
);

NAND3xp33_ASAP7_75t_L g3018 ( 
.A(n_2991),
.B(n_2970),
.C(n_2982),
.Y(n_3018)
);

AND2x2_ASAP7_75t_L g3019 ( 
.A(n_2987),
.B(n_2886),
.Y(n_3019)
);

OAI221xp5_ASAP7_75t_L g3020 ( 
.A1(n_2989),
.A2(n_2850),
.B1(n_2738),
.B2(n_2903),
.C(n_2944),
.Y(n_3020)
);

AND2x2_ASAP7_75t_L g3021 ( 
.A(n_2984),
.B(n_2888),
.Y(n_3021)
);

NAND3xp33_ASAP7_75t_L g3022 ( 
.A(n_2976),
.B(n_2958),
.C(n_2985),
.Y(n_3022)
);

OAI22xp5_ASAP7_75t_L g3023 ( 
.A1(n_3000),
.A2(n_2913),
.B1(n_2939),
.B2(n_2914),
.Y(n_3023)
);

AND4x1_ASAP7_75t_L g3024 ( 
.A(n_2997),
.B(n_2746),
.C(n_2720),
.D(n_2728),
.Y(n_3024)
);

AOI211xp5_ASAP7_75t_L g3025 ( 
.A1(n_2986),
.A2(n_2914),
.B(n_2993),
.C(n_2762),
.Y(n_3025)
);

OAI22xp5_ASAP7_75t_L g3026 ( 
.A1(n_2996),
.A2(n_2933),
.B1(n_2557),
.B2(n_2919),
.Y(n_3026)
);

NOR2xp33_ASAP7_75t_R g3027 ( 
.A(n_3007),
.B(n_2757),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_SL g3028 ( 
.A(n_2972),
.B(n_2945),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2960),
.B(n_2890),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2955),
.B(n_2894),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2976),
.B(n_2895),
.Y(n_3031)
);

NAND3xp33_ASAP7_75t_L g3032 ( 
.A(n_2982),
.B(n_2846),
.C(n_2769),
.Y(n_3032)
);

OAI22xp5_ASAP7_75t_L g3033 ( 
.A1(n_2969),
.A2(n_2557),
.B1(n_2891),
.B2(n_2915),
.Y(n_3033)
);

OAI22xp5_ASAP7_75t_L g3034 ( 
.A1(n_2995),
.A2(n_2945),
.B1(n_2728),
.B2(n_2818),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2965),
.B(n_2924),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2965),
.B(n_2968),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2971),
.B(n_2925),
.Y(n_3037)
);

NOR2xp33_ASAP7_75t_L g3038 ( 
.A(n_2957),
.B(n_2820),
.Y(n_3038)
);

AND2x2_ASAP7_75t_L g3039 ( 
.A(n_2967),
.B(n_2953),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_3008),
.B(n_2910),
.Y(n_3040)
);

NOR3xp33_ASAP7_75t_L g3041 ( 
.A(n_2963),
.B(n_2629),
.C(n_2672),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2981),
.B(n_2910),
.Y(n_3042)
);

AND2x2_ASAP7_75t_L g3043 ( 
.A(n_2990),
.B(n_2897),
.Y(n_3043)
);

AND2x2_ASAP7_75t_L g3044 ( 
.A(n_2966),
.B(n_2951),
.Y(n_3044)
);

OA211x2_ASAP7_75t_L g3045 ( 
.A1(n_2973),
.A2(n_2974),
.B(n_2980),
.C(n_2977),
.Y(n_3045)
);

AOI211xp5_ASAP7_75t_L g3046 ( 
.A1(n_2998),
.A2(n_2671),
.B(n_2517),
.C(n_2550),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2994),
.B(n_2853),
.Y(n_3047)
);

AND2x2_ASAP7_75t_L g3048 ( 
.A(n_2956),
.B(n_2853),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_3003),
.B(n_2855),
.Y(n_3049)
);

HB1xp67_ASAP7_75t_L g3050 ( 
.A(n_3031),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_3044),
.B(n_3006),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_L g3052 ( 
.A(n_3047),
.B(n_2952),
.Y(n_3052)
);

AND2x2_ASAP7_75t_L g3053 ( 
.A(n_3039),
.B(n_2964),
.Y(n_3053)
);

AOI21xp33_ASAP7_75t_L g3054 ( 
.A1(n_3011),
.A2(n_2701),
.B(n_2695),
.Y(n_3054)
);

OR2x2_ASAP7_75t_L g3055 ( 
.A(n_3029),
.B(n_3001),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_3043),
.B(n_2975),
.Y(n_3056)
);

HB1xp67_ASAP7_75t_L g3057 ( 
.A(n_3022),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_3049),
.B(n_2959),
.Y(n_3058)
);

AND2x2_ASAP7_75t_L g3059 ( 
.A(n_3019),
.B(n_2988),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_3036),
.B(n_2992),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_3012),
.B(n_3002),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_3035),
.B(n_3004),
.Y(n_3062)
);

AND2x2_ASAP7_75t_L g3063 ( 
.A(n_3021),
.B(n_3005),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_3030),
.Y(n_3064)
);

INVx3_ASAP7_75t_L g3065 ( 
.A(n_3014),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_3048),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_3016),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_3040),
.B(n_2974),
.Y(n_3068)
);

OR2x2_ASAP7_75t_L g3069 ( 
.A(n_3042),
.B(n_2977),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_3037),
.Y(n_3070)
);

HB1xp67_ASAP7_75t_L g3071 ( 
.A(n_3009),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_3045),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_3025),
.Y(n_3073)
);

INVx2_ASAP7_75t_SL g3074 ( 
.A(n_3027),
.Y(n_3074)
);

INVx2_ASAP7_75t_SL g3075 ( 
.A(n_3013),
.Y(n_3075)
);

INVxp67_ASAP7_75t_SL g3076 ( 
.A(n_3023),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_3033),
.Y(n_3077)
);

HB1xp67_ASAP7_75t_L g3078 ( 
.A(n_3017),
.Y(n_3078)
);

HB1xp67_ASAP7_75t_L g3079 ( 
.A(n_3034),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_3015),
.B(n_2938),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_3026),
.Y(n_3081)
);

AND2x2_ASAP7_75t_L g3082 ( 
.A(n_3028),
.B(n_2872),
.Y(n_3082)
);

AND2x2_ASAP7_75t_L g3083 ( 
.A(n_3038),
.B(n_2922),
.Y(n_3083)
);

AND2x4_ASAP7_75t_L g3084 ( 
.A(n_3010),
.B(n_2922),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_3041),
.Y(n_3085)
);

OR2x2_ASAP7_75t_L g3086 ( 
.A(n_3069),
.B(n_2937),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_3050),
.Y(n_3087)
);

INVx2_ASAP7_75t_L g3088 ( 
.A(n_3053),
.Y(n_3088)
);

NOR2xp33_ASAP7_75t_L g3089 ( 
.A(n_3074),
.B(n_3024),
.Y(n_3089)
);

AND2x2_ASAP7_75t_L g3090 ( 
.A(n_3083),
.B(n_3032),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_3085),
.B(n_3018),
.Y(n_3091)
);

INVx2_ASAP7_75t_L g3092 ( 
.A(n_3056),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_3060),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_3062),
.Y(n_3094)
);

OR2x2_ASAP7_75t_L g3095 ( 
.A(n_3068),
.B(n_2912),
.Y(n_3095)
);

AND2x4_ASAP7_75t_L g3096 ( 
.A(n_3065),
.B(n_3032),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_L g3097 ( 
.A(n_3077),
.B(n_3046),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_3062),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_3071),
.B(n_2873),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_3052),
.Y(n_3100)
);

INVx2_ASAP7_75t_SL g3101 ( 
.A(n_3061),
.Y(n_3101)
);

HB1xp67_ASAP7_75t_L g3102 ( 
.A(n_3078),
.Y(n_3102)
);

OAI22xp5_ASAP7_75t_L g3103 ( 
.A1(n_3073),
.A2(n_3020),
.B1(n_2983),
.B2(n_2759),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_3058),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_3094),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_3098),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_3088),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_3093),
.Y(n_3108)
);

OAI21xp5_ASAP7_75t_SL g3109 ( 
.A1(n_3089),
.A2(n_3079),
.B(n_3076),
.Y(n_3109)
);

HB1xp67_ASAP7_75t_L g3110 ( 
.A(n_3102),
.Y(n_3110)
);

AND2x2_ASAP7_75t_L g3111 ( 
.A(n_3096),
.B(n_3072),
.Y(n_3111)
);

AND2x2_ASAP7_75t_L g3112 ( 
.A(n_3090),
.B(n_3081),
.Y(n_3112)
);

NOR2x1_ASAP7_75t_SL g3113 ( 
.A(n_3101),
.B(n_3075),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_3097),
.B(n_3057),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_3087),
.Y(n_3115)
);

INVx2_ASAP7_75t_SL g3116 ( 
.A(n_3092),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_3095),
.Y(n_3117)
);

AOI22xp5_ASAP7_75t_L g3118 ( 
.A1(n_3103),
.A2(n_3084),
.B1(n_3054),
.B2(n_3067),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_3100),
.Y(n_3119)
);

INVxp67_ASAP7_75t_SL g3120 ( 
.A(n_3091),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_3104),
.Y(n_3121)
);

AOI22xp5_ASAP7_75t_L g3122 ( 
.A1(n_3099),
.A2(n_3080),
.B1(n_3064),
.B2(n_3070),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_3086),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_3094),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_3094),
.Y(n_3125)
);

OR2x2_ASAP7_75t_L g3126 ( 
.A(n_3094),
.B(n_3055),
.Y(n_3126)
);

AND2x2_ASAP7_75t_L g3127 ( 
.A(n_3111),
.B(n_3051),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_3120),
.B(n_3082),
.Y(n_3128)
);

AOI21xp5_ASAP7_75t_L g3129 ( 
.A1(n_3113),
.A2(n_3059),
.B(n_3063),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_3110),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_L g3131 ( 
.A(n_3112),
.B(n_3066),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_3126),
.Y(n_3132)
);

INVx1_ASAP7_75t_SL g3133 ( 
.A(n_3114),
.Y(n_3133)
);

INVxp67_ASAP7_75t_L g3134 ( 
.A(n_3118),
.Y(n_3134)
);

INVxp67_ASAP7_75t_SL g3135 ( 
.A(n_3116),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_3117),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_3105),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_3107),
.Y(n_3138)
);

OR2x2_ASAP7_75t_L g3139 ( 
.A(n_3106),
.B(n_2255),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_3108),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_3124),
.Y(n_3141)
);

OR2x2_ASAP7_75t_L g3142 ( 
.A(n_3125),
.B(n_2216),
.Y(n_3142)
);

AND2x2_ASAP7_75t_L g3143 ( 
.A(n_3119),
.B(n_2722),
.Y(n_3143)
);

AND2x2_ASAP7_75t_L g3144 ( 
.A(n_3121),
.B(n_2816),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_3115),
.B(n_2221),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_3123),
.Y(n_3146)
);

NAND2xp33_ASAP7_75t_SL g3147 ( 
.A(n_3122),
.B(n_2816),
.Y(n_3147)
);

AND2x4_ASAP7_75t_L g3148 ( 
.A(n_3113),
.B(n_2709),
.Y(n_3148)
);

NOR3xp33_ASAP7_75t_L g3149 ( 
.A(n_3109),
.B(n_2639),
.C(n_2681),
.Y(n_3149)
);

NOR2xp67_ASAP7_75t_L g3150 ( 
.A(n_3118),
.B(n_637),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_3113),
.Y(n_3151)
);

AND2x2_ASAP7_75t_L g3152 ( 
.A(n_3111),
.B(n_2823),
.Y(n_3152)
);

NOR2xp33_ASAP7_75t_L g3153 ( 
.A(n_3134),
.B(n_637),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_3130),
.Y(n_3154)
);

OAI22xp33_ASAP7_75t_L g3155 ( 
.A1(n_3151),
.A2(n_2896),
.B1(n_2833),
.B2(n_2567),
.Y(n_3155)
);

NOR2xp33_ASAP7_75t_L g3156 ( 
.A(n_3133),
.B(n_638),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_3132),
.Y(n_3157)
);

O2A1O1Ixp33_ASAP7_75t_L g3158 ( 
.A1(n_3135),
.A2(n_2704),
.B(n_2551),
.C(n_2668),
.Y(n_3158)
);

OR2x6_ASAP7_75t_L g3159 ( 
.A(n_3148),
.B(n_2533),
.Y(n_3159)
);

AND2x2_ASAP7_75t_L g3160 ( 
.A(n_3127),
.B(n_2785),
.Y(n_3160)
);

AOI222xp33_ASAP7_75t_L g3161 ( 
.A1(n_3150),
.A2(n_2677),
.B1(n_2636),
.B2(n_2682),
.C1(n_2637),
.C2(n_2699),
.Y(n_3161)
);

AND2x4_ASAP7_75t_L g3162 ( 
.A(n_3148),
.B(n_2703),
.Y(n_3162)
);

AOI221xp5_ASAP7_75t_L g3163 ( 
.A1(n_3136),
.A2(n_2513),
.B1(n_2664),
.B2(n_2498),
.C(n_2535),
.Y(n_3163)
);

AOI21xp5_ASAP7_75t_L g3164 ( 
.A1(n_3128),
.A2(n_3147),
.B(n_3129),
.Y(n_3164)
);

OAI221xp5_ASAP7_75t_L g3165 ( 
.A1(n_3149),
.A2(n_2653),
.B1(n_2661),
.B2(n_2643),
.C(n_2642),
.Y(n_3165)
);

AOI221xp5_ASAP7_75t_L g3166 ( 
.A1(n_3146),
.A2(n_2663),
.B1(n_2203),
.B2(n_2433),
.C(n_2432),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_3154),
.B(n_3137),
.Y(n_3167)
);

CKINVDCx14_ASAP7_75t_R g3168 ( 
.A(n_3156),
.Y(n_3168)
);

INVxp67_ASAP7_75t_L g3169 ( 
.A(n_3157),
.Y(n_3169)
);

NOR2xp33_ASAP7_75t_L g3170 ( 
.A(n_3164),
.B(n_3138),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_3161),
.B(n_3140),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_3162),
.B(n_3141),
.Y(n_3172)
);

AND2x2_ASAP7_75t_L g3173 ( 
.A(n_3159),
.B(n_3152),
.Y(n_3173)
);

NAND2xp33_ASAP7_75t_L g3174 ( 
.A(n_3160),
.B(n_3144),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_3158),
.B(n_3131),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_3159),
.Y(n_3176)
);

BUFx2_ASAP7_75t_L g3177 ( 
.A(n_3155),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_3163),
.B(n_3143),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_3166),
.B(n_3145),
.Y(n_3179)
);

OR2x2_ASAP7_75t_L g3180 ( 
.A(n_3165),
.B(n_3142),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_3153),
.B(n_3139),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_3153),
.B(n_638),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_3153),
.B(n_639),
.Y(n_3183)
);

AOI221xp5_ASAP7_75t_L g3184 ( 
.A1(n_3170),
.A2(n_2436),
.B1(n_2440),
.B2(n_2437),
.C(n_2422),
.Y(n_3184)
);

OAI211xp5_ASAP7_75t_L g3185 ( 
.A1(n_3168),
.A2(n_3171),
.B(n_3169),
.C(n_3175),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_SL g3186 ( 
.A(n_3177),
.B(n_2833),
.Y(n_3186)
);

AOI221xp5_ASAP7_75t_L g3187 ( 
.A1(n_3178),
.A2(n_2442),
.B1(n_2458),
.B2(n_2443),
.C(n_2441),
.Y(n_3187)
);

NOR3xp33_ASAP7_75t_L g3188 ( 
.A(n_3182),
.B(n_2471),
.C(n_2462),
.Y(n_3188)
);

NOR2xp33_ASAP7_75t_SL g3189 ( 
.A(n_3176),
.B(n_2833),
.Y(n_3189)
);

AOI221xp5_ASAP7_75t_L g3190 ( 
.A1(n_3179),
.A2(n_2602),
.B1(n_2597),
.B2(n_2596),
.C(n_2327),
.Y(n_3190)
);

NAND3xp33_ASAP7_75t_L g3191 ( 
.A(n_3183),
.B(n_2184),
.C(n_2403),
.Y(n_3191)
);

AOI221xp5_ASAP7_75t_L g3192 ( 
.A1(n_3167),
.A2(n_2193),
.B1(n_2274),
.B2(n_2268),
.C(n_2931),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_3172),
.Y(n_3193)
);

AOI221xp5_ASAP7_75t_L g3194 ( 
.A1(n_3181),
.A2(n_2935),
.B1(n_2920),
.B2(n_2936),
.C(n_2692),
.Y(n_3194)
);

AOI21xp5_ASAP7_75t_L g3195 ( 
.A1(n_3174),
.A2(n_3180),
.B(n_3173),
.Y(n_3195)
);

AOI221xp5_ASAP7_75t_L g3196 ( 
.A1(n_3170),
.A2(n_2935),
.B1(n_2920),
.B2(n_2936),
.C(n_2679),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_3193),
.Y(n_3197)
);

NAND3xp33_ASAP7_75t_L g3198 ( 
.A(n_3186),
.B(n_2659),
.C(n_2658),
.Y(n_3198)
);

NAND3xp33_ASAP7_75t_SL g3199 ( 
.A(n_3189),
.B(n_643),
.C(n_644),
.Y(n_3199)
);

NAND4xp75_ASAP7_75t_L g3200 ( 
.A(n_3187),
.B(n_3184),
.C(n_3194),
.D(n_3190),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_SL g3201 ( 
.A(n_3196),
.B(n_3188),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3191),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_3192),
.B(n_647),
.Y(n_3203)
);

NAND4xp75_ASAP7_75t_L g3204 ( 
.A(n_3195),
.B(n_652),
.C(n_650),
.D(n_651),
.Y(n_3204)
);

NOR3x1_ASAP7_75t_L g3205 ( 
.A(n_3185),
.B(n_2423),
.C(n_2404),
.Y(n_3205)
);

NOR2x1_ASAP7_75t_L g3206 ( 
.A(n_3204),
.B(n_3197),
.Y(n_3206)
);

NAND4xp25_ASAP7_75t_L g3207 ( 
.A(n_3205),
.B(n_658),
.C(n_656),
.D(n_657),
.Y(n_3207)
);

AOI221xp5_ASAP7_75t_L g3208 ( 
.A1(n_3202),
.A2(n_2705),
.B1(n_661),
.B2(n_659),
.C(n_660),
.Y(n_3208)
);

NOR4xp75_ASAP7_75t_L g3209 ( 
.A(n_3200),
.B(n_3203),
.C(n_3201),
.D(n_3199),
.Y(n_3209)
);

NAND3xp33_ASAP7_75t_SL g3210 ( 
.A(n_3198),
.B(n_663),
.C(n_664),
.Y(n_3210)
);

AND2x4_ASAP7_75t_L g3211 ( 
.A(n_3209),
.B(n_665),
.Y(n_3211)
);

AO22x1_ASAP7_75t_L g3212 ( 
.A1(n_3206),
.A2(n_669),
.B1(n_666),
.B2(n_668),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3210),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3207),
.Y(n_3214)
);

NOR3xp33_ASAP7_75t_L g3215 ( 
.A(n_3208),
.B(n_670),
.C(n_671),
.Y(n_3215)
);

AND2x2_ASAP7_75t_L g3216 ( 
.A(n_3211),
.B(n_674),
.Y(n_3216)
);

AOI21xp5_ASAP7_75t_L g3217 ( 
.A1(n_3212),
.A2(n_674),
.B(n_675),
.Y(n_3217)
);

BUFx4f_ASAP7_75t_SL g3218 ( 
.A(n_3211),
.Y(n_3218)
);

NAND4xp75_ASAP7_75t_L g3219 ( 
.A(n_3214),
.B(n_679),
.C(n_677),
.D(n_678),
.Y(n_3219)
);

NAND3xp33_ASAP7_75t_SL g3220 ( 
.A(n_3215),
.B(n_678),
.C(n_679),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_SL g3221 ( 
.A(n_3218),
.B(n_3213),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3216),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_3219),
.Y(n_3223)
);

AOI22xp5_ASAP7_75t_L g3224 ( 
.A1(n_3220),
.A2(n_2406),
.B1(n_2449),
.B2(n_2364),
.Y(n_3224)
);

OR2x2_ASAP7_75t_L g3225 ( 
.A(n_3217),
.B(n_682),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_3225),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3221),
.Y(n_3227)
);

NOR3xp33_ASAP7_75t_L g3228 ( 
.A(n_3227),
.B(n_3223),
.C(n_3222),
.Y(n_3228)
);

OAI22xp5_ASAP7_75t_SL g3229 ( 
.A1(n_3226),
.A2(n_3224),
.B1(n_685),
.B2(n_683),
.Y(n_3229)
);

AOI21xp5_ASAP7_75t_L g3230 ( 
.A1(n_3229),
.A2(n_686),
.B(n_687),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_3230),
.B(n_3228),
.Y(n_3231)
);

OAI22xp5_ASAP7_75t_L g3232 ( 
.A1(n_3231),
.A2(n_2259),
.B1(n_2321),
.B2(n_2297),
.Y(n_3232)
);

AOI21xp33_ASAP7_75t_SL g3233 ( 
.A1(n_3231),
.A2(n_689),
.B(n_690),
.Y(n_3233)
);

NAND3xp33_ASAP7_75t_SL g3234 ( 
.A(n_3233),
.B(n_691),
.C(n_692),
.Y(n_3234)
);

OAI21xp5_ASAP7_75t_L g3235 ( 
.A1(n_3232),
.A2(n_691),
.B(n_692),
.Y(n_3235)
);

INVx4_ASAP7_75t_L g3236 ( 
.A(n_3234),
.Y(n_3236)
);

AOI221xp5_ASAP7_75t_L g3237 ( 
.A1(n_3236),
.A2(n_3235),
.B1(n_695),
.B2(n_693),
.C(n_694),
.Y(n_3237)
);

AOI211xp5_ASAP7_75t_L g3238 ( 
.A1(n_3237),
.A2(n_700),
.B(n_698),
.C(n_699),
.Y(n_3238)
);


endmodule