module fake_jpeg_11366_n_53 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_53);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_53;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

AND2x2_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_15),
.B1(n_12),
.B2(n_9),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_28),
.B1(n_19),
.B2(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_34),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_26),
.B1(n_29),
.B2(n_22),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_20),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_40),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_20),
.B1(n_23),
.B2(n_30),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_42),
.B1(n_35),
.B2(n_33),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_46),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_32),
.C(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_1),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_38),
.C(n_3),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_45),
.Y(n_50)
);

AO221x1_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_49),
.B1(n_7),
.B2(n_8),
.C(n_18),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_42),
.C(n_3),
.Y(n_52)
);

AOI322xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_30),
.C2(n_43),
.Y(n_53)
);


endmodule