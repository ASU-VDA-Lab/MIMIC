module fake_ariane_2255_n_1419 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_367, n_345, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_221, n_321, n_86, n_361, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_359, n_155, n_127, n_1419);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_359;
input n_155;
input n_127;

output n_1419;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_1295;
wire n_1013;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_965;
wire n_934;
wire n_1220;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1414;
wire n_1134;
wire n_647;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1218;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_608;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_1361;
wire n_1057;
wire n_1011;
wire n_978;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_241),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_143),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_196),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_242),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_285),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_137),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_141),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_24),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_232),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_159),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_35),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_235),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_125),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_13),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_272),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_281),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_110),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_4),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_297),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_361),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_80),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_9),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_129),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_11),
.Y(n_391)
);

INVxp33_ASAP7_75t_SL g392 ( 
.A(n_8),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_79),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_273),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_178),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_158),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_247),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_345),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_210),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_65),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_307),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_123),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_320),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_31),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_315),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_66),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_10),
.Y(n_407)
);

BUFx8_ASAP7_75t_SL g408 ( 
.A(n_108),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_310),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_68),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_190),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_142),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_278),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_202),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_L g415 ( 
.A(n_316),
.B(n_339),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_92),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_305),
.Y(n_417)
);

BUFx10_ASAP7_75t_L g418 ( 
.A(n_77),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_96),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_119),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_189),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_161),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_233),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_211),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_123),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_238),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_146),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_344),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_88),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_186),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_290),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_20),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_87),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_65),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_110),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_306),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_96),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_171),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_127),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_183),
.B(n_145),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_322),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_95),
.Y(n_442)
);

BUFx5_ASAP7_75t_L g443 ( 
.A(n_35),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_93),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_126),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_148),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_100),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_216),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_329),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_46),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_165),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_299),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_269),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_114),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_93),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_282),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_101),
.Y(n_457)
);

BUFx10_ASAP7_75t_L g458 ( 
.A(n_197),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_117),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_135),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_364),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_89),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_139),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_348),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_167),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_304),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_219),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_40),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_203),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_121),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_66),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_337),
.Y(n_472)
);

BUFx10_ASAP7_75t_L g473 ( 
.A(n_116),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_108),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_150),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_38),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_173),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_338),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_151),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_266),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_44),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_217),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_43),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_45),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_200),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_182),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_317),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_51),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_363),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_21),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_L g491 ( 
.A(n_231),
.B(n_357),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_187),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_286),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_34),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_326),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_280),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_207),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_223),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_6),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_79),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_101),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_225),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_82),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_48),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_132),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_204),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_239),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_19),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_292),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_31),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_29),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_58),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_13),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_122),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_57),
.Y(n_515)
);

BUFx2_ASAP7_75t_SL g516 ( 
.A(n_55),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_362),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_122),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_140),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_16),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_358),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_249),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_279),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_212),
.Y(n_524)
);

BUFx10_ASAP7_75t_L g525 ( 
.A(n_7),
.Y(n_525)
);

CKINVDCx14_ASAP7_75t_R g526 ( 
.A(n_170),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_147),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_131),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_149),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_246),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_209),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_111),
.Y(n_532)
);

BUFx10_ASAP7_75t_L g533 ( 
.A(n_26),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_46),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_69),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_59),
.Y(n_536)
);

BUFx10_ASAP7_75t_L g537 ( 
.A(n_97),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_251),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_71),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_342),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_162),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_72),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_152),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_81),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_398),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_398),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_442),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_402),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_442),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_376),
.B(n_0),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_376),
.B(n_0),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_389),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_402),
.A2(n_526),
.B1(n_453),
.B2(n_375),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_389),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_443),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_499),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_398),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_423),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_385),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_432),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_499),
.B(n_4),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_443),
.Y(n_562)
);

OA21x2_ASAP7_75t_L g563 ( 
.A1(n_373),
.A2(n_5),
.B(n_6),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_390),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_430),
.A2(n_8),
.B1(n_5),
.B2(n_7),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_403),
.B(n_9),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_501),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_398),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_443),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_443),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_509),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_515),
.B(n_393),
.Y(n_572)
);

INVx5_ASAP7_75t_L g573 ( 
.A(n_509),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_443),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_464),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_403),
.B(n_12),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_443),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_390),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_509),
.Y(n_579)
);

OA21x2_ASAP7_75t_L g580 ( 
.A1(n_374),
.A2(n_14),
.B(n_15),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_509),
.Y(n_581)
);

BUFx12f_ASAP7_75t_L g582 ( 
.A(n_458),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_494),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_494),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_505),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_368),
.Y(n_586)
);

CKINVDCx6p67_ASAP7_75t_R g587 ( 
.A(n_458),
.Y(n_587)
);

OAI22x1_ASAP7_75t_R g588 ( 
.A1(n_444),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_480),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_384),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_480),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_380),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_505),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_380),
.B(n_17),
.Y(n_594)
);

INVx5_ASAP7_75t_L g595 ( 
.A(n_412),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_388),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_496),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_391),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_505),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_418),
.Y(n_600)
);

OA21x2_ASAP7_75t_L g601 ( 
.A1(n_379),
.A2(n_17),
.B(n_18),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_381),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_377),
.A2(n_138),
.B(n_136),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_R g604 ( 
.A1(n_392),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_465),
.B(n_22),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_506),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_606)
);

CKINVDCx6p67_ASAP7_75t_R g607 ( 
.A(n_418),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_507),
.Y(n_608)
);

OA21x2_ASAP7_75t_L g609 ( 
.A1(n_382),
.A2(n_395),
.B(n_386),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_487),
.B(n_23),
.Y(n_610)
);

INVxp33_ASAP7_75t_SL g611 ( 
.A(n_378),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_526),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_507),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_473),
.B(n_25),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_505),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_396),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_397),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_406),
.Y(n_618)
);

BUFx8_ASAP7_75t_SL g619 ( 
.A(n_408),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_473),
.B(n_27),
.Y(n_620)
);

INVx6_ASAP7_75t_L g621 ( 
.A(n_525),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_399),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_462),
.Y(n_623)
);

AOI22x1_ASAP7_75t_SL g624 ( 
.A1(n_459),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_409),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_416),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_462),
.B(n_28),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_419),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_545),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_552),
.B(n_525),
.Y(n_630)
);

BUFx6f_ASAP7_75t_SL g631 ( 
.A(n_608),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_545),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_568),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_612),
.B(n_560),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_572),
.A2(n_534),
.B1(n_504),
.B2(n_400),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_586),
.B(n_413),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_548),
.B(n_377),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_L g638 ( 
.A(n_576),
.B(n_404),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_548),
.B(n_611),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_545),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_555),
.Y(n_641)
);

AOI21x1_ASAP7_75t_L g642 ( 
.A1(n_555),
.A2(n_387),
.B(n_383),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_562),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_545),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_562),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_568),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_569),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_546),
.Y(n_648)
);

AND3x2_ASAP7_75t_L g649 ( 
.A(n_547),
.B(n_387),
.C(n_383),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_546),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_546),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_616),
.B(n_417),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_557),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_557),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_621),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_557),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_573),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_571),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_611),
.B(n_414),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_585),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_586),
.B(n_531),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_587),
.Y(n_662)
);

AOI21x1_ASAP7_75t_L g663 ( 
.A1(n_570),
.A2(n_427),
.B(n_414),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_579),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_570),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_621),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_579),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_553),
.B(n_427),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_579),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_581),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_574),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_581),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_621),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_574),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_585),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_661),
.B(n_595),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_630),
.B(n_655),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_637),
.B(n_582),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_630),
.B(n_636),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_659),
.B(n_582),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_641),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_635),
.A2(n_551),
.B1(n_566),
.B2(n_550),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_655),
.B(n_605),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_666),
.B(n_610),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_641),
.B(n_643),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_666),
.B(n_610),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_673),
.B(n_639),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_673),
.B(n_600),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_645),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_668),
.B(n_608),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_647),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_665),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_671),
.B(n_674),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_671),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_635),
.B(n_620),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_638),
.B(n_607),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_662),
.B(n_614),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_652),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_652),
.A2(n_609),
.B(n_577),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_629),
.A2(n_609),
.B(n_577),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_634),
.A2(n_561),
.B1(n_584),
.B2(n_583),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_662),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_SL g703 ( 
.A(n_631),
.B(n_619),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_660),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_660),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_649),
.B(n_567),
.Y(n_706)
);

INVx8_ASAP7_75t_L g707 ( 
.A(n_631),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_675),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_648),
.Y(n_709)
);

NAND2xp33_ASAP7_75t_L g710 ( 
.A(n_648),
.B(n_369),
.Y(n_710)
);

AND2x6_ASAP7_75t_SL g711 ( 
.A(n_634),
.B(n_604),
.Y(n_711)
);

NAND2xp33_ASAP7_75t_L g712 ( 
.A(n_648),
.B(n_370),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_642),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_634),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_642),
.Y(n_715)
);

INVx8_ASAP7_75t_L g716 ( 
.A(n_634),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_629),
.B(n_589),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_646),
.B(n_549),
.Y(n_718)
);

AOI221xp5_ASAP7_75t_L g719 ( 
.A1(n_634),
.A2(n_556),
.B1(n_547),
.B2(n_627),
.C(n_565),
.Y(n_719)
);

NOR2x2_ASAP7_75t_L g720 ( 
.A(n_632),
.B(n_588),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_640),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_663),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_640),
.B(n_589),
.Y(n_723)
);

OAI22xp33_ASAP7_75t_L g724 ( 
.A1(n_663),
.A2(n_575),
.B1(n_606),
.B2(n_558),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_644),
.B(n_556),
.C(n_594),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_644),
.B(n_591),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_650),
.B(n_591),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_650),
.B(n_592),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_646),
.B(n_554),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_651),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_648),
.B(n_627),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_653),
.B(n_591),
.Y(n_732)
);

OAI22xp33_ASAP7_75t_SL g733 ( 
.A1(n_654),
.A2(n_433),
.B1(n_407),
.B2(n_410),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_646),
.B(n_564),
.Y(n_734)
);

OAI21xp33_ASAP7_75t_L g735 ( 
.A1(n_658),
.A2(n_596),
.B(n_590),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_698),
.B(n_616),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_681),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_685),
.A2(n_603),
.B(n_609),
.Y(n_738)
);

INVx1_ASAP7_75t_SL g739 ( 
.A(n_702),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_714),
.B(n_592),
.Y(n_740)
);

AND2x2_ASAP7_75t_SL g741 ( 
.A(n_703),
.B(n_563),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_693),
.A2(n_646),
.B(n_633),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_714),
.B(n_701),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_719),
.A2(n_696),
.B(n_699),
.C(n_691),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_704),
.Y(n_745)
);

O2A1O1Ixp5_ASAP7_75t_L g746 ( 
.A1(n_684),
.A2(n_449),
.B(n_451),
.C(n_438),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_707),
.Y(n_747)
);

A2O1A1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_719),
.A2(n_425),
.B(n_429),
.C(n_420),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_L g749 ( 
.A1(n_700),
.A2(n_699),
.B(n_713),
.Y(n_749)
);

INVx5_ASAP7_75t_L g750 ( 
.A(n_707),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_695),
.A2(n_622),
.B1(n_625),
.B2(n_617),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_690),
.B(n_617),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_692),
.A2(n_694),
.B(n_683),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_676),
.A2(n_657),
.B(n_580),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_724),
.A2(n_625),
.B1(n_622),
.B2(n_580),
.Y(n_755)
);

OAI22x1_ASAP7_75t_L g756 ( 
.A1(n_711),
.A2(n_559),
.B1(n_624),
.B2(n_623),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_L g757 ( 
.A1(n_700),
.A2(n_722),
.B(n_715),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_689),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_728),
.Y(n_759)
);

AO22x1_ASAP7_75t_L g760 ( 
.A1(n_680),
.A2(n_623),
.B1(n_602),
.B2(n_445),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_686),
.A2(n_657),
.B(n_601),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_706),
.B(n_602),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_707),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_718),
.B(n_435),
.Y(n_764)
);

OAI21xp5_ASAP7_75t_L g765 ( 
.A1(n_705),
.A2(n_460),
.B(n_452),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_678),
.B(n_559),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_677),
.B(n_578),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_716),
.A2(n_447),
.B1(n_455),
.B2(n_450),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_687),
.A2(n_470),
.B1(n_471),
.B2(n_457),
.Y(n_769)
);

BUFx12f_ASAP7_75t_L g770 ( 
.A(n_709),
.Y(n_770)
);

BUFx4f_ASAP7_75t_L g771 ( 
.A(n_716),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_708),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_729),
.A2(n_434),
.B(n_439),
.C(n_437),
.Y(n_773)
);

A2O1A1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_734),
.A2(n_468),
.B(n_474),
.C(n_454),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_716),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_731),
.B(n_597),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_697),
.B(n_619),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_709),
.Y(n_778)
);

OAI21xp33_ASAP7_75t_L g779 ( 
.A1(n_725),
.A2(n_488),
.B(n_483),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_709),
.Y(n_780)
);

O2A1O1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_733),
.A2(n_481),
.B(n_484),
.C(n_476),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_717),
.A2(n_667),
.B(n_664),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_688),
.B(n_598),
.Y(n_783)
);

NOR3xp33_ASAP7_75t_L g784 ( 
.A(n_735),
.B(n_503),
.C(n_490),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_721),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_723),
.A2(n_669),
.B(n_667),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_726),
.A2(n_670),
.B(n_669),
.Y(n_787)
);

AO22x1_ASAP7_75t_L g788 ( 
.A1(n_720),
.A2(n_500),
.B1(n_514),
.B2(n_510),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_730),
.A2(n_463),
.B(n_461),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_727),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_SL g791 ( 
.A(n_732),
.B(n_533),
.Y(n_791)
);

A2O1A1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_710),
.A2(n_511),
.B(n_512),
.C(n_508),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_R g793 ( 
.A(n_712),
.B(n_372),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_698),
.B(n_613),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_698),
.B(n_613),
.Y(n_795)
);

O2A1O1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_682),
.A2(n_518),
.B(n_528),
.C(n_513),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_698),
.A2(n_672),
.B(n_475),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_698),
.B(n_613),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_698),
.B(n_371),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_698),
.A2(n_477),
.B(n_472),
.Y(n_800)
);

OAI21xp33_ASAP7_75t_L g801 ( 
.A1(n_682),
.A2(n_536),
.B(n_520),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_704),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_698),
.A2(n_479),
.B(n_478),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_698),
.A2(n_489),
.B(n_485),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_698),
.A2(n_497),
.B(n_492),
.Y(n_805)
);

AO32x1_ASAP7_75t_L g806 ( 
.A1(n_682),
.A2(n_593),
.A3(n_428),
.B1(n_431),
.B2(n_495),
.Y(n_806)
);

O2A1O1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_682),
.A2(n_535),
.B(n_532),
.C(n_618),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_679),
.A2(n_539),
.B1(n_544),
.B2(n_542),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_714),
.Y(n_809)
);

O2A1O1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_682),
.A2(n_626),
.B(n_628),
.C(n_593),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_728),
.B(n_599),
.Y(n_811)
);

AOI21x1_ASAP7_75t_L g812 ( 
.A1(n_700),
.A2(n_491),
.B(n_415),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_704),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_698),
.A2(n_519),
.B(n_524),
.C(n_521),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_679),
.A2(n_516),
.B1(n_529),
.B2(n_527),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_698),
.A2(n_530),
.B(n_440),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_704),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_679),
.B(n_533),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_698),
.B(n_394),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_L g820 ( 
.A1(n_700),
.A2(n_446),
.B(n_431),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_682),
.A2(n_537),
.B1(n_495),
.B2(n_498),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_702),
.B(n_537),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_679),
.B(n_401),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_704),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_700),
.A2(n_411),
.B(n_405),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_775),
.B(n_599),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_757),
.A2(n_422),
.B(n_421),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_743),
.B(n_615),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_770),
.Y(n_829)
);

AOI21x1_ASAP7_75t_L g830 ( 
.A1(n_812),
.A2(n_573),
.B(n_656),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_744),
.A2(n_426),
.B1(n_436),
.B2(n_424),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_747),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_825),
.A2(n_448),
.B(n_441),
.Y(n_833)
);

AO31x2_ASAP7_75t_L g834 ( 
.A1(n_738),
.A2(n_814),
.A3(n_754),
.B(n_761),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_737),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_762),
.B(n_30),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_740),
.B(n_32),
.Y(n_837)
);

O2A1O1Ixp5_ASAP7_75t_L g838 ( 
.A1(n_816),
.A2(n_36),
.B(n_33),
.C(n_34),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_753),
.A2(n_466),
.B(n_456),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_799),
.B(n_467),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_739),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_SL g842 ( 
.A(n_766),
.B(n_469),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_771),
.B(n_482),
.Y(n_843)
);

NOR2xp67_ASAP7_75t_SL g844 ( 
.A(n_750),
.B(n_486),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_742),
.A2(n_502),
.B(n_493),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_818),
.B(n_517),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_736),
.B(n_522),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_772),
.Y(n_848)
);

NOR2x1_ASAP7_75t_SL g849 ( 
.A(n_750),
.B(n_656),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_771),
.B(n_523),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_809),
.B(n_33),
.Y(n_851)
);

A2O1A1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_796),
.A2(n_540),
.B(n_541),
.C(n_538),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_821),
.A2(n_543),
.B1(n_38),
.B2(n_36),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_SL g854 ( 
.A1(n_768),
.A2(n_40),
.B1(n_37),
.B2(n_39),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_764),
.A2(n_41),
.B1(n_37),
.B2(n_39),
.Y(n_855)
);

NOR2x1_ASAP7_75t_SL g856 ( 
.A(n_778),
.B(n_656),
.Y(n_856)
);

OAI21xp33_ASAP7_75t_L g857 ( 
.A1(n_801),
.A2(n_41),
.B(n_42),
.Y(n_857)
);

INVx4_ASAP7_75t_SL g858 ( 
.A(n_822),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_794),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_859)
);

OAI21x1_ASAP7_75t_SL g860 ( 
.A1(n_807),
.A2(n_45),
.B(n_47),
.Y(n_860)
);

AO21x1_ASAP7_75t_L g861 ( 
.A1(n_820),
.A2(n_581),
.B(n_144),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_778),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_768),
.B(n_47),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_795),
.A2(n_52),
.B1(n_49),
.B2(n_50),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_745),
.B(n_50),
.Y(n_865)
);

CKINVDCx16_ASAP7_75t_R g866 ( 
.A(n_777),
.Y(n_866)
);

NAND2x1p5_ASAP7_75t_L g867 ( 
.A(n_745),
.B(n_52),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_811),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_760),
.B(n_53),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_758),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_811),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_752),
.B(n_53),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_759),
.B(n_54),
.Y(n_873)
);

AOI221x1_ASAP7_75t_L g874 ( 
.A1(n_789),
.A2(n_57),
.B1(n_54),
.B2(n_56),
.C(n_58),
.Y(n_874)
);

INVx1_ASAP7_75t_SL g875 ( 
.A(n_763),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_815),
.A2(n_60),
.B1(n_56),
.B2(n_59),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_808),
.B(n_60),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_798),
.Y(n_878)
);

BUFx8_ASAP7_75t_L g879 ( 
.A(n_783),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_778),
.Y(n_880)
);

AO31x2_ASAP7_75t_L g881 ( 
.A1(n_790),
.A2(n_63),
.A3(n_61),
.B(n_62),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_797),
.A2(n_154),
.B(n_153),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_L g883 ( 
.A(n_780),
.B(n_61),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_755),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_813),
.B(n_64),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_788),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_765),
.A2(n_70),
.B(n_67),
.C(n_68),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_800),
.A2(n_71),
.B(n_67),
.C(n_70),
.Y(n_888)
);

OAI21x1_ASAP7_75t_L g889 ( 
.A1(n_782),
.A2(n_787),
.B(n_786),
.Y(n_889)
);

NAND2x1_ASAP7_75t_L g890 ( 
.A(n_780),
.B(n_155),
.Y(n_890)
);

OAI21x1_ASAP7_75t_SL g891 ( 
.A1(n_803),
.A2(n_72),
.B(n_73),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_813),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_804),
.A2(n_157),
.B(n_156),
.Y(n_893)
);

AO31x2_ASAP7_75t_L g894 ( 
.A1(n_806),
.A2(n_773),
.A3(n_774),
.B(n_805),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_SL g895 ( 
.A1(n_756),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_748),
.A2(n_76),
.B(n_74),
.C(n_75),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_802),
.Y(n_897)
);

INVx6_ASAP7_75t_SL g898 ( 
.A(n_791),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_767),
.B(n_76),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_817),
.A2(n_824),
.B(n_776),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_779),
.B(n_77),
.Y(n_901)
);

INVxp67_ASAP7_75t_SL g902 ( 
.A(n_780),
.Y(n_902)
);

OAI21x1_ASAP7_75t_L g903 ( 
.A1(n_810),
.A2(n_163),
.B(n_160),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_785),
.B(n_78),
.Y(n_904)
);

AO31x2_ASAP7_75t_L g905 ( 
.A1(n_806),
.A2(n_81),
.A3(n_78),
.B(n_80),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_751),
.B(n_82),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_741),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_793),
.B(n_83),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_746),
.A2(n_166),
.B(n_164),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_792),
.A2(n_169),
.B(n_168),
.Y(n_910)
);

AOI211x1_ASAP7_75t_L g911 ( 
.A1(n_769),
.A2(n_86),
.B(n_84),
.C(n_85),
.Y(n_911)
);

AO31x2_ASAP7_75t_L g912 ( 
.A1(n_806),
.A2(n_87),
.A3(n_85),
.B(n_86),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_784),
.B(n_88),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_781),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_823),
.B(n_89),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_747),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_762),
.B(n_90),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_823),
.B(n_91),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_744),
.A2(n_97),
.B1(n_94),
.B2(n_95),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_823),
.B(n_94),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_825),
.A2(n_174),
.B(n_172),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_757),
.A2(n_176),
.B(n_175),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_823),
.B(n_98),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_744),
.A2(n_100),
.B(n_98),
.C(n_99),
.Y(n_924)
);

NAND2x1p5_ASAP7_75t_L g925 ( 
.A(n_775),
.B(n_99),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_766),
.B(n_102),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_744),
.A2(n_104),
.B(n_102),
.C(n_103),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_737),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_770),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_825),
.A2(n_179),
.B(n_177),
.Y(n_930)
);

NAND3xp33_ASAP7_75t_L g931 ( 
.A(n_823),
.B(n_104),
.C(n_105),
.Y(n_931)
);

OA22x2_ASAP7_75t_L g932 ( 
.A1(n_768),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_825),
.A2(n_181),
.B(n_180),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_823),
.B(n_106),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_825),
.A2(n_185),
.B(n_184),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_823),
.B(n_107),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_744),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_750),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_823),
.B(n_109),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_SL g940 ( 
.A1(n_766),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_940)
);

NAND2x1p5_ASAP7_75t_L g941 ( 
.A(n_775),
.B(n_113),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_762),
.B(n_115),
.Y(n_942)
);

OA21x2_ASAP7_75t_L g943 ( 
.A1(n_749),
.A2(n_191),
.B(n_188),
.Y(n_943)
);

AOI221x1_ASAP7_75t_L g944 ( 
.A1(n_744),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.C(n_118),
.Y(n_944)
);

OAI21x1_ASAP7_75t_SL g945 ( 
.A1(n_816),
.A2(n_118),
.B(n_120),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_825),
.A2(n_193),
.B(n_192),
.Y(n_946)
);

AO21x1_ASAP7_75t_L g947 ( 
.A1(n_820),
.A2(n_195),
.B(n_194),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_762),
.B(n_120),
.Y(n_948)
);

AOI21x1_ASAP7_75t_SL g949 ( 
.A1(n_819),
.A2(n_121),
.B(n_124),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_823),
.B(n_124),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_825),
.A2(n_199),
.B(n_198),
.Y(n_951)
);

AO21x1_ASAP7_75t_L g952 ( 
.A1(n_820),
.A2(n_367),
.B(n_201),
.Y(n_952)
);

O2A1O1Ixp5_ASAP7_75t_L g953 ( 
.A1(n_825),
.A2(n_125),
.B(n_126),
.C(n_127),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_744),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_823),
.B(n_128),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_823),
.B(n_130),
.Y(n_956)
);

NAND3xp33_ASAP7_75t_L g957 ( 
.A(n_823),
.B(n_131),
.C(n_132),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_739),
.B(n_133),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_770),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_747),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_757),
.A2(n_206),
.B(n_205),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_762),
.B(n_133),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_737),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_775),
.B(n_134),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_823),
.B(n_208),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_809),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_966),
.Y(n_967)
);

AO21x2_ASAP7_75t_L g968 ( 
.A1(n_921),
.A2(n_213),
.B(n_214),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_842),
.B(n_215),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_828),
.B(n_218),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_959),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_835),
.Y(n_972)
);

NOR2xp67_ASAP7_75t_L g973 ( 
.A(n_880),
.B(n_220),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_928),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_963),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_930),
.A2(n_221),
.B(n_222),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_870),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_926),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_978)
);

BUFx2_ASAP7_75t_R g979 ( 
.A(n_886),
.Y(n_979)
);

AO31x2_ASAP7_75t_L g980 ( 
.A1(n_861),
.A2(n_228),
.A3(n_229),
.B(n_230),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_929),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_915),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_982)
);

AO31x2_ASAP7_75t_L g983 ( 
.A1(n_947),
.A2(n_240),
.A3(n_243),
.B(n_244),
.Y(n_983)
);

INVxp67_ASAP7_75t_SL g984 ( 
.A(n_907),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_858),
.B(n_245),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_935),
.A2(n_248),
.B(n_250),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_836),
.B(n_366),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_940),
.A2(n_901),
.B1(n_854),
.B2(n_863),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_866),
.B(n_252),
.Y(n_989)
);

AO21x2_ASAP7_75t_L g990 ( 
.A1(n_946),
.A2(n_253),
.B(n_254),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_929),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_868),
.Y(n_992)
);

AO31x2_ASAP7_75t_L g993 ( 
.A1(n_952),
.A2(n_255),
.A3(n_256),
.B(n_257),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_951),
.A2(n_258),
.B(n_259),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_953),
.A2(n_260),
.B(n_261),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_916),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_853),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_848),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_873),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_965),
.A2(n_265),
.B(n_267),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_846),
.B(n_268),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_885),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_917),
.B(n_270),
.Y(n_1003)
);

AO31x2_ASAP7_75t_L g1004 ( 
.A1(n_944),
.A2(n_271),
.A3(n_274),
.B(n_275),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_885),
.Y(n_1005)
);

NOR2x1_ASAP7_75t_SL g1006 ( 
.A(n_938),
.B(n_276),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_875),
.B(n_277),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_897),
.Y(n_1008)
);

NAND3xp33_ASAP7_75t_L g1009 ( 
.A(n_920),
.B(n_283),
.C(n_284),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_862),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_914),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_857),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_1012)
);

OAI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_877),
.A2(n_365),
.B1(n_291),
.B2(n_293),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_878),
.B(n_294),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_913),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_858),
.B(n_295),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_872),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_923),
.A2(n_296),
.B(n_298),
.C(n_300),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_899),
.B(n_301),
.Y(n_1019)
);

BUFx4f_ASAP7_75t_SL g1020 ( 
.A(n_960),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_929),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_832),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_837),
.B(n_302),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_829),
.B(n_303),
.Y(n_1024)
);

INVx2_ASAP7_75t_SL g1025 ( 
.A(n_879),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_892),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_862),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_829),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_906),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_867),
.Y(n_1030)
);

AOI21x1_ASAP7_75t_L g1031 ( 
.A1(n_934),
.A2(n_308),
.B(n_309),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_879),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_871),
.B(n_314),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_851),
.B(n_318),
.Y(n_1034)
);

NAND3xp33_ASAP7_75t_L g1035 ( 
.A(n_936),
.B(n_319),
.C(n_321),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_964),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_898),
.Y(n_1037)
);

AOI221xp5_ASAP7_75t_L g1038 ( 
.A1(n_884),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.C(n_327),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_826),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_964),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_840),
.B(n_328),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_826),
.B(n_330),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_942),
.B(n_331),
.Y(n_1043)
);

OR2x6_ASAP7_75t_L g1044 ( 
.A(n_938),
.B(n_332),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_925),
.Y(n_1045)
);

AOI22x1_ASAP7_75t_L g1046 ( 
.A1(n_833),
.A2(n_827),
.B1(n_961),
.B2(n_922),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_945),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_948),
.B(n_360),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_962),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_1049)
);

AOI31xp67_ASAP7_75t_L g1050 ( 
.A1(n_939),
.A2(n_336),
.A3(n_340),
.B(n_341),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_R g1051 ( 
.A(n_880),
.B(n_343),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_950),
.B(n_346),
.Y(n_1052)
);

BUFx8_ASAP7_75t_L g1053 ( 
.A(n_862),
.Y(n_1053)
);

INVx3_ASAP7_75t_SL g1054 ( 
.A(n_958),
.Y(n_1054)
);

AO21x2_ASAP7_75t_L g1055 ( 
.A1(n_882),
.A2(n_347),
.B(n_349),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_SL g1056 ( 
.A1(n_895),
.A2(n_869),
.B1(n_932),
.B2(n_956),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_849),
.B(n_350),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_955),
.A2(n_351),
.B(n_352),
.Y(n_1058)
);

OAI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_876),
.A2(n_359),
.B1(n_354),
.B2(n_355),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_865),
.Y(n_1060)
);

OR3x4_ASAP7_75t_SL g1061 ( 
.A(n_898),
.B(n_353),
.C(n_356),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_908),
.A2(n_855),
.B1(n_831),
.B2(n_931),
.Y(n_1062)
);

CKINVDCx6p67_ASAP7_75t_R g1063 ( 
.A(n_843),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_904),
.B(n_941),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_957),
.A2(n_937),
.B1(n_954),
.B2(n_919),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_900),
.B(n_847),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_924),
.A2(n_927),
.B(n_903),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_860),
.A2(n_910),
.B1(n_864),
.B2(n_859),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_883),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_891),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_838),
.A2(n_909),
.B(n_852),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_850),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_896),
.B(n_887),
.Y(n_1073)
);

AO21x2_ASAP7_75t_L g1074 ( 
.A1(n_893),
.A2(n_845),
.B(n_856),
.Y(n_1074)
);

NAND2x1p5_ASAP7_75t_L g1075 ( 
.A(n_844),
.B(n_890),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_888),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_881),
.B(n_894),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_902),
.A2(n_943),
.B1(n_839),
.B2(n_874),
.Y(n_1078)
);

CKINVDCx16_ASAP7_75t_R g1079 ( 
.A(n_911),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_949),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_SL g1081 ( 
.A1(n_856),
.A2(n_834),
.B(n_905),
.C(n_912),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_889),
.A2(n_749),
.B(n_830),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_842),
.B(n_766),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_889),
.A2(n_749),
.B(n_830),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_889),
.A2(n_749),
.B(n_830),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_835),
.Y(n_1086)
);

AO21x2_ASAP7_75t_L g1087 ( 
.A1(n_921),
.A2(n_933),
.B(n_930),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_926),
.A2(n_766),
.B1(n_719),
.B2(n_743),
.Y(n_1088)
);

AO21x2_ASAP7_75t_L g1089 ( 
.A1(n_921),
.A2(n_933),
.B(n_930),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_842),
.B(n_841),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_926),
.A2(n_915),
.B1(n_920),
.B2(n_918),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_835),
.Y(n_1092)
);

NOR2x1_ASAP7_75t_SL g1093 ( 
.A(n_938),
.B(n_770),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_835),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_835),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_926),
.A2(n_766),
.B1(n_719),
.B2(n_743),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_L g1097 ( 
.A(n_926),
.B(n_842),
.C(n_915),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_SL g1098 ( 
.A1(n_842),
.A2(n_766),
.B1(n_559),
.B2(n_926),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_836),
.B(n_714),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_959),
.B(n_775),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_972),
.Y(n_1101)
);

OR2x2_ASAP7_75t_L g1102 ( 
.A(n_967),
.B(n_1088),
.Y(n_1102)
);

OA21x2_ASAP7_75t_L g1103 ( 
.A1(n_1082),
.A2(n_1085),
.B(n_1084),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1011),
.B(n_1017),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_1053),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_974),
.Y(n_1106)
);

OAI21xp33_ASAP7_75t_SL g1107 ( 
.A1(n_976),
.A2(n_994),
.B(n_986),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_1096),
.B(n_1036),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_975),
.Y(n_1109)
);

INVx6_ASAP7_75t_L g1110 ( 
.A(n_1053),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1086),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1092),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1094),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1091),
.A2(n_1097),
.B(n_1083),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1095),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_1022),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_992),
.B(n_1040),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_971),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1098),
.B(n_1099),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1056),
.B(n_984),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_977),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_998),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1002),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1005),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1008),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1015),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1042),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_985),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_1100),
.Y(n_1129)
);

BUFx2_ASAP7_75t_SL g1130 ( 
.A(n_996),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1091),
.A2(n_1097),
.B(n_1065),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_1100),
.Y(n_1132)
);

OR2x6_ASAP7_75t_L g1133 ( 
.A(n_985),
.B(n_1016),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1026),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1010),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1039),
.B(n_979),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_999),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1060),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1029),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_1090),
.B(n_1064),
.Y(n_1140)
);

INVx8_ASAP7_75t_L g1141 ( 
.A(n_1044),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_988),
.A2(n_1073),
.B1(n_1076),
.B2(n_1079),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1030),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_970),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1010),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1027),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1027),
.Y(n_1147)
);

INVxp67_ASAP7_75t_L g1148 ( 
.A(n_1033),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1047),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1054),
.B(n_989),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1044),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1044),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_988),
.A2(n_1062),
.B1(n_1087),
.B2(n_1089),
.Y(n_1153)
);

AO21x2_ASAP7_75t_L g1154 ( 
.A1(n_1087),
.A2(n_1089),
.B(n_1081),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1020),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1093),
.B(n_1045),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1070),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1025),
.B(n_1037),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_987),
.A2(n_1003),
.B1(n_1048),
.B2(n_1068),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1069),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1014),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1072),
.A2(n_1063),
.B1(n_1001),
.B2(n_997),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1028),
.B(n_991),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1014),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_973),
.B(n_1057),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1034),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_1021),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1077),
.Y(n_1168)
);

BUFx2_ASAP7_75t_SL g1169 ( 
.A(n_981),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1080),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_969),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1051),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1007),
.B(n_1023),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1051),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1066),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1023),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_1067),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1066),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1019),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1067),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1032),
.B(n_1043),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_973),
.Y(n_1182)
);

CKINVDCx16_ASAP7_75t_R g1183 ( 
.A(n_1061),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1052),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1024),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1006),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1041),
.B(n_1004),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1050),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1075),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1078),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1031),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_997),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1078),
.B(n_1074),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1004),
.B(n_1049),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1071),
.B(n_1013),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1071),
.B(n_1035),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_1018),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1004),
.Y(n_1198)
);

INVxp67_ASAP7_75t_L g1199 ( 
.A(n_1012),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_982),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_986),
.A2(n_978),
.B1(n_1046),
.B2(n_1038),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_982),
.Y(n_1202)
);

AO21x2_ASAP7_75t_L g1203 ( 
.A1(n_995),
.A2(n_968),
.B(n_990),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1009),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1035),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1173),
.B(n_1059),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1101),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1142),
.B(n_1153),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1106),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1109),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1133),
.B(n_993),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1111),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1153),
.B(n_993),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1118),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1131),
.B(n_983),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1118),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_1130),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1112),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1114),
.B(n_968),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1163),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1104),
.B(n_1148),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1168),
.B(n_983),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1113),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1104),
.B(n_1058),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1148),
.B(n_1000),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1102),
.B(n_980),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1115),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1121),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_1108),
.B(n_1055),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1177),
.B(n_990),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1117),
.B(n_1140),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1177),
.B(n_1180),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1180),
.B(n_1192),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1137),
.B(n_1179),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1190),
.B(n_1139),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1176),
.B(n_1126),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1122),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1187),
.B(n_1175),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1120),
.B(n_1119),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_1167),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1183),
.B(n_1150),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1138),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1134),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1162),
.B(n_1127),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1128),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1123),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1124),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_1143),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1178),
.B(n_1149),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1166),
.B(n_1129),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1157),
.B(n_1160),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1184),
.B(n_1200),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1202),
.B(n_1159),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1159),
.B(n_1144),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1132),
.B(n_1172),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1110),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1199),
.A2(n_1181),
.B1(n_1107),
.B2(n_1195),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1125),
.Y(n_1258)
);

AND2x2_ASAP7_75t_SL g1259 ( 
.A(n_1195),
.B(n_1196),
.Y(n_1259)
);

BUFx12f_ASAP7_75t_L g1260 ( 
.A(n_1110),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1152),
.B(n_1161),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1145),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1174),
.B(n_1141),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1141),
.B(n_1171),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_1110),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1164),
.B(n_1151),
.Y(n_1266)
);

AND2x2_ASAP7_75t_SL g1267 ( 
.A(n_1196),
.B(n_1194),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1136),
.B(n_1116),
.Y(n_1268)
);

NOR2x1_ASAP7_75t_L g1269 ( 
.A(n_1170),
.B(n_1189),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1197),
.A2(n_1201),
.B1(n_1203),
.B2(n_1165),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1189),
.B(n_1105),
.Y(n_1271)
);

NAND2x1_ASAP7_75t_L g1272 ( 
.A(n_1186),
.B(n_1182),
.Y(n_1272)
);

INVx4_ASAP7_75t_L g1273 ( 
.A(n_1245),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1232),
.B(n_1198),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1232),
.B(n_1198),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1221),
.B(n_1116),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1243),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1258),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1242),
.Y(n_1279)
);

INVxp67_ASAP7_75t_L g1280 ( 
.A(n_1231),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1261),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1233),
.B(n_1193),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1235),
.B(n_1193),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1251),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1251),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1267),
.B(n_1154),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1207),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1214),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1234),
.B(n_1135),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1238),
.B(n_1253),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1209),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1257),
.A2(n_1201),
.B(n_1204),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1234),
.B(n_1135),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1210),
.Y(n_1294)
);

INVx1_ASAP7_75t_SL g1295 ( 
.A(n_1214),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1261),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1216),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1212),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1236),
.B(n_1146),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1218),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1223),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1227),
.Y(n_1302)
);

NOR2x1p5_ASAP7_75t_L g1303 ( 
.A(n_1260),
.B(n_1105),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1216),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1236),
.B(n_1147),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1211),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1266),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1228),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1237),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1249),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1235),
.B(n_1103),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1252),
.B(n_1103),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1249),
.B(n_1103),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_SL g1314 ( 
.A(n_1260),
.B(n_1155),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1213),
.B(n_1205),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1281),
.B(n_1226),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1296),
.B(n_1259),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1290),
.B(n_1248),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1277),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1278),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1292),
.A2(n_1257),
.B(n_1219),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1315),
.B(n_1230),
.Y(n_1322)
);

NOR2xp67_ASAP7_75t_L g1323 ( 
.A(n_1311),
.B(n_1265),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1284),
.B(n_1259),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1279),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1315),
.B(n_1230),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1287),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1291),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_SL g1329 ( 
.A1(n_1286),
.A2(n_1219),
.B(n_1270),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1313),
.B(n_1213),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1294),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1298),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1313),
.B(n_1215),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1300),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1290),
.B(n_1215),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1283),
.B(n_1254),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1295),
.B(n_1240),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1301),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1312),
.B(n_1222),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1285),
.B(n_1254),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1307),
.B(n_1268),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1302),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1311),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1280),
.B(n_1266),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1283),
.B(n_1229),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1288),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1276),
.B(n_1246),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1325),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1327),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1328),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1347),
.B(n_1312),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1343),
.B(n_1282),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1333),
.B(n_1306),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1331),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1343),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1335),
.B(n_1304),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1343),
.B(n_1282),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1333),
.B(n_1274),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1330),
.B(n_1274),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1330),
.B(n_1275),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1332),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1337),
.B(n_1217),
.Y(n_1362)
);

AOI33xp33_ASAP7_75t_L g1363 ( 
.A1(n_1319),
.A2(n_1308),
.A3(n_1309),
.B1(n_1208),
.B2(n_1158),
.B3(n_1310),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1334),
.Y(n_1364)
);

INVxp67_ASAP7_75t_L g1365 ( 
.A(n_1337),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1339),
.B(n_1286),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1318),
.B(n_1314),
.Y(n_1367)
);

NAND2x1_ASAP7_75t_L g1368 ( 
.A(n_1346),
.B(n_1273),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1338),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1355),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1353),
.B(n_1341),
.Y(n_1371)
);

XOR2x2_ASAP7_75t_L g1372 ( 
.A(n_1362),
.B(n_1241),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1365),
.B(n_1367),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1348),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1363),
.A2(n_1321),
.B(n_1329),
.Y(n_1375)
);

O2A1O1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1363),
.A2(n_1206),
.B(n_1244),
.C(n_1225),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1352),
.B(n_1335),
.Y(n_1377)
);

AOI21xp33_ASAP7_75t_L g1378 ( 
.A1(n_1349),
.A2(n_1269),
.B(n_1320),
.Y(n_1378)
);

INVxp67_ASAP7_75t_L g1379 ( 
.A(n_1356),
.Y(n_1379)
);

AOI221xp5_ASAP7_75t_L g1380 ( 
.A1(n_1350),
.A2(n_1239),
.B1(n_1342),
.B2(n_1326),
.C(n_1322),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1354),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1358),
.B(n_1322),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1358),
.B(n_1326),
.Y(n_1383)
);

AOI21xp33_ASAP7_75t_L g1384 ( 
.A1(n_1361),
.A2(n_1317),
.B(n_1272),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1364),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1369),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1375),
.A2(n_1323),
.B1(n_1357),
.B2(n_1352),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1376),
.A2(n_1379),
.B1(n_1377),
.B2(n_1383),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1371),
.B(n_1359),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1374),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1381),
.Y(n_1391)
);

XNOR2x2_ASAP7_75t_L g1392 ( 
.A(n_1372),
.B(n_1264),
.Y(n_1392)
);

INVx6_ASAP7_75t_L g1393 ( 
.A(n_1373),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1376),
.A2(n_1357),
.B(n_1353),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1391),
.Y(n_1395)
);

AO22x1_ASAP7_75t_L g1396 ( 
.A1(n_1394),
.A2(n_1386),
.B1(n_1385),
.B2(n_1370),
.Y(n_1396)
);

AOI211x1_ASAP7_75t_L g1397 ( 
.A1(n_1388),
.A2(n_1384),
.B(n_1378),
.C(n_1382),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1387),
.A2(n_1380),
.B1(n_1340),
.B2(n_1324),
.Y(n_1398)
);

NAND4xp25_ASAP7_75t_L g1399 ( 
.A(n_1390),
.B(n_1380),
.C(n_1351),
.D(n_1271),
.Y(n_1399)
);

NAND3xp33_ASAP7_75t_SL g1400 ( 
.A(n_1398),
.B(n_1392),
.C(n_1393),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1396),
.A2(n_1368),
.B(n_1393),
.Y(n_1401)
);

OAI21xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1395),
.A2(n_1389),
.B(n_1360),
.Y(n_1402)
);

XOR2x2_ASAP7_75t_L g1403 ( 
.A(n_1397),
.B(n_1256),
.Y(n_1403)
);

OAI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1399),
.A2(n_1336),
.B1(n_1316),
.B2(n_1345),
.Y(n_1404)
);

AOI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1396),
.A2(n_1366),
.B1(n_1271),
.B2(n_1265),
.Y(n_1405)
);

NOR4xp25_ASAP7_75t_L g1406 ( 
.A(n_1400),
.B(n_1255),
.C(n_1263),
.D(n_1344),
.Y(n_1406)
);

NOR3x1_ASAP7_75t_L g1407 ( 
.A(n_1403),
.B(n_1346),
.C(n_1289),
.Y(n_1407)
);

NOR2x1_ASAP7_75t_L g1408 ( 
.A(n_1401),
.B(n_1303),
.Y(n_1408)
);

NOR2x1_ASAP7_75t_L g1409 ( 
.A(n_1408),
.B(n_1404),
.Y(n_1409)
);

NOR2x1_ASAP7_75t_L g1410 ( 
.A(n_1406),
.B(n_1256),
.Y(n_1410)
);

NAND2x1_ASAP7_75t_L g1411 ( 
.A(n_1409),
.B(n_1405),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1411),
.A2(n_1410),
.B1(n_1402),
.B2(n_1407),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1412),
.A2(n_1185),
.B(n_1156),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1413),
.A2(n_1288),
.B1(n_1297),
.B2(n_1293),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1414),
.A2(n_1297),
.B1(n_1305),
.B2(n_1299),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_R g1416 ( 
.A1(n_1415),
.A2(n_1247),
.B1(n_1262),
.B2(n_1191),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1416),
.A2(n_1169),
.B1(n_1224),
.B2(n_1220),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1417),
.B(n_1360),
.Y(n_1418)
);

AOI211xp5_ASAP7_75t_L g1419 ( 
.A1(n_1418),
.A2(n_1250),
.B(n_1188),
.C(n_1191),
.Y(n_1419)
);


endmodule