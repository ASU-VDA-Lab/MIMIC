module real_jpeg_6112_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_0),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_0),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_0),
.Y(n_151)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_0),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_0),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_1),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_1),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_1),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_1),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_1),
.B(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_1),
.Y(n_236)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_3),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_3),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_3),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_3),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_3),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_3),
.B(n_241),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_3),
.B(n_385),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_4),
.B(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_4),
.A2(n_233),
.B(n_235),
.Y(n_232)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_4),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_4),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_4),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_4),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_4),
.B(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_4),
.B(n_394),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_5),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_6),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_6),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_6),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_6),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_6),
.B(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_6),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_6),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_6),
.B(n_408),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_7),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_7),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_7),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_7),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_7),
.B(n_256),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_7),
.B(n_241),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_7),
.B(n_390),
.Y(n_389)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_9),
.Y(n_146)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_9),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_9),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_10),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_10),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_10),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_10),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_10),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_10),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_10),
.B(n_303),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_11),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_11),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_11),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_11),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_11),
.B(n_177),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_12),
.Y(n_111)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_12),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_12),
.Y(n_234)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_14),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_14),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_14),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_14),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_14),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_14),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_15),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_15),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_199),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_197),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_164),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_19),
.B(n_164),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_92),
.C(n_122),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_20),
.B(n_92),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_57),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_39),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_22),
.B(n_39),
.C(n_57),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_33),
.C(n_37),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_23),
.B(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_26),
.C(n_30),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_49),
.C(n_53),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_24),
.A2(n_53),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_24),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_24),
.A2(n_30),
.B1(n_88),
.B2(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_24),
.A2(n_88),
.B1(n_366),
.B2(n_368),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_24),
.B(n_368),
.Y(n_410)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_25),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_26),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_26),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_26),
.A2(n_125),
.B1(n_192),
.B2(n_196),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_29),
.Y(n_149)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_29),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_30),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_30),
.B(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_30),
.A2(n_128),
.B1(n_263),
.B2(n_264),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_31),
.Y(n_359)
);

INVx8_ASAP7_75t_L g383 ( 
.A(n_31),
.Y(n_383)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g392 ( 
.A(n_32),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_33),
.A2(n_37),
.B1(n_47),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_33),
.Y(n_163)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_41),
.B1(n_42),
.B2(n_47),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_48),
.B1(n_55),
.B2(n_56),
.Y(n_39)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_42),
.B(n_47),
.C(n_56),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_45),
.Y(n_214)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_46),
.Y(n_133)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_46),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_46),
.Y(n_323)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_49),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_49),
.B(n_222),
.C(n_226),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_49),
.A2(n_90),
.B1(n_222),
.B2(n_293),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_76),
.C(n_86),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_58),
.B(n_76),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_64),
.B2(n_65),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_67),
.C(n_71),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_59),
.A2(n_60),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_59),
.B(n_115),
.C(n_121),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_59),
.A2(n_60),
.B1(n_141),
.B2(n_142),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_60),
.B(n_142),
.Y(n_300)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_71),
.B2(n_75),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_70),
.Y(n_173)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_70),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_70),
.Y(n_349)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.C(n_84),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_77),
.B(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_80),
.B(n_84),
.Y(n_138)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_83),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_86),
.B(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_112),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_94),
.B(n_95),
.C(n_112),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_109),
.B2(n_110),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_102),
.Y(n_225)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_103),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_104),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_104),
.B(n_107),
.C(n_110),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_104),
.B(n_131),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_130),
.C(n_134),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_111),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_121),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_115),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_118),
.A2(n_121),
.B1(n_176),
.B2(n_179),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_118),
.B(n_255),
.C(n_259),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_118),
.A2(n_121),
.B1(n_259),
.B2(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_122),
.B(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_139),
.C(n_161),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_123),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.C(n_137),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_124),
.Y(n_248)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_129),
.B(n_137),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_134),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_139),
.B(n_161),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_152),
.C(n_156),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_140),
.B(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_147),
.C(n_150),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_141),
.A2(n_142),
.B1(n_150),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_146),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_146),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_147),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_147),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_150),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_152),
.A2(n_156),
.B1(n_157),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_152),
.Y(n_246)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_155),
.Y(n_326)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_160),
.Y(n_243)
);

BUFx24_ASAP7_75t_SL g442 ( 
.A(n_164),
.Y(n_442)
);

FAx1_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_166),
.CI(n_180),
.CON(n_164),
.SN(n_164)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_210),
.C(n_215),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_171),
.A2(n_172),
.B1(n_210),
.B2(n_211),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_176),
.Y(n_179)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI221xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_338),
.B1(n_434),
.B2(n_439),
.C(n_440),
.Y(n_200)
);

NOR3xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_281),
.C(n_285),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_202),
.A2(n_435),
.B(n_438),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_274),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_203),
.B(n_274),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_247),
.C(n_250),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_204),
.B(n_247),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_230),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_205),
.B(n_231),
.C(n_244),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.C(n_220),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_207),
.B(n_221),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_209),
.B(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_214),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_215),
.B(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g367 ( 
.A(n_219),
.Y(n_367)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_222),
.Y(n_293)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_226),
.B(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_244),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_240),
.C(n_242),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_273),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_232),
.A2(n_235),
.B(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_242),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_250),
.B(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_267),
.C(n_272),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_251),
.B(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.C(n_261),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_252),
.B(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_254),
.A2(n_261),
.B1(n_262),
.B2(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_254),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_255),
.B(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_259),
.Y(n_318)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_260),
.Y(n_330)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_272),
.Y(n_289)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_280),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_278),
.C(n_280),
.Y(n_282)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_281),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_282),
.B(n_283),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_311),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_286),
.A2(n_436),
.B(n_437),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_309),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_287),
.B(n_309),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.C(n_307),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_288),
.B(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_290),
.B(n_307),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_294),
.C(n_298),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_294),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_296),
.B(n_372),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.C(n_304),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_299),
.A2(n_300),
.B1(n_422),
.B2(n_423),
.Y(n_421)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_301),
.A2(n_302),
.B1(n_304),
.B2(n_305),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_336),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_312),
.B(n_336),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.C(n_333),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_313),
.B(n_432),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_315),
.B(n_333),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.C(n_331),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_316),
.B(n_425),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_319),
.A2(n_331),
.B1(n_332),
.B2(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_319),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_324),
.C(n_327),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_320),
.A2(n_321),
.B1(n_327),
.B2(n_328),
.Y(n_414)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_324),
.B(n_414),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_325),
.B(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_339),
.A2(n_429),
.B(n_433),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_416),
.B(n_428),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_403),
.B(n_415),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_377),
.B(n_402),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_369),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_343),
.B(n_369),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_355),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_344),
.B(n_356),
.C(n_365),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_350),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_345),
.B(n_351),
.C(n_352),
.Y(n_412)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_365),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_360),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_360),
.Y(n_370)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx8_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_366),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.C(n_375),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_399),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_371),
.A2(n_375),
.B1(n_376),
.B2(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_371),
.Y(n_400)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_396),
.B(n_401),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_388),
.B(n_395),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_387),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_387),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_384),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_384),
.Y(n_397)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_SL g385 ( 
.A(n_386),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_393),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_391),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_397),
.B(n_398),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_404),
.B(n_405),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_411),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_406),
.A2(n_419),
.B1(n_420),
.B2(n_421),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_406),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_406),
.B(n_412),
.C(n_413),
.Y(n_427)
);

FAx1_ASAP7_75t_SL g406 ( 
.A(n_407),
.B(n_409),
.CI(n_410),
.CON(n_406),
.SN(n_406)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_427),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_417),
.B(n_427),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_424),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_421),
.C(n_424),
.Y(n_430)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_422),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_430),
.B(n_431),
.Y(n_433)
);


endmodule