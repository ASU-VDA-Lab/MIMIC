module real_aes_2600_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_764, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_765, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_764;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_765;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_532;
wire n_316;
wire n_284;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_753;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g183 ( .A(n_0), .B(n_157), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_1), .B(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_2), .B(n_127), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_3), .B(n_141), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_4), .B(n_159), .Y(n_480) );
INVx1_ASAP7_75t_L g148 ( .A(n_5), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_6), .B(n_141), .Y(n_210) );
NAND2xp33_ASAP7_75t_SL g253 ( .A(n_7), .B(n_147), .Y(n_253) );
XNOR2xp5_ASAP7_75t_L g743 ( .A(n_8), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g245 ( .A(n_9), .Y(n_245) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_10), .Y(n_120) );
AND2x2_ASAP7_75t_L g208 ( .A(n_11), .B(n_165), .Y(n_208) );
AND2x2_ASAP7_75t_L g482 ( .A(n_12), .B(n_161), .Y(n_482) );
AND2x2_ASAP7_75t_L g492 ( .A(n_13), .B(n_251), .Y(n_492) );
INVx2_ASAP7_75t_L g163 ( .A(n_14), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_15), .B(n_159), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_16), .Y(n_113) );
AOI221x1_ASAP7_75t_L g248 ( .A1(n_17), .A2(n_150), .B1(n_249), .B2(n_251), .C(n_252), .Y(n_248) );
AOI22xp5_ASAP7_75t_SL g744 ( .A1(n_18), .A2(n_75), .B1(n_745), .B2(n_746), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_18), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_19), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_20), .B(n_141), .Y(n_537) );
INVx1_ASAP7_75t_L g117 ( .A(n_21), .Y(n_117) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_22), .A2(n_91), .B1(n_141), .B2(n_194), .Y(n_496) );
AOI221xp5_ASAP7_75t_SL g172 ( .A1(n_23), .A2(n_39), .B1(n_141), .B2(n_150), .C(n_173), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_24), .A2(n_150), .B(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_25), .B(n_157), .Y(n_213) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_26), .A2(n_90), .B(n_163), .Y(n_162) );
OR2x2_ASAP7_75t_L g166 ( .A(n_26), .B(n_90), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_27), .B(n_159), .Y(n_158) );
INVxp67_ASAP7_75t_L g247 ( .A(n_28), .Y(n_247) );
AND2x2_ASAP7_75t_L g234 ( .A(n_29), .B(n_171), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_30), .A2(n_150), .B(n_182), .Y(n_181) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_31), .A2(n_251), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_32), .B(n_159), .Y(n_174) );
OAI22xp5_ASAP7_75t_SL g447 ( .A1(n_33), .A2(n_72), .B1(n_448), .B2(n_449), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_33), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_34), .A2(n_150), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_35), .B(n_159), .Y(n_552) );
AND2x2_ASAP7_75t_L g147 ( .A(n_36), .B(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g151 ( .A(n_36), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g202 ( .A(n_36), .Y(n_202) );
OR2x6_ASAP7_75t_L g115 ( .A(n_37), .B(n_116), .Y(n_115) );
AOI221xp5_ASAP7_75t_L g102 ( .A1(n_38), .A2(n_103), .B1(n_121), .B2(n_124), .C(n_452), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_38), .A2(n_131), .B1(n_132), .B2(n_450), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_38), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_40), .B(n_141), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_41), .A2(n_83), .B1(n_150), .B2(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_42), .B(n_159), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_43), .B(n_141), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_44), .B(n_755), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_45), .B(n_157), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_46), .A2(n_150), .B(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g186 ( .A(n_47), .B(n_171), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_48), .B(n_157), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_49), .B(n_171), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_50), .B(n_141), .Y(n_529) );
INVx1_ASAP7_75t_L g144 ( .A(n_51), .Y(n_144) );
INVx1_ASAP7_75t_L g154 ( .A(n_51), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_52), .B(n_159), .Y(n_490) );
AND2x2_ASAP7_75t_L g519 ( .A(n_53), .B(n_171), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_54), .B(n_141), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_55), .B(n_157), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_56), .B(n_157), .Y(n_551) );
AND2x2_ASAP7_75t_L g225 ( .A(n_57), .B(n_171), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_58), .B(n_141), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_59), .B(n_159), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_60), .B(n_141), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_61), .A2(n_150), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_62), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_63), .B(n_157), .Y(n_222) );
AND2x2_ASAP7_75t_L g543 ( .A(n_64), .B(n_165), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_65), .A2(n_150), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_66), .B(n_159), .Y(n_214) );
AND2x2_ASAP7_75t_SL g205 ( .A(n_67), .B(n_161), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_68), .B(n_157), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_69), .B(n_157), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_70), .A2(n_93), .B1(n_150), .B2(n_200), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_71), .B(n_159), .Y(n_540) );
INVx1_ASAP7_75t_L g448 ( .A(n_72), .Y(n_448) );
INVx1_ASAP7_75t_L g146 ( .A(n_73), .Y(n_146) );
INVx1_ASAP7_75t_L g152 ( .A(n_73), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_74), .B(n_157), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_75), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_76), .A2(n_150), .B(n_523), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_77), .A2(n_150), .B(n_470), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_78), .A2(n_150), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g554 ( .A(n_79), .B(n_165), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_80), .B(n_171), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_81), .A2(n_85), .B1(n_141), .B2(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_82), .B(n_141), .Y(n_223) );
INVx1_ASAP7_75t_L g118 ( .A(n_84), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_86), .B(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_87), .B(n_157), .Y(n_175) );
AND2x2_ASAP7_75t_L g473 ( .A(n_88), .B(n_161), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_89), .A2(n_150), .B(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_92), .B(n_159), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_94), .A2(n_150), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_95), .B(n_159), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_96), .B(n_141), .Y(n_185) );
INVxp67_ASAP7_75t_L g250 ( .A(n_97), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_98), .B(n_159), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_99), .A2(n_150), .B(n_155), .Y(n_149) );
BUFx2_ASAP7_75t_L g542 ( .A(n_100), .Y(n_542) );
BUFx2_ASAP7_75t_SL g109 ( .A(n_101), .Y(n_109) );
BUFx2_ASAP7_75t_L g123 ( .A(n_101), .Y(n_123) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_110), .B(n_119), .Y(n_106) );
CKINVDCx11_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx8_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx3_ASAP7_75t_L g128 ( .A(n_112), .Y(n_128) );
BUFx2_ASAP7_75t_L g762 ( .A(n_112), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AND2x6_ASAP7_75t_SL g456 ( .A(n_113), .B(n_115), .Y(n_456) );
OR2x6_ASAP7_75t_SL g742 ( .A(n_113), .B(n_114), .Y(n_742) );
OR2x2_ASAP7_75t_L g756 ( .A(n_113), .B(n_115), .Y(n_756) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
OR2x2_ASAP7_75t_SL g122 ( .A(n_119), .B(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g761 ( .A(n_119), .Y(n_761) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g760 ( .A(n_123), .B(n_761), .Y(n_760) );
OAI21xp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_129), .B(n_451), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
CKINVDCx11_ASAP7_75t_R g126 ( .A(n_127), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_128), .Y(n_127) );
INVxp33_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g450 ( .A(n_132), .Y(n_450) );
XNOR2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_447), .Y(n_132) );
AOI22xp5_ASAP7_75t_SL g455 ( .A1(n_133), .A2(n_456), .B1(n_457), .B2(n_741), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_133), .A2(n_457), .B1(n_750), .B2(n_753), .Y(n_749) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_339), .Y(n_133) );
NOR3xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_267), .C(n_317), .Y(n_134) );
OAI211xp5_ASAP7_75t_SL g135 ( .A1(n_136), .A2(n_187), .B(n_235), .C(n_256), .Y(n_135) );
OR2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_167), .Y(n_136) );
AND2x2_ASAP7_75t_L g266 ( .A(n_137), .B(n_168), .Y(n_266) );
INVx1_ASAP7_75t_L g397 ( .A(n_137), .Y(n_397) );
NOR2x1p5_ASAP7_75t_L g429 ( .A(n_137), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g240 ( .A(n_138), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g288 ( .A(n_138), .Y(n_288) );
OR2x2_ASAP7_75t_L g292 ( .A(n_138), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_138), .B(n_170), .Y(n_304) );
OR2x2_ASAP7_75t_L g326 ( .A(n_138), .B(n_170), .Y(n_326) );
AND2x4_ASAP7_75t_L g332 ( .A(n_138), .B(n_296), .Y(n_332) );
OR2x2_ASAP7_75t_L g349 ( .A(n_138), .B(n_242), .Y(n_349) );
INVx1_ASAP7_75t_L g384 ( .A(n_138), .Y(n_384) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_138), .Y(n_406) );
OR2x2_ASAP7_75t_L g420 ( .A(n_138), .B(n_353), .Y(n_420) );
AND2x4_ASAP7_75t_SL g424 ( .A(n_138), .B(n_242), .Y(n_424) );
OR2x6_ASAP7_75t_L g138 ( .A(n_139), .B(n_164), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_149), .B(n_161), .Y(n_139) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_147), .Y(n_141) );
INVx1_ASAP7_75t_L g254 ( .A(n_142), .Y(n_254) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
AND2x6_ASAP7_75t_L g157 ( .A(n_143), .B(n_152), .Y(n_157) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_L g159 ( .A(n_145), .B(n_154), .Y(n_159) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx5_ASAP7_75t_L g160 ( .A(n_147), .Y(n_160) );
AND2x2_ASAP7_75t_L g153 ( .A(n_148), .B(n_154), .Y(n_153) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_148), .Y(n_197) );
AND2x6_ASAP7_75t_L g150 ( .A(n_151), .B(n_153), .Y(n_150) );
BUFx3_ASAP7_75t_L g198 ( .A(n_151), .Y(n_198) );
INVx2_ASAP7_75t_L g204 ( .A(n_152), .Y(n_204) );
AND2x4_ASAP7_75t_L g200 ( .A(n_153), .B(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g196 ( .A(n_154), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_158), .B(n_160), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_157), .B(n_542), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_160), .A2(n_174), .B(n_175), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_160), .A2(n_183), .B(n_184), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_160), .A2(n_213), .B(n_214), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_160), .A2(n_221), .B(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_160), .A2(n_231), .B(n_232), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_160), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_160), .A2(n_479), .B(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_160), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_160), .A2(n_524), .B(n_525), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_160), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_160), .A2(n_540), .B(n_541), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_160), .A2(n_551), .B(n_552), .Y(n_550) );
INVx2_ASAP7_75t_SL g191 ( .A(n_161), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_161), .A2(n_537), .B(n_538), .Y(n_536) );
BUFx4f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx3_ASAP7_75t_L g179 ( .A(n_162), .Y(n_179) );
AND2x2_ASAP7_75t_SL g165 ( .A(n_163), .B(n_166), .Y(n_165) );
AND2x4_ASAP7_75t_L g215 ( .A(n_163), .B(n_166), .Y(n_215) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_165), .Y(n_171) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g376 ( .A(n_168), .B(n_332), .Y(n_376) );
AND2x2_ASAP7_75t_L g423 ( .A(n_168), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_177), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g239 ( .A(n_170), .Y(n_239) );
AND2x2_ASAP7_75t_L g286 ( .A(n_170), .B(n_177), .Y(n_286) );
INVx2_ASAP7_75t_L g293 ( .A(n_170), .Y(n_293) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_170), .Y(n_414) );
BUFx3_ASAP7_75t_L g430 ( .A(n_170), .Y(n_430) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_176), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_171), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_171), .A2(n_468), .B(n_469), .Y(n_467) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_171), .A2(n_496), .B(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g255 ( .A(n_177), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_177), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g353 ( .A(n_177), .B(n_293), .Y(n_353) );
INVx1_ASAP7_75t_L g371 ( .A(n_177), .Y(n_371) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_177), .Y(n_387) );
INVx1_ASAP7_75t_L g409 ( .A(n_177), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_177), .B(n_288), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_177), .B(n_242), .Y(n_446) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AOI21x1_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_186), .Y(n_178) );
INVx4_ASAP7_75t_L g251 ( .A(n_179), .Y(n_251) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_179), .A2(n_486), .B(n_492), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_181), .B(n_185), .Y(n_180) );
INVx1_ASAP7_75t_SL g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_206), .Y(n_188) );
AND2x4_ASAP7_75t_L g260 ( .A(n_189), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g271 ( .A(n_189), .Y(n_271) );
AND2x2_ASAP7_75t_L g276 ( .A(n_189), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g311 ( .A(n_189), .B(n_216), .Y(n_311) );
AND2x2_ASAP7_75t_L g321 ( .A(n_189), .B(n_217), .Y(n_321) );
OR2x2_ASAP7_75t_L g401 ( .A(n_189), .B(n_316), .Y(n_401) );
OAI322xp33_ASAP7_75t_L g431 ( .A1(n_189), .A2(n_344), .A3(n_383), .B1(n_416), .B2(n_432), .C1(n_433), .C2(n_434), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_189), .B(n_414), .Y(n_432) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g265 ( .A(n_190), .Y(n_265) );
AOI21x1_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_205), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_199), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_194), .A2(n_200), .B1(n_244), .B2(n_246), .Y(n_243) );
AND2x4_ASAP7_75t_L g194 ( .A(n_195), .B(n_198), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
NOR2x1p5_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
INVx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_206), .A2(n_378), .B1(n_382), .B2(n_385), .Y(n_377) );
AOI211xp5_ASAP7_75t_L g437 ( .A1(n_206), .A2(n_438), .B(n_439), .C(n_442), .Y(n_437) );
AND2x4_ASAP7_75t_SL g206 ( .A(n_207), .B(n_216), .Y(n_206) );
AND2x4_ASAP7_75t_L g259 ( .A(n_207), .B(n_227), .Y(n_259) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_207), .Y(n_263) );
INVx5_ASAP7_75t_L g275 ( .A(n_207), .Y(n_275) );
INVx2_ASAP7_75t_L g284 ( .A(n_207), .Y(n_284) );
AND2x2_ASAP7_75t_L g307 ( .A(n_207), .B(n_217), .Y(n_307) );
AND2x2_ASAP7_75t_L g336 ( .A(n_207), .B(n_226), .Y(n_336) );
OR2x2_ASAP7_75t_L g345 ( .A(n_207), .B(n_265), .Y(n_345) );
OR2x2_ASAP7_75t_L g360 ( .A(n_207), .B(n_274), .Y(n_360) );
OR2x6_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_215), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_215), .B(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_215), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_215), .B(n_250), .Y(n_249) );
NOR3xp33_ASAP7_75t_L g252 ( .A(n_215), .B(n_253), .C(n_254), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_215), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_215), .A2(n_529), .B(n_530), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_216), .B(n_236), .Y(n_235) );
INVx3_ASAP7_75t_SL g344 ( .A(n_216), .Y(n_344) );
AND2x2_ASAP7_75t_L g367 ( .A(n_216), .B(n_275), .Y(n_367) );
AND2x4_ASAP7_75t_L g216 ( .A(n_217), .B(n_226), .Y(n_216) );
INVx2_ASAP7_75t_L g261 ( .A(n_217), .Y(n_261) );
AND2x2_ASAP7_75t_L g264 ( .A(n_217), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g278 ( .A(n_217), .B(n_227), .Y(n_278) );
INVx1_ASAP7_75t_L g282 ( .A(n_217), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_217), .B(n_227), .Y(n_316) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_217), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_217), .B(n_275), .Y(n_391) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_224), .B(n_225), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_223), .Y(n_218) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_224), .A2(n_228), .B(n_234), .Y(n_227) );
AO21x2_ASAP7_75t_L g274 ( .A1(n_224), .A2(n_228), .B(n_234), .Y(n_274) );
AOI21x1_ASAP7_75t_L g475 ( .A1(n_224), .A2(n_476), .B(n_482), .Y(n_475) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_227), .Y(n_297) );
AND2x2_ASAP7_75t_L g381 ( .A(n_227), .B(n_265), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_233), .Y(n_228) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_240), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_237), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OR2x6_ASAP7_75t_SL g445 ( .A(n_238), .B(n_446), .Y(n_445) );
INVxp67_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_239), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_239), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g393 ( .A(n_239), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_240), .A2(n_302), .B1(n_305), .B2(n_312), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_241), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g337 ( .A(n_241), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_241), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_SL g392 ( .A(n_241), .B(n_393), .Y(n_392) );
AND2x4_ASAP7_75t_L g241 ( .A(n_242), .B(n_255), .Y(n_241) );
AND2x2_ASAP7_75t_L g287 ( .A(n_242), .B(n_288), .Y(n_287) );
INVx3_ASAP7_75t_L g296 ( .A(n_242), .Y(n_296) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_242), .A2(n_303), .B1(n_355), .B2(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g362 ( .A(n_242), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_242), .B(n_356), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_242), .B(n_286), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_242), .B(n_293), .Y(n_435) );
AND2x4_ASAP7_75t_L g242 ( .A(n_243), .B(n_248), .Y(n_242) );
INVx3_ASAP7_75t_L g547 ( .A(n_251), .Y(n_547) );
OAI21xp33_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_262), .B(n_266), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
NAND4xp25_ASAP7_75t_SL g305 ( .A(n_258), .B(n_306), .C(n_308), .D(n_310), .Y(n_305) );
INVx2_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_259), .B(n_366), .Y(n_395) );
AND2x2_ASAP7_75t_L g422 ( .A(n_259), .B(n_260), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_259), .B(n_282), .Y(n_433) );
INVx1_ASAP7_75t_L g298 ( .A(n_260), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_260), .A2(n_323), .B1(n_334), .B2(n_337), .Y(n_333) );
NAND3xp33_ASAP7_75t_L g355 ( .A(n_260), .B(n_273), .C(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_260), .B(n_275), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_260), .B(n_283), .Y(n_426) );
AND2x2_ASAP7_75t_L g358 ( .A(n_261), .B(n_265), .Y(n_358) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_261), .Y(n_419) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g314 ( .A(n_263), .Y(n_314) );
INVx1_ASAP7_75t_L g404 ( .A(n_264), .Y(n_404) );
AND2x2_ASAP7_75t_L g411 ( .A(n_264), .B(n_275), .Y(n_411) );
BUFx2_ASAP7_75t_L g366 ( .A(n_265), .Y(n_366) );
NAND3xp33_ASAP7_75t_SL g267 ( .A(n_268), .B(n_289), .C(n_301), .Y(n_267) );
OAI31xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_276), .A3(n_279), .B(n_285), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g322 ( .A1(n_269), .A2(n_323), .B1(n_327), .B2(n_328), .Y(n_322) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
OR2x2_ASAP7_75t_L g308 ( .A(n_271), .B(n_309), .Y(n_308) );
NOR2x1_ASAP7_75t_L g334 ( .A(n_271), .B(n_335), .Y(n_334) );
O2A1O1Ixp33_ASAP7_75t_L g403 ( .A1(n_272), .A2(n_374), .B(n_404), .C(n_405), .Y(n_403) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_273), .B(n_419), .Y(n_418) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_274), .B(n_282), .Y(n_309) );
AND2x2_ASAP7_75t_L g327 ( .A(n_274), .B(n_307), .Y(n_327) );
AND2x2_ASAP7_75t_L g444 ( .A(n_277), .B(n_366), .Y(n_444) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g300 ( .A(n_278), .B(n_284), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_283), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g375 ( .A(n_283), .B(n_358), .Y(n_375) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_284), .B(n_358), .Y(n_364) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx2_ASAP7_75t_L g356 ( .A(n_286), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_287), .B(n_387), .Y(n_386) );
AOI32xp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_297), .A3(n_298), .B1(n_299), .B2(n_764), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_290), .A2(n_375), .B1(n_411), .B2(n_412), .C(n_415), .Y(n_410) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_294), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_293), .Y(n_338) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g303 ( .A(n_295), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g408 ( .A(n_296), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_297), .B(n_319), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_299), .A2(n_342), .B1(n_346), .B2(n_350), .C(n_354), .Y(n_341) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI211xp5_ASAP7_75t_L g317 ( .A1(n_304), .A2(n_318), .B(n_322), .C(n_333), .Y(n_317) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI322xp33_ASAP7_75t_L g415 ( .A1(n_310), .A2(n_320), .A3(n_369), .B1(n_416), .B2(n_417), .C1(n_418), .C2(n_420), .Y(n_415) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AOI21xp33_ASAP7_75t_L g442 ( .A1(n_313), .A2(n_443), .B(n_445), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_L g399 ( .A1(n_319), .A2(n_400), .B(n_402), .C(n_403), .Y(n_399) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g441 ( .A(n_326), .B(n_407), .Y(n_441) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_332), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g416 ( .A(n_332), .Y(n_416) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI31xp33_ASAP7_75t_L g372 ( .A1(n_336), .A2(n_373), .A3(n_375), .B(n_376), .Y(n_372) );
NOR2x1_ASAP7_75t_L g339 ( .A(n_340), .B(n_398), .Y(n_339) );
NAND5xp2_ASAP7_75t_L g340 ( .A(n_341), .B(n_361), .C(n_372), .D(n_377), .E(n_388), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AOI21xp33_ASAP7_75t_L g439 ( .A1(n_344), .A2(n_440), .B(n_441), .Y(n_439) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g412 ( .A(n_348), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
A2O1A1Ixp33_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_363), .B(n_365), .C(n_368), .Y(n_361) );
INVxp33_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
OR2x2_ASAP7_75t_L g390 ( .A(n_366), .B(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_369), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_SL g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g440 ( .A(n_381), .Y(n_440) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_392), .B(n_394), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI21xp33_ASAP7_75t_L g394 ( .A1(n_390), .A2(n_395), .B(n_396), .Y(n_394) );
NAND4xp25_ASAP7_75t_L g398 ( .A(n_399), .B(n_410), .C(n_421), .D(n_437), .Y(n_398) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_408), .B(n_429), .Y(n_428) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g438 ( .A(n_420), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B1(n_425), .B2(n_427), .C(n_431), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI31xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_747), .A3(n_754), .B(n_757), .Y(n_452) );
INVxp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_743), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g752 ( .A(n_456), .Y(n_752) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_654), .Y(n_457) );
NOR4xp75_ASAP7_75t_L g458 ( .A(n_459), .B(n_577), .C(n_602), .D(n_629), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_514), .B(n_555), .Y(n_459) );
NOR4xp25_ASAP7_75t_L g460 ( .A(n_461), .B(n_498), .C(n_505), .D(n_509), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_483), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_474), .Y(n_464) );
NAND2x1p5_ASAP7_75t_L g617 ( .A(n_465), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_465), .B(n_502), .Y(n_648) );
AND2x2_ASAP7_75t_L g673 ( .A(n_465), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g698 ( .A(n_465), .B(n_493), .Y(n_698) );
AND2x2_ASAP7_75t_L g739 ( .A(n_465), .B(n_507), .Y(n_739) );
INVx4_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_SL g511 ( .A(n_466), .B(n_504), .Y(n_511) );
AND2x2_ASAP7_75t_L g513 ( .A(n_466), .B(n_485), .Y(n_513) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_466), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g574 ( .A(n_466), .Y(n_574) );
AND2x2_ASAP7_75t_L g580 ( .A(n_466), .B(n_507), .Y(n_580) );
BUFx2_ASAP7_75t_L g593 ( .A(n_466), .Y(n_593) );
AND2x4_ASAP7_75t_L g624 ( .A(n_466), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g671 ( .A(n_466), .B(n_672), .Y(n_671) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_473), .Y(n_466) );
INVx1_ASAP7_75t_L g665 ( .A(n_474), .Y(n_665) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g504 ( .A(n_475), .Y(n_504) );
AND2x2_ASAP7_75t_L g507 ( .A(n_475), .B(n_485), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_481), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_483), .B(n_683), .Y(n_736) );
INVx2_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
OR2x2_ASAP7_75t_L g573 ( .A(n_484), .B(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_493), .Y(n_484) );
INVx2_ASAP7_75t_L g503 ( .A(n_485), .Y(n_503) );
INVx2_ASAP7_75t_L g564 ( .A(n_485), .Y(n_564) );
AND2x2_ASAP7_75t_L g674 ( .A(n_485), .B(n_504), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_491), .Y(n_486) );
INVx2_ASAP7_75t_L g562 ( .A(n_493), .Y(n_562) );
BUFx3_ASAP7_75t_L g579 ( .A(n_493), .Y(n_579) );
AND2x2_ASAP7_75t_L g606 ( .A(n_493), .B(n_607), .Y(n_606) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
AND2x4_ASAP7_75t_L g500 ( .A(n_494), .B(n_495), .Y(n_500) );
NOR2x1_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
INVx2_ASAP7_75t_L g508 ( .A(n_499), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_499), .B(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g677 ( .A(n_499), .B(n_617), .Y(n_677) );
AND2x2_ASAP7_75t_L g701 ( .A(n_499), .B(n_511), .Y(n_701) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g597 ( .A(n_500), .B(n_503), .Y(n_597) );
AND2x2_ASAP7_75t_L g679 ( .A(n_500), .B(n_672), .Y(n_679) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_SL g722 ( .A(n_502), .Y(n_722) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
INVx1_ASAP7_75t_L g607 ( .A(n_503), .Y(n_607) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_504), .Y(n_611) );
INVx2_ASAP7_75t_L g619 ( .A(n_504), .Y(n_619) );
INVx1_ASAP7_75t_L g625 ( .A(n_504), .Y(n_625) );
AOI222xp33_ASAP7_75t_SL g555 ( .A1(n_505), .A2(n_556), .B1(n_560), .B2(n_565), .C1(n_572), .C2(n_575), .Y(n_555) );
INVx1_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g632 ( .A(n_507), .Y(n_632) );
BUFx2_ASAP7_75t_L g661 ( .A(n_507), .Y(n_661) );
OAI211xp5_ASAP7_75t_L g655 ( .A1(n_508), .A2(n_656), .B(n_660), .C(n_668), .Y(n_655) );
OR2x2_ASAP7_75t_L g726 ( .A(n_508), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g734 ( .A(n_508), .B(n_639), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_512), .Y(n_509) );
INVx2_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_SL g691 ( .A(n_511), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g709 ( .A(n_511), .B(n_597), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_511), .B(n_689), .Y(n_716) );
OR2x2_ASAP7_75t_L g717 ( .A(n_512), .B(n_579), .Y(n_717) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g639 ( .A(n_513), .B(n_611), .Y(n_639) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_534), .Y(n_515) );
INVx1_ASAP7_75t_L g733 ( .A(n_516), .Y(n_733) );
NOR2xp67_ASAP7_75t_L g516 ( .A(n_517), .B(n_526), .Y(n_516) );
AND2x2_ASAP7_75t_L g576 ( .A(n_517), .B(n_535), .Y(n_576) );
INVx1_ASAP7_75t_L g653 ( .A(n_517), .Y(n_653) );
OR2x2_ASAP7_75t_L g712 ( .A(n_517), .B(n_535), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_517), .B(n_584), .Y(n_718) );
INVx4_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g559 ( .A(n_518), .Y(n_559) );
OR2x2_ASAP7_75t_L g591 ( .A(n_518), .B(n_545), .Y(n_591) );
AND2x2_ASAP7_75t_L g600 ( .A(n_518), .B(n_527), .Y(n_600) );
NAND2x1_ASAP7_75t_L g628 ( .A(n_518), .B(n_535), .Y(n_628) );
AND2x2_ASAP7_75t_L g675 ( .A(n_518), .B(n_570), .Y(n_675) );
OR2x6_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g558 ( .A(n_527), .Y(n_558) );
INVx1_ASAP7_75t_L g568 ( .A(n_527), .Y(n_568) );
AND2x2_ASAP7_75t_L g584 ( .A(n_527), .B(n_571), .Y(n_584) );
INVx2_ASAP7_75t_L g589 ( .A(n_527), .Y(n_589) );
OR2x2_ASAP7_75t_L g685 ( .A(n_527), .B(n_535), .Y(n_685) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_544), .Y(n_534) );
NOR2x1_ASAP7_75t_SL g570 ( .A(n_535), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g588 ( .A(n_535), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g601 ( .A(n_535), .B(n_545), .Y(n_601) );
BUFx2_ASAP7_75t_L g620 ( .A(n_535), .Y(n_620) );
INVx2_ASAP7_75t_SL g647 ( .A(n_535), .Y(n_647) );
OR2x6_ASAP7_75t_L g535 ( .A(n_536), .B(n_543), .Y(n_535) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g557 ( .A(n_545), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g703 ( .A(n_545), .B(n_645), .Y(n_703) );
INVx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B(n_554), .Y(n_546) );
AO21x1_ASAP7_75t_SL g571 ( .A1(n_547), .A2(n_548), .B(n_554), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_553), .Y(n_548) );
AOI211xp5_ASAP7_75t_L g719 ( .A1(n_556), .A2(n_580), .B(n_720), .C(n_724), .Y(n_719) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_557), .B(n_635), .Y(n_670) );
BUFx2_ASAP7_75t_L g634 ( .A(n_558), .Y(n_634) );
OR2x2_ASAP7_75t_L g582 ( .A(n_559), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g667 ( .A(n_559), .B(n_601), .Y(n_667) );
AND2x2_ASAP7_75t_L g688 ( .A(n_559), .B(n_644), .Y(n_688) );
INVx2_ASAP7_75t_L g695 ( .A(n_559), .Y(n_695) );
OAI21xp5_ASAP7_75t_SL g700 ( .A1(n_560), .A2(n_701), .B(n_702), .Y(n_700) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
AND2x2_ASAP7_75t_L g642 ( .A(n_561), .B(n_624), .Y(n_642) );
OR2x2_ASAP7_75t_L g721 ( .A(n_561), .B(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_562), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_564), .Y(n_595) );
AND2x2_ASAP7_75t_L g672 ( .A(n_564), .B(n_619), .Y(n_672) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
AND2x2_ASAP7_75t_L g657 ( .A(n_567), .B(n_658), .Y(n_657) );
AND2x4_ASAP7_75t_SL g666 ( .A(n_567), .B(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_567), .B(n_576), .Y(n_699) );
INVx3_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g575 ( .A(n_568), .B(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g694 ( .A(n_569), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g644 ( .A(n_570), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g614 ( .A(n_571), .B(n_589), .Y(n_614) );
OAI31xp33_ASAP7_75t_L g621 ( .A1(n_572), .A2(n_622), .A3(n_624), .B(n_626), .Y(n_621) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_574), .B(n_597), .Y(n_623) );
AO21x1_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .B(n_585), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
OR2x2_ASAP7_75t_L g633 ( .A(n_579), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g738 ( .A(n_579), .Y(n_738) );
INVx2_ASAP7_75t_SL g723 ( .A(n_580), .Y(n_723) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g627 ( .A(n_583), .B(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g711 ( .A(n_583), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_584), .B(n_647), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_592), .B1(n_596), .B2(n_598), .Y(n_585) );
AOI21xp33_ASAP7_75t_L g704 ( .A1(n_586), .A2(n_705), .B(n_706), .Y(n_704) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x4_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx1_ASAP7_75t_L g645 ( .A(n_589), .Y(n_645) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g659 ( .A(n_591), .B(n_620), .Y(n_659) );
OR2x2_ASAP7_75t_L g684 ( .A(n_591), .B(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_593), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_593), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g683 ( .A(n_593), .Y(n_683) );
INVx2_ASAP7_75t_L g612 ( .A(n_594), .Y(n_612) );
INVx1_ASAP7_75t_L g692 ( .A(n_595), .Y(n_692) );
AND2x2_ASAP7_75t_L g615 ( .A(n_597), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g689 ( .A(n_597), .Y(n_689) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_603), .B(n_621), .Y(n_602) );
OAI321xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_608), .A3(n_613), .B1(n_614), .B2(n_615), .C(n_620), .Y(n_603) );
AOI322xp5_ASAP7_75t_L g729 ( .A1(n_604), .A2(n_635), .A3(n_730), .B1(n_732), .B2(n_734), .C1(n_735), .C2(n_740), .Y(n_729) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_L g682 ( .A(n_607), .Y(n_682) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_612), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_609), .B(n_689), .Y(n_706) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g714 ( .A(n_612), .Y(n_714) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp33_ASAP7_75t_SL g646 ( .A(n_614), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OAI21xp33_ASAP7_75t_SL g713 ( .A1(n_617), .A2(n_623), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx3_ASAP7_75t_L g635 ( .A(n_628), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_649), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_635), .B1(n_636), .B2(n_637), .C(n_640), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_632), .Y(n_651) );
AND2x2_ASAP7_75t_L g636 ( .A(n_634), .B(n_635), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI22xp33_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_643), .B1(n_646), .B2(n_648), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g652 ( .A(n_644), .B(n_653), .Y(n_652) );
OAI21xp33_ASAP7_75t_L g735 ( .A1(n_647), .A2(n_736), .B(n_737), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NOR3xp33_ASAP7_75t_SL g654 ( .A(n_655), .B(n_686), .C(n_707), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_659), .A2(n_694), .B1(n_721), .B2(n_723), .Y(n_720) );
OAI21xp33_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_662), .B(n_666), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_661), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_667), .A2(n_709), .B1(n_710), .B2(n_713), .C(n_715), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B1(n_673), .B2(n_675), .C(n_676), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g705 ( .A(n_671), .Y(n_705) );
INVx1_ASAP7_75t_L g727 ( .A(n_672), .Y(n_727) );
INVx1_ASAP7_75t_SL g725 ( .A(n_673), .Y(n_725) );
AOI31xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .A3(n_680), .B(n_684), .Y(n_676) );
OAI221xp5_ASAP7_75t_L g686 ( .A1(n_677), .A2(n_687), .B1(n_689), .B2(n_690), .C(n_765), .Y(n_686) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI211xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_693), .B(n_696), .C(n_704), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g702 ( .A(n_695), .B(n_703), .Y(n_702) );
OAI21xp5_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_699), .B(n_700), .Y(n_696) );
INVx1_ASAP7_75t_L g731 ( .A(n_703), .Y(n_731) );
BUFx2_ASAP7_75t_SL g740 ( .A(n_703), .Y(n_740) );
NAND3xp33_ASAP7_75t_SL g707 ( .A(n_708), .B(n_719), .C(n_729), .Y(n_707) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI21xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B(n_718), .Y(n_715) );
AOI21xp33_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .B(n_728), .Y(n_724) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVxp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx1_ASAP7_75t_SL g753 ( .A(n_741), .Y(n_753) );
CKINVDCx11_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g748 ( .A(n_743), .B(n_749), .Y(n_748) );
INVxp33_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx4_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVx3_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx3_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_762), .Y(n_758) );
INVxp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
endmodule