module real_aes_9036_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g265 ( .A1(n_0), .A2(n_266), .B(n_267), .C(n_270), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_1), .B(n_254), .Y(n_271) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_2), .B(n_108), .C(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g123 ( .A(n_2), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_3), .B(n_182), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_4), .A2(n_143), .B(n_146), .C(n_526), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_5), .A2(n_138), .B(n_550), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_6), .A2(n_138), .B(n_248), .Y(n_247) );
AOI222xp33_ASAP7_75t_SL g126 ( .A1(n_7), .A2(n_61), .B1(n_127), .B2(n_732), .C1(n_733), .C2(n_737), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_8), .B(n_254), .Y(n_556) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_9), .A2(n_173), .B(n_210), .Y(n_209) );
AND2x6_ASAP7_75t_L g143 ( .A(n_10), .B(n_144), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_11), .A2(n_143), .B(n_146), .C(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g494 ( .A(n_12), .Y(n_494) );
INVx1_ASAP7_75t_L g105 ( .A(n_13), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_13), .B(n_39), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_14), .B(n_230), .Y(n_528) );
INVx1_ASAP7_75t_L g164 ( .A(n_15), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_16), .B(n_182), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_17), .A2(n_183), .B(n_512), .C(n_514), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_18), .B(n_254), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_19), .B(n_158), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g145 ( .A1(n_20), .A2(n_146), .B(n_149), .C(n_157), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_21), .A2(n_218), .B(n_269), .C(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_22), .B(n_230), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_23), .B(n_230), .Y(n_467) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_24), .Y(n_541) );
INVx1_ASAP7_75t_L g466 ( .A(n_25), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_26), .A2(n_146), .B(n_157), .C(n_213), .Y(n_212) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_27), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_28), .Y(n_524) );
INVx1_ASAP7_75t_L g482 ( .A(n_29), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_30), .A2(n_138), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g141 ( .A(n_31), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_32), .A2(n_186), .B(n_195), .C(n_197), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_33), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_34), .A2(n_269), .B(n_553), .C(n_555), .Y(n_552) );
INVxp67_ASAP7_75t_L g483 ( .A(n_35), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_36), .B(n_215), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_37), .A2(n_146), .B(n_157), .C(n_465), .Y(n_464) );
CKINVDCx14_ASAP7_75t_R g551 ( .A(n_38), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_39), .B(n_105), .Y(n_104) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_40), .A2(n_270), .B(n_492), .C(n_493), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_41), .B(n_137), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_42), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_43), .B(n_182), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_44), .B(n_138), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_45), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_46), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_47), .A2(n_186), .B(n_195), .C(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g268 ( .A(n_48), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_49), .A2(n_128), .B1(n_735), .B2(n_744), .Y(n_743) );
CKINVDCx16_ASAP7_75t_R g744 ( .A(n_49), .Y(n_744) );
INVx1_ASAP7_75t_L g240 ( .A(n_50), .Y(n_240) );
INVx1_ASAP7_75t_L g500 ( .A(n_51), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_52), .B(n_138), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_53), .Y(n_166) );
CKINVDCx14_ASAP7_75t_R g490 ( .A(n_54), .Y(n_490) );
INVx1_ASAP7_75t_L g144 ( .A(n_55), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_56), .B(n_138), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_57), .B(n_254), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_58), .A2(n_156), .B(n_179), .C(n_251), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_59), .Y(n_125) );
INVx1_ASAP7_75t_L g163 ( .A(n_60), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_61), .Y(n_732) );
INVx1_ASAP7_75t_SL g554 ( .A(n_62), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_63), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_64), .B(n_182), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_65), .B(n_254), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_66), .B(n_183), .Y(n_228) );
INVx1_ASAP7_75t_L g544 ( .A(n_67), .Y(n_544) );
CKINVDCx16_ASAP7_75t_R g264 ( .A(n_68), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_69), .B(n_151), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_70), .A2(n_146), .B(n_177), .C(n_186), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_71), .A2(n_100), .B1(n_112), .B2(n_745), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g249 ( .A(n_72), .Y(n_249) );
INVx1_ASAP7_75t_L g111 ( .A(n_73), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_74), .A2(n_138), .B(n_489), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_75), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_76), .A2(n_138), .B(n_509), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_77), .A2(n_137), .B(n_478), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g463 ( .A(n_78), .Y(n_463) );
INVx1_ASAP7_75t_L g510 ( .A(n_79), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_80), .B(n_154), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_81), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_82), .A2(n_138), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g513 ( .A(n_83), .Y(n_513) );
INVx2_ASAP7_75t_L g161 ( .A(n_84), .Y(n_161) );
INVx1_ASAP7_75t_L g527 ( .A(n_85), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_86), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_87), .B(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g108 ( .A(n_88), .Y(n_108) );
OR2x2_ASAP7_75t_L g120 ( .A(n_88), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g455 ( .A(n_88), .B(n_122), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_89), .A2(n_146), .B(n_186), .C(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_90), .B(n_138), .Y(n_193) );
INVx1_ASAP7_75t_L g198 ( .A(n_91), .Y(n_198) );
INVxp67_ASAP7_75t_L g252 ( .A(n_92), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_93), .B(n_173), .Y(n_495) );
INVx2_ASAP7_75t_L g503 ( .A(n_94), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_95), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g178 ( .A(n_96), .Y(n_178) );
INVx1_ASAP7_75t_L g224 ( .A(n_97), .Y(n_224) );
AND2x2_ASAP7_75t_L g242 ( .A(n_98), .B(n_160), .Y(n_242) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_SL g745 ( .A(n_102), .Y(n_745) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g731 ( .A(n_108), .B(n_122), .Y(n_731) );
NOR2x2_ASAP7_75t_L g739 ( .A(n_108), .B(n_121), .Y(n_739) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AOI22x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_126), .B1(n_740), .B2(n_742), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_117), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g741 ( .A(n_116), .Y(n_741) );
AOI21xp5_ASAP7_75t_L g742 ( .A1(n_117), .A2(n_120), .B(n_743), .Y(n_742) );
NOR2xp33_ASAP7_75t_SL g117 ( .A(n_118), .B(n_125), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_453), .B1(n_456), .B2(n_729), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx2_ASAP7_75t_L g735 ( .A(n_129), .Y(n_735) );
AND3x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_357), .C(n_414), .Y(n_129) );
NOR3xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_302), .C(n_338), .Y(n_130) );
OAI211xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_204), .B(n_256), .C(n_289), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_168), .Y(n_132) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g259 ( .A(n_134), .B(n_260), .Y(n_259) );
INVx5_ASAP7_75t_L g288 ( .A(n_134), .Y(n_288) );
AND2x2_ASAP7_75t_L g361 ( .A(n_134), .B(n_277), .Y(n_361) );
AND2x2_ASAP7_75t_L g399 ( .A(n_134), .B(n_305), .Y(n_399) );
AND2x2_ASAP7_75t_L g419 ( .A(n_134), .B(n_261), .Y(n_419) );
OR2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_165), .Y(n_134) );
AOI21xp5_ASAP7_75t_SL g135 ( .A1(n_136), .A2(n_145), .B(n_158), .Y(n_135) );
BUFx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
NAND2x1p5_ASAP7_75t_L g225 ( .A(n_139), .B(n_143), .Y(n_225) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g156 ( .A(n_140), .Y(n_156) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
INVx1_ASAP7_75t_L g219 ( .A(n_141), .Y(n_219) );
INVx1_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_142), .Y(n_152) );
INVx3_ASAP7_75t_L g183 ( .A(n_142), .Y(n_183) );
INVx1_ASAP7_75t_L g215 ( .A(n_142), .Y(n_215) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_142), .Y(n_230) );
BUFx3_ASAP7_75t_L g157 ( .A(n_143), .Y(n_157) );
INVx4_ASAP7_75t_SL g187 ( .A(n_143), .Y(n_187) );
INVx5_ASAP7_75t_L g196 ( .A(n_146), .Y(n_196) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_147), .Y(n_185) );
BUFx3_ASAP7_75t_L g201 ( .A(n_147), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_153), .B(n_155), .Y(n_149) );
INVx2_ASAP7_75t_L g154 ( .A(n_151), .Y(n_154) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx4_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_154), .A2(n_198), .B(n_199), .C(n_200), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g239 ( .A1(n_154), .A2(n_200), .B(n_240), .C(n_241), .Y(n_239) );
O2A1O1Ixp5_ASAP7_75t_L g526 ( .A1(n_154), .A2(n_527), .B(n_528), .C(n_529), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_154), .A2(n_529), .B(n_544), .C(n_545), .Y(n_543) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_155), .A2(n_182), .B(n_466), .C(n_467), .Y(n_465) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_156), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_159), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g167 ( .A(n_160), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_160), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_160), .A2(n_237), .B(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_160), .A2(n_225), .B(n_463), .C(n_464), .Y(n_462) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_160), .A2(n_488), .B(n_495), .Y(n_487) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AND2x2_ASAP7_75t_L g174 ( .A(n_161), .B(n_162), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_167), .A2(n_523), .B(n_530), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_168), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_191), .Y(n_168) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_169), .Y(n_300) );
AND2x2_ASAP7_75t_L g314 ( .A(n_169), .B(n_260), .Y(n_314) );
INVx1_ASAP7_75t_L g337 ( .A(n_169), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_169), .B(n_288), .Y(n_376) );
OR2x2_ASAP7_75t_L g413 ( .A(n_169), .B(n_258), .Y(n_413) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_170), .Y(n_349) );
AND2x2_ASAP7_75t_L g356 ( .A(n_170), .B(n_261), .Y(n_356) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g277 ( .A(n_171), .B(n_261), .Y(n_277) );
BUFx2_ASAP7_75t_L g305 ( .A(n_171), .Y(n_305) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B(n_189), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_172), .B(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_172), .B(n_203), .Y(n_202) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_172), .A2(n_223), .B(n_231), .Y(n_222) );
INVx3_ASAP7_75t_L g254 ( .A(n_172), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_172), .B(n_469), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_172), .B(n_531), .Y(n_530) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_172), .A2(n_540), .B(n_546), .Y(n_539) );
INVx4_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_173), .A2(n_211), .B(n_212), .Y(n_210) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_173), .Y(n_246) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g233 ( .A(n_174), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_188), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_181), .C(n_184), .Y(n_177) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
OAI22xp33_ASAP7_75t_L g481 ( .A1(n_180), .A2(n_182), .B1(n_482), .B2(n_483), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_180), .B(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_180), .B(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_182), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g266 ( .A(n_182), .Y(n_266) );
INVx5_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_183), .B(n_494), .Y(n_493) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx3_ASAP7_75t_L g555 ( .A(n_185), .Y(n_555) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_187), .A2(n_196), .B(n_249), .C(n_250), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_SL g263 ( .A1(n_187), .A2(n_196), .B(n_264), .C(n_265), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_SL g478 ( .A1(n_187), .A2(n_196), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_SL g489 ( .A1(n_187), .A2(n_196), .B(n_490), .C(n_491), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_SL g499 ( .A1(n_187), .A2(n_196), .B(n_500), .C(n_501), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_SL g509 ( .A1(n_187), .A2(n_196), .B(n_510), .C(n_511), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g550 ( .A1(n_187), .A2(n_196), .B(n_551), .C(n_552), .Y(n_550) );
INVx5_ASAP7_75t_L g258 ( .A(n_191), .Y(n_258) );
BUFx2_ASAP7_75t_L g281 ( .A(n_191), .Y(n_281) );
AND2x2_ASAP7_75t_L g438 ( .A(n_191), .B(n_292), .Y(n_438) );
OR2x6_ASAP7_75t_L g191 ( .A(n_192), .B(n_202), .Y(n_191) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g270 ( .A(n_201), .Y(n_270) );
INVx1_ASAP7_75t_L g514 ( .A(n_201), .Y(n_514) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp33_ASAP7_75t_L g205 ( .A(n_206), .B(n_243), .Y(n_205) );
OAI221xp5_ASAP7_75t_L g338 ( .A1(n_206), .A2(n_339), .B1(n_346), .B2(n_347), .C(n_350), .Y(n_338) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_220), .Y(n_206) );
AND2x2_ASAP7_75t_L g244 ( .A(n_207), .B(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_207), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g273 ( .A(n_208), .B(n_221), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_208), .B(n_222), .Y(n_283) );
OR2x2_ASAP7_75t_L g294 ( .A(n_208), .B(n_245), .Y(n_294) );
AND2x2_ASAP7_75t_L g297 ( .A(n_208), .B(n_285), .Y(n_297) );
AND2x2_ASAP7_75t_L g313 ( .A(n_208), .B(n_234), .Y(n_313) );
OR2x2_ASAP7_75t_L g329 ( .A(n_208), .B(n_222), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_208), .B(n_245), .Y(n_391) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_209), .B(n_234), .Y(n_383) );
AND2x2_ASAP7_75t_L g386 ( .A(n_209), .B(n_222), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_216), .B(n_217), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_217), .A2(n_228), .B(n_229), .Y(n_227) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_L g307 ( .A(n_220), .B(n_294), .Y(n_307) );
INVx2_ASAP7_75t_L g333 ( .A(n_220), .Y(n_333) );
OR2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_234), .Y(n_220) );
AND2x2_ASAP7_75t_L g255 ( .A(n_221), .B(n_235), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_221), .B(n_245), .Y(n_312) );
OR2x2_ASAP7_75t_L g323 ( .A(n_221), .B(n_235), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_221), .B(n_285), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g415 ( .A1(n_221), .A2(n_416), .B1(n_418), .B2(n_420), .C(n_423), .Y(n_415) );
INVx5_ASAP7_75t_SL g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_222), .B(n_245), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_226), .Y(n_223) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_225), .A2(n_524), .B(n_525), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_225), .A2(n_541), .B(n_542), .Y(n_540) );
INVx4_ASAP7_75t_L g269 ( .A(n_230), .Y(n_269) );
INVx2_ASAP7_75t_L g492 ( .A(n_230), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g475 ( .A(n_233), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_234), .B(n_285), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_234), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g301 ( .A(n_234), .B(n_273), .Y(n_301) );
OR2x2_ASAP7_75t_L g345 ( .A(n_234), .B(n_245), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_234), .B(n_297), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_234), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g410 ( .A(n_234), .B(n_411), .Y(n_410) );
INVx5_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_SL g274 ( .A(n_235), .B(n_244), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_SL g278 ( .A1(n_235), .A2(n_279), .B(n_282), .C(n_286), .Y(n_278) );
OR2x2_ASAP7_75t_L g316 ( .A(n_235), .B(n_312), .Y(n_316) );
OR2x2_ASAP7_75t_L g352 ( .A(n_235), .B(n_294), .Y(n_352) );
OAI311xp33_ASAP7_75t_L g358 ( .A1(n_235), .A2(n_297), .A3(n_359), .B1(n_362), .C1(n_369), .Y(n_358) );
AND2x2_ASAP7_75t_L g409 ( .A(n_235), .B(n_245), .Y(n_409) );
AND2x2_ASAP7_75t_L g417 ( .A(n_235), .B(n_272), .Y(n_417) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_235), .Y(n_435) );
AND2x2_ASAP7_75t_L g452 ( .A(n_235), .B(n_273), .Y(n_452) );
OR2x6_ASAP7_75t_L g235 ( .A(n_236), .B(n_242), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_255), .Y(n_243) );
AND2x2_ASAP7_75t_L g280 ( .A(n_244), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g436 ( .A(n_244), .Y(n_436) );
AND2x2_ASAP7_75t_L g272 ( .A(n_245), .B(n_273), .Y(n_272) );
INVx3_ASAP7_75t_L g285 ( .A(n_245), .Y(n_285) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_245), .Y(n_328) );
INVxp67_ASAP7_75t_L g367 ( .A(n_245), .Y(n_367) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_247), .B(n_253), .Y(n_245) );
OA21x2_ASAP7_75t_L g497 ( .A1(n_246), .A2(n_498), .B(n_504), .Y(n_497) );
OA21x2_ASAP7_75t_L g507 ( .A1(n_246), .A2(n_508), .B(n_515), .Y(n_507) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_246), .A2(n_549), .B(n_556), .Y(n_548) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_254), .A2(n_262), .B(n_271), .Y(n_261) );
AND2x2_ASAP7_75t_L g445 ( .A(n_255), .B(n_293), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_272), .B1(n_274), .B2(n_275), .C(n_278), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_258), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g298 ( .A(n_258), .B(n_288), .Y(n_298) );
AND2x2_ASAP7_75t_L g306 ( .A(n_258), .B(n_260), .Y(n_306) );
OR2x2_ASAP7_75t_L g318 ( .A(n_258), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g336 ( .A(n_258), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g360 ( .A(n_258), .B(n_361), .Y(n_360) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_258), .Y(n_380) );
AND2x2_ASAP7_75t_L g432 ( .A(n_258), .B(n_356), .Y(n_432) );
OAI31xp33_ASAP7_75t_L g440 ( .A1(n_258), .A2(n_309), .A3(n_408), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_259), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g404 ( .A(n_259), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_259), .B(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g292 ( .A(n_260), .B(n_288), .Y(n_292) );
INVx1_ASAP7_75t_L g379 ( .A(n_260), .Y(n_379) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g429 ( .A(n_261), .B(n_288), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_269), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g529 ( .A(n_270), .Y(n_529) );
INVx1_ASAP7_75t_SL g439 ( .A(n_272), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_273), .B(n_344), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_274), .A2(n_386), .B1(n_424), .B2(n_427), .Y(n_423) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g287 ( .A(n_277), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g346 ( .A(n_277), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_277), .B(n_298), .Y(n_451) );
INVx1_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g421 ( .A(n_280), .B(n_422), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_281), .A2(n_340), .B(n_342), .Y(n_339) );
OR2x2_ASAP7_75t_L g347 ( .A(n_281), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g368 ( .A(n_281), .B(n_356), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_281), .B(n_379), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_281), .B(n_419), .Y(n_418) );
OAI221xp5_ASAP7_75t_SL g395 ( .A1(n_282), .A2(n_396), .B1(n_401), .B2(n_404), .C(n_405), .Y(n_395) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
OR2x2_ASAP7_75t_L g372 ( .A(n_283), .B(n_345), .Y(n_372) );
INVx1_ASAP7_75t_L g411 ( .A(n_283), .Y(n_411) );
INVx2_ASAP7_75t_L g387 ( .A(n_284), .Y(n_387) );
INVx1_ASAP7_75t_L g321 ( .A(n_285), .Y(n_321) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g326 ( .A(n_288), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_288), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g355 ( .A(n_288), .B(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g443 ( .A(n_288), .B(n_413), .Y(n_443) );
AOI222xp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_293), .B1(n_295), .B2(n_298), .C1(n_299), .C2(n_301), .Y(n_289) );
INVxp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g299 ( .A(n_292), .B(n_300), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_292), .A2(n_342), .B1(n_370), .B2(n_371), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_292), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
OAI21xp33_ASAP7_75t_SL g330 ( .A1(n_301), .A2(n_331), .B(n_334), .Y(n_330) );
OAI211xp5_ASAP7_75t_SL g302 ( .A1(n_303), .A2(n_307), .B(n_308), .C(n_330), .Y(n_302) );
INVxp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AOI221xp5_ASAP7_75t_L g308 ( .A1(n_306), .A2(n_309), .B1(n_314), .B2(n_315), .C(n_317), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_306), .B(n_394), .Y(n_393) );
INVxp67_ASAP7_75t_L g400 ( .A(n_306), .Y(n_400) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
AND2x2_ASAP7_75t_L g402 ( .A(n_311), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g319 ( .A(n_314), .Y(n_319) );
AND2x2_ASAP7_75t_L g325 ( .A(n_314), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_320), .B1(n_324), .B2(n_327), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_321), .B(n_333), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_322), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g422 ( .A(n_326), .Y(n_422) );
AND2x2_ASAP7_75t_L g441 ( .A(n_326), .B(n_356), .Y(n_441) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_333), .B(n_390), .Y(n_449) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_336), .B(n_404), .Y(n_447) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g370 ( .A(n_348), .Y(n_370) );
BUFx2_ASAP7_75t_L g394 ( .A(n_349), .Y(n_394) );
OAI21xp5_ASAP7_75t_SL g350 ( .A1(n_351), .A2(n_353), .B(n_355), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR3xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_373), .C(n_395), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI21xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_365), .B(n_368), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
A2O1A1Ixp33_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_377), .B(n_381), .C(n_384), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_374), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NOR2xp67_ASAP7_75t_SL g378 ( .A(n_379), .B(n_380), .Y(n_378) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_SL g403 ( .A(n_383), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_388), .B(n_392), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
AND2x2_ASAP7_75t_L g408 ( .A(n_386), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_400), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B1(n_410), .B2(n_412), .Y(n_405) );
INVx2_ASAP7_75t_SL g426 ( .A(n_413), .Y(n_426) );
NOR3xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_430), .C(n_442), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVxp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_426), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B1(n_437), .B2(n_439), .C(n_440), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g442 ( .A1(n_431), .A2(n_443), .B(n_444), .C(n_446), .Y(n_442) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B1(n_450), .B2(n_452), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g734 ( .A(n_454), .Y(n_734) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g736 ( .A(n_456), .Y(n_736) );
OR5x1_ASAP7_75t_L g456 ( .A(n_457), .B(n_623), .C(n_687), .D(n_703), .E(n_718), .Y(n_456) );
NAND4xp25_ASAP7_75t_L g457 ( .A(n_458), .B(n_557), .C(n_584), .D(n_607), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_505), .B(n_516), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_470), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx3_ASAP7_75t_SL g536 ( .A(n_461), .Y(n_536) );
AND2x4_ASAP7_75t_L g570 ( .A(n_461), .B(n_559), .Y(n_570) );
OR2x2_ASAP7_75t_L g580 ( .A(n_461), .B(n_538), .Y(n_580) );
OR2x2_ASAP7_75t_L g626 ( .A(n_461), .B(n_473), .Y(n_626) );
AND2x2_ASAP7_75t_L g640 ( .A(n_461), .B(n_537), .Y(n_640) );
AND2x2_ASAP7_75t_L g683 ( .A(n_461), .B(n_573), .Y(n_683) );
AND2x2_ASAP7_75t_L g690 ( .A(n_461), .B(n_548), .Y(n_690) );
AND2x2_ASAP7_75t_L g709 ( .A(n_461), .B(n_599), .Y(n_709) );
AND2x2_ASAP7_75t_L g727 ( .A(n_461), .B(n_569), .Y(n_727) );
OR2x6_ASAP7_75t_L g461 ( .A(n_462), .B(n_468), .Y(n_461) );
INVx1_ASAP7_75t_L g692 ( .A(n_470), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_486), .Y(n_470) );
AND2x2_ASAP7_75t_L g602 ( .A(n_471), .B(n_537), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_471), .B(n_622), .Y(n_621) );
AOI32xp33_ASAP7_75t_L g635 ( .A1(n_471), .A2(n_636), .A3(n_639), .B1(n_641), .B2(n_645), .Y(n_635) );
AND2x2_ASAP7_75t_L g705 ( .A(n_471), .B(n_599), .Y(n_705) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g569 ( .A(n_473), .B(n_538), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_473), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g611 ( .A(n_473), .B(n_558), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_473), .B(n_690), .Y(n_689) );
AO21x2_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_476), .B(n_484), .Y(n_473) );
INVx1_ASAP7_75t_L g574 ( .A(n_474), .Y(n_574) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OA21x2_ASAP7_75t_L g573 ( .A1(n_477), .A2(n_485), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g576 ( .A(n_486), .B(n_520), .Y(n_576) );
AND2x2_ASAP7_75t_L g652 ( .A(n_486), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g724 ( .A(n_486), .Y(n_724) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_496), .Y(n_486) );
OR2x2_ASAP7_75t_L g519 ( .A(n_487), .B(n_497), .Y(n_519) );
AND2x2_ASAP7_75t_L g533 ( .A(n_487), .B(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_487), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g583 ( .A(n_487), .Y(n_583) );
AND2x2_ASAP7_75t_L g610 ( .A(n_487), .B(n_497), .Y(n_610) );
BUFx3_ASAP7_75t_L g613 ( .A(n_487), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_487), .B(n_588), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_487), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g564 ( .A(n_496), .Y(n_564) );
AND2x2_ASAP7_75t_L g582 ( .A(n_496), .B(n_562), .Y(n_582) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g593 ( .A(n_497), .B(n_507), .Y(n_593) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_497), .Y(n_606) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_506), .B(n_613), .Y(n_663) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_SL g534 ( .A(n_507), .Y(n_534) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_507), .B(n_582), .C(n_583), .Y(n_581) );
OR2x2_ASAP7_75t_L g589 ( .A(n_507), .B(n_562), .Y(n_589) );
AND2x2_ASAP7_75t_L g609 ( .A(n_507), .B(n_562), .Y(n_609) );
AND2x2_ASAP7_75t_L g653 ( .A(n_507), .B(n_522), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_532), .B(n_535), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_518), .B(n_520), .Y(n_517) );
AND2x2_ASAP7_75t_L g728 ( .A(n_518), .B(n_653), .Y(n_728) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_519), .A2(n_626), .B1(n_668), .B2(n_670), .Y(n_667) );
OR2x2_ASAP7_75t_L g674 ( .A(n_519), .B(n_589), .Y(n_674) );
OR2x2_ASAP7_75t_L g698 ( .A(n_519), .B(n_699), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_519), .B(n_618), .Y(n_711) );
AND2x2_ASAP7_75t_L g604 ( .A(n_520), .B(n_605), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_520), .A2(n_677), .B(n_692), .Y(n_691) );
AOI32xp33_ASAP7_75t_L g712 ( .A1(n_520), .A2(n_602), .A3(n_713), .B1(n_715), .B2(n_716), .Y(n_712) );
OR2x2_ASAP7_75t_L g723 ( .A(n_520), .B(n_724), .Y(n_723) );
CKINVDCx16_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
OR2x2_ASAP7_75t_L g591 ( .A(n_521), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_521), .B(n_605), .Y(n_670) );
BUFx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx4_ASAP7_75t_L g562 ( .A(n_522), .Y(n_562) );
AND2x2_ASAP7_75t_L g628 ( .A(n_522), .B(n_593), .Y(n_628) );
AND3x2_ASAP7_75t_L g637 ( .A(n_522), .B(n_533), .C(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g563 ( .A(n_534), .B(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_534), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_534), .B(n_562), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
AND2x2_ASAP7_75t_L g558 ( .A(n_536), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g598 ( .A(n_536), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g616 ( .A(n_536), .B(n_548), .Y(n_616) );
AND2x2_ASAP7_75t_L g634 ( .A(n_536), .B(n_538), .Y(n_634) );
OR2x2_ASAP7_75t_L g648 ( .A(n_536), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g694 ( .A(n_536), .B(n_622), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_537), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_548), .Y(n_537) );
AND2x2_ASAP7_75t_L g595 ( .A(n_538), .B(n_573), .Y(n_595) );
OR2x2_ASAP7_75t_L g649 ( .A(n_538), .B(n_573), .Y(n_649) );
AND2x2_ASAP7_75t_L g702 ( .A(n_538), .B(n_559), .Y(n_702) );
INVx2_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
BUFx2_ASAP7_75t_L g600 ( .A(n_539), .Y(n_600) );
AND2x2_ASAP7_75t_L g622 ( .A(n_539), .B(n_548), .Y(n_622) );
INVx2_ASAP7_75t_L g559 ( .A(n_548), .Y(n_559) );
INVx1_ASAP7_75t_L g579 ( .A(n_548), .Y(n_579) );
AOI211xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_560), .B(n_565), .C(n_577), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_558), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g721 ( .A(n_558), .Y(n_721) );
AND2x2_ASAP7_75t_L g599 ( .A(n_559), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_562), .B(n_563), .Y(n_571) );
INVx1_ASAP7_75t_L g656 ( .A(n_562), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_562), .B(n_583), .Y(n_680) );
AND2x2_ASAP7_75t_L g696 ( .A(n_562), .B(n_610), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_563), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g587 ( .A(n_564), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_571), .B1(n_572), .B2(n_575), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_568), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_569), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g594 ( .A(n_570), .B(n_595), .Y(n_594) );
AOI221xp5_ASAP7_75t_SL g659 ( .A1(n_570), .A2(n_612), .B1(n_660), .B2(n_665), .C(n_667), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_570), .B(n_633), .Y(n_666) );
INVx1_ASAP7_75t_L g726 ( .A(n_572), .Y(n_726) );
BUFx3_ASAP7_75t_L g633 ( .A(n_573), .Y(n_633) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AOI21xp33_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_580), .B(n_581), .Y(n_577) );
INVx1_ASAP7_75t_L g642 ( .A(n_579), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_579), .B(n_633), .Y(n_686) );
INVx1_ASAP7_75t_L g643 ( .A(n_580), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_580), .B(n_633), .Y(n_644) );
INVxp67_ASAP7_75t_L g664 ( .A(n_582), .Y(n_664) );
AND2x2_ASAP7_75t_L g605 ( .A(n_583), .B(n_606), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_590), .B(n_594), .C(n_596), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_SL g619 ( .A(n_587), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_588), .B(n_619), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_588), .B(n_610), .Y(n_661) );
INVx2_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_591), .A2(n_597), .B1(n_601), .B2(n_603), .Y(n_596) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g612 ( .A(n_593), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g657 ( .A(n_593), .B(n_658), .Y(n_657) );
OAI21xp33_ASAP7_75t_L g660 ( .A1(n_595), .A2(n_661), .B(n_662), .Y(n_660) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
AOI221xp5_ASAP7_75t_L g607 ( .A1(n_599), .A2(n_608), .B1(n_611), .B2(n_612), .C(n_614), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_599), .B(n_633), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_599), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g715 ( .A(n_605), .Y(n_715) );
INVxp67_ASAP7_75t_L g638 ( .A(n_606), .Y(n_638) );
INVx1_ASAP7_75t_L g645 ( .A(n_608), .Y(n_645) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
AND2x2_ASAP7_75t_L g684 ( .A(n_609), .B(n_613), .Y(n_684) );
INVx1_ASAP7_75t_L g658 ( .A(n_613), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_613), .B(n_628), .Y(n_688) );
OAI32xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_617), .A3(n_619), .B1(n_620), .B2(n_621), .Y(n_614) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_SL g627 ( .A(n_622), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_622), .B(n_654), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_622), .B(n_683), .Y(n_714) );
NAND2x1p5_ASAP7_75t_L g722 ( .A(n_622), .B(n_633), .Y(n_722) );
NAND5xp2_ASAP7_75t_L g623 ( .A(n_624), .B(n_646), .C(n_659), .D(n_671), .E(n_672), .Y(n_623) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_628), .B1(n_629), .B2(n_631), .C(n_635), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp33_ASAP7_75t_SL g650 ( .A(n_630), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_633), .B(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_634), .A2(n_647), .B1(n_650), .B2(n_654), .Y(n_646) );
INVx2_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
OAI211xp5_ASAP7_75t_SL g641 ( .A1(n_637), .A2(n_642), .B(n_643), .C(n_644), .Y(n_641) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g669 ( .A(n_649), .Y(n_669) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_658), .B(n_707), .Y(n_717) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI222xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_675), .B1(n_677), .B2(n_681), .C1(n_684), .C2(n_685), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI221xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B1(n_691), .B2(n_693), .C(n_695), .Y(n_687) );
INVx1_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
OAI21xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B(n_700), .Y(n_695) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g707 ( .A(n_699), .Y(n_707) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_706), .B1(n_708), .B2(n_710), .C(n_712), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_722), .B(n_723), .C(n_725), .Y(n_718) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OAI21xp33_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B(n_728), .Y(n_725) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_731), .A2(n_734), .B1(n_735), .B2(n_736), .Y(n_733) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
endmodule