module real_jpeg_32302_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_0),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_0),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_1),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_1),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_1),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_1),
.B(n_352),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_1),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_1),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_1),
.B(n_447),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_2),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_2),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_2),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_2),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_2),
.B(n_189),
.Y(n_188)
);

NAND2xp33_ASAP7_75t_SL g209 ( 
.A(n_2),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_2),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_2),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_3),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_3),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_3),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_3),
.B(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_3),
.Y(n_171)
);

NAND2x1_ASAP7_75t_L g308 ( 
.A(n_3),
.B(n_85),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_3),
.B(n_354),
.Y(n_353)
);

NAND2x1_ASAP7_75t_L g412 ( 
.A(n_3),
.B(n_413),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_4),
.A2(n_19),
.B(n_477),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_4),
.B(n_478),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_5),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_5),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_5),
.Y(n_472)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_7),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_7),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_7),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_7),
.B(n_304),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_7),
.B(n_304),
.Y(n_309)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_7),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_7),
.B(n_427),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_7),
.B(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_8),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_8),
.Y(n_169)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_8),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_9),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_9),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_9),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_9),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_9),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_9),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_9),
.B(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_10),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_10),
.Y(n_193)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_10),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_11),
.Y(n_395)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_12),
.Y(n_109)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_12),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_13),
.B(n_92),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_13),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_13),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_13),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_13),
.B(n_287),
.Y(n_463)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_14),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_15),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_15),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_16),
.B(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_16),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_16),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_16),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_16),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_16),
.B(n_336),
.Y(n_335)
);

AND2x4_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_17),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_17),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_17),
.B(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_17),
.B(n_287),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_17),
.B(n_340),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_17),
.B(n_393),
.Y(n_392)
);

AND2x2_ASAP7_75t_SL g469 ( 
.A(n_17),
.B(n_470),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_431),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_368),
.B(n_429),
.Y(n_20)
);

NOR2xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_364),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_256),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_158),
.B(n_255),
.Y(n_23)
);

NOR2xp67_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_112),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_25),
.B(n_112),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_73),
.C(n_94),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_26),
.B(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_44),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_27),
.B(n_56),
.C(n_71),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_39),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_29),
.B(n_38),
.C(n_39),
.Y(n_119)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_32),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_33),
.A2(n_38),
.B1(n_467),
.B2(n_473),
.Y(n_466)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_43),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_56),
.B1(n_71),
.B2(n_72),
.Y(n_44)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_46),
.B(n_51),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_46),
.A2(n_47),
.B1(n_96),
.B2(n_97),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

MAJx2_ASAP7_75t_L g386 ( 
.A(n_47),
.B(n_97),
.C(n_326),
.Y(n_386)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_55),
.Y(n_139)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_55),
.Y(n_270)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_55),
.Y(n_355)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.C(n_66),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_57),
.B(n_66),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_61),
.Y(n_342)
);

XNOR2x2_ASAP7_75t_SL g243 ( 
.A(n_62),
.B(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_69),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_70),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_70),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_73),
.A2(n_74),
.B1(n_94),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_83),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_75),
.B(n_88),
.C(n_93),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

AO22x1_ASAP7_75t_SL g110 ( 
.A1(n_76),
.A2(n_80),
.B1(n_81),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_76),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_76),
.A2(n_111),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_76),
.B(n_282),
.C(n_286),
.Y(n_358)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_78),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_79),
.B(n_426),
.C(n_465),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_79),
.A2(n_80),
.B1(n_468),
.B2(n_469),
.Y(n_467)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22x1_ASAP7_75t_L g425 ( 
.A1(n_80),
.A2(n_81),
.B1(n_426),
.B2(n_428),
.Y(n_425)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_88),
.B1(n_89),
.B2(n_93),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_94),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_103),
.C(n_110),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_95),
.B(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_96),
.A2(n_97),
.B1(n_411),
.B2(n_412),
.Y(n_410)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_97),
.B(n_99),
.Y(n_185)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_97),
.Y(n_450)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_102),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_103),
.A2(n_104),
.B1(n_110),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_108),
.Y(n_222)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_108),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_109),
.Y(n_203)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_109),
.Y(n_276)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_110),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_134),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_114),
.B(n_134),
.C(n_259),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_115),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2x1_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_118),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_119),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_120),
.B(n_263),
.C(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_131),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_SL g293 ( 
.A(n_123),
.B(n_127),
.C(n_131),
.Y(n_293)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx8_ASAP7_75t_L g448 ( 
.A(n_126),
.Y(n_448)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_130),
.Y(n_352)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g310 ( 
.A(n_135),
.B(n_142),
.C(n_156),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_142),
.B1(n_156),
.B2(n_157),
.Y(n_136)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_140),
.B(n_141),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_140),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_141),
.B(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_141),
.B(n_271),
.C(n_277),
.Y(n_348)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

XNOR2x1_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_149),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_144),
.B(n_152),
.C(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_148),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_150),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_150),
.B(n_410),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_150),
.B(n_412),
.C(n_450),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_154),
.B(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI21x1_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_249),
.B(n_254),
.Y(n_158)
);

OAI21x1_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_237),
.B(n_248),
.Y(n_159)
);

AOI21x1_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_206),
.B(n_236),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_180),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g236 ( 
.A(n_162),
.B(n_180),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_174),
.C(n_177),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_163),
.A2(n_164),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_170),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_174),
.A2(n_177),
.B1(n_178),
.B2(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_174),
.Y(n_216)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_186),
.B1(n_204),
.B2(n_205),
.Y(n_180)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_182),
.B(n_185),
.C(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_194),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_188),
.B(n_195),
.C(n_199),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

OAI21x1_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_217),
.B(n_235),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_213),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_211),
.Y(n_219)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_223),
.B(n_234),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_220),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_228),
.Y(n_301)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_240),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_245),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_243),
.C(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

NOR2xp67_ASAP7_75t_SL g254 ( 
.A(n_250),
.B(n_253),
.Y(n_254)
);

NOR2x1_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_312),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_258),
.B(n_260),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_289),
.Y(n_260)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_261),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_262),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_278),
.Y(n_265)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_266),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_271),
.B1(n_272),
.B2(n_277),
.Y(n_267)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_278),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_285),
.B2(n_288),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_284),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_310),
.B2(n_311),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_296),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_293),
.B(n_294),
.C(n_297),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_302),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_298),
.B(n_308),
.C(n_344),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_303),
.A2(n_309),
.B1(n_462),
.B2(n_463),
.Y(n_461)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx5_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_306),
.Y(n_424)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_309),
.Y(n_344)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_310),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_314),
.C(n_315),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_312),
.A2(n_366),
.B(n_367),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_313),
.B(n_316),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_321),
.Y(n_316)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_317),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.C(n_320),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_345),
.B1(n_346),
.B2(n_360),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_343),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_330),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_324),
.B(n_361),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_324),
.B(n_330),
.C(n_363),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_330),
.A2(n_343),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_330),
.Y(n_362)
);

XOR2x2_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_339),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_334),
.B1(n_335),
.B2(n_338),
.Y(n_331)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_332),
.Y(n_338)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_335),
.Y(n_418)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_338),
.B(n_339),
.C(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_341),
.Y(n_427)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_343),
.Y(n_363)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_346),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_359),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

HB1xp67_ASAP7_75t_SL g405 ( 
.A(n_348),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_349),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_358),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_353),
.B1(n_356),
.B2(n_357),
.Y(n_350)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_351),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_353),
.Y(n_357)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_355),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_356),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_357),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_358),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_359),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_360),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_375),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_371),
.B(n_377),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.C(n_374),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_377),
.Y(n_376)
);

XNOR2x1_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_402),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_379),
.B(n_407),
.C(n_435),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_399),
.B1(n_400),
.B2(n_401),
.Y(n_379)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_380),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_385),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_381),
.B(n_399),
.C(n_438),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.C(n_384),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_385),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_386),
.A2(n_452),
.B(n_453),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_392),
.B1(n_396),
.B2(n_398),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_390),
.Y(n_397)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_392),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_392),
.A2(n_398),
.B1(n_445),
.B2(n_446),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_392),
.B(n_396),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_392),
.B(n_396),
.Y(n_453)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2x1_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_407),
.Y(n_402)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_403),
.Y(n_435)
);

MAJx2_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.C(n_406),
.Y(n_403)
);

XOR2x2_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_416),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_409),
.B(n_417),
.C(n_419),
.Y(n_454)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_419),
.Y(n_416)
);

XNOR2x1_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_425),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_420),
.Y(n_465)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_426),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_475),
.Y(n_431)
);

INVxp33_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_436),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_434),
.B(n_436),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_439),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_441),
.B1(n_455),
.B2(n_474),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_454),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_451),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_449),
.Y(n_443)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_455),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_466),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_464),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_461),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_467),
.Y(n_473)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);


endmodule