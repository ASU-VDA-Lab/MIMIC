module fake_ariane_1362_n_1762 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1762);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1762;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx2_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_98),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_115),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_51),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_4),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_37),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_74),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_155),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_14),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_86),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_44),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_92),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_151),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_88),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_134),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_27),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_85),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_96),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_62),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_65),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_30),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_57),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_105),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_13),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_109),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_123),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_121),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_131),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_9),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_45),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_46),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_0),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_64),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_17),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_89),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_136),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_28),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_2),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_8),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_19),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_55),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_52),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_12),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_0),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_25),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_9),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_152),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_72),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_70),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_112),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_93),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_76),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_139),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_29),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_41),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_15),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_132),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_17),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_68),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_23),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_42),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_71),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_154),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_146),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_100),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_128),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_101),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_81),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_153),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_56),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_145),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_84),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_18),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_80),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_12),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_15),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_91),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_77),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_13),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_79),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_58),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_90),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_78),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_28),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_16),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_38),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_1),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_35),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_111),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_144),
.Y(n_251)
);

CKINVDCx11_ASAP7_75t_R g252 ( 
.A(n_6),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_87),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_108),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_110),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_82),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_34),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_46),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_26),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_36),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_126),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_61),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_24),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_40),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_18),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_29),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_33),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_133),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_6),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_113),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_35),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_5),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_116),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_16),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_75),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_118),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_106),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_37),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_43),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_25),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_142),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_33),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_44),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_50),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_53),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_43),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_66),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_67),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_47),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_48),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_24),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_83),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_3),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_38),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_40),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_22),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_8),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_104),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_114),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_14),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_95),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_45),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_60),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_125),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_7),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_122),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_148),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_135),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_69),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_201),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_252),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_202),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_201),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_174),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_178),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_182),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_191),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_196),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_206),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_207),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_215),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_215),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_270),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_220),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_309),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_215),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_215),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_215),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_156),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_217),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_266),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_266),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_175),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_222),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_234),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g336 ( 
.A(n_212),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_285),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_217),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_266),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_231),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_236),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_237),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_245),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_280),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_246),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_257),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_266),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_301),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_260),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_269),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_266),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_264),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_286),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_200),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_272),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_295),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_200),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_216),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_280),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_216),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_285),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_285),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_158),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_158),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_249),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_159),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_161),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_249),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_296),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_296),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_302),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_294),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_302),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_305),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_177),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_159),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_177),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_166),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_225),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_221),
.Y(n_380)
);

INVxp33_ASAP7_75t_SL g381 ( 
.A(n_161),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_221),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_170),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_221),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_367),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_314),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_325),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_315),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_350),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_351),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_337),
.B(n_170),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_321),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_318),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_322),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_322),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_326),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_326),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_310),
.B(n_287),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_327),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_313),
.B(n_287),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_336),
.A2(n_162),
.B1(n_300),
.B2(n_297),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_327),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_353),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_328),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_339),
.B(n_157),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_328),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_375),
.B(n_163),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_331),
.Y(n_411)
);

NOR2x1_ASAP7_75t_L g412 ( 
.A(n_383),
.B(n_375),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_336),
.B(n_307),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_363),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_332),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_347),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_383),
.Y(n_418)
);

OAI21x1_ASAP7_75t_L g419 ( 
.A1(n_347),
.A2(n_307),
.B(n_165),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_354),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_354),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_357),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_316),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_363),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_358),
.Y(n_425)
);

AND2x6_ASAP7_75t_L g426 ( 
.A(n_317),
.B(n_307),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_360),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_325),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_380),
.B(n_179),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_319),
.B(n_164),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_365),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_368),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_369),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_370),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_320),
.B(n_168),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_371),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_372),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_373),
.B(n_279),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_334),
.B(n_173),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_335),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_341),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_342),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_343),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_345),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_346),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_364),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_349),
.B(n_352),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_355),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_312),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_337),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_356),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_330),
.B(n_180),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_324),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_450),
.B(n_364),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_398),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_409),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_393),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_418),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_393),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_396),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_393),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_398),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_396),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_393),
.Y(n_464)
);

BUFx10_ASAP7_75t_L g465 ( 
.A(n_413),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_399),
.Y(n_466)
);

INVx8_ASAP7_75t_L g467 ( 
.A(n_426),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_393),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_397),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_450),
.B(n_366),
.Y(n_470)
);

CKINVDCx6p67_ASAP7_75t_R g471 ( 
.A(n_449),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_397),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_397),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_390),
.Y(n_474)
);

BUFx4f_ASAP7_75t_L g475 ( 
.A(n_426),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_413),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_438),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_450),
.B(n_366),
.Y(n_478)
);

BUFx4f_ASAP7_75t_L g479 ( 
.A(n_426),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_397),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_397),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_396),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_399),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_415),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_414),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_415),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_415),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_410),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_423),
.B(n_448),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_418),
.Y(n_490)
);

AOI21x1_ASAP7_75t_L g491 ( 
.A1(n_419),
.A2(n_203),
.B(n_194),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_396),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_415),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_392),
.A2(n_379),
.B1(n_381),
.B2(n_329),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_387),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_438),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_425),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_415),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_450),
.B(n_376),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_423),
.B(n_361),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_410),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_409),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_450),
.B(n_376),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_392),
.A2(n_381),
.B1(n_329),
.B2(n_333),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_446),
.B(n_323),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_411),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_388),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_391),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_391),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_396),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_446),
.B(n_378),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_411),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_391),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_416),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_391),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_403),
.A2(n_333),
.B1(n_377),
.B2(n_382),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_423),
.B(n_361),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_440),
.B(n_384),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_416),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_417),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_438),
.B(n_378),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_388),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_440),
.B(n_441),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_390),
.B(n_374),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_396),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_388),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_426),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_428),
.Y(n_528)
);

AO22x2_ASAP7_75t_L g529 ( 
.A1(n_403),
.A2(n_278),
.B1(n_359),
.B2(n_344),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_414),
.B(n_362),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_425),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_417),
.Y(n_532)
);

NOR2x1p5_ASAP7_75t_L g533 ( 
.A(n_448),
.B(n_362),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_417),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_417),
.Y(n_535)
);

NOR2x1p5_ASAP7_75t_L g536 ( 
.A(n_452),
.B(n_162),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_429),
.A2(n_282),
.B1(n_283),
.B2(n_291),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_394),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_396),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_429),
.B(n_338),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_407),
.B(n_160),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_394),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_394),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_407),
.B(n_166),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_440),
.B(n_418),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_401),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_401),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_401),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_440),
.B(n_171),
.Y(n_549)
);

NOR3xp33_ASAP7_75t_L g550 ( 
.A(n_385),
.B(n_169),
.C(n_167),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_396),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_404),
.Y(n_552)
);

INVx5_ASAP7_75t_L g553 ( 
.A(n_426),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_R g554 ( 
.A(n_449),
.B(n_389),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_404),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_408),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_408),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_424),
.B(n_171),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_385),
.B(n_340),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_424),
.B(n_172),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_406),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_406),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_428),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_406),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_425),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_406),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_440),
.B(n_172),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_408),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_400),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_406),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_428),
.B(n_181),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_395),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_406),
.Y(n_573)
);

INVxp67_ASAP7_75t_SL g574 ( 
.A(n_447),
.Y(n_574)
);

INVx6_ASAP7_75t_L g575 ( 
.A(n_425),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_420),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_418),
.B(n_181),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_452),
.B(n_183),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_420),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_420),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_406),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_425),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_426),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_406),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_400),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_420),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_426),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_421),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_453),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_421),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_386),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_386),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_421),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_386),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_386),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_426),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_386),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_426),
.B(n_183),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_421),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_L g600 ( 
.A(n_447),
.B(n_169),
.C(n_167),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_425),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_L g602 ( 
.A(n_442),
.B(n_185),
.C(n_176),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_458),
.Y(n_603)
);

BUFx5_ASAP7_75t_L g604 ( 
.A(n_583),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_474),
.B(n_400),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_465),
.B(n_442),
.Y(n_606)
);

BUFx4_ASAP7_75t_L g607 ( 
.A(n_471),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_518),
.A2(n_426),
.B1(n_445),
.B2(n_451),
.Y(n_608)
);

O2A1O1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_574),
.A2(n_451),
.B(n_445),
.C(n_430),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_465),
.B(n_430),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_507),
.B(n_402),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_455),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_508),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_508),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_465),
.B(n_435),
.Y(n_615)
);

AND2x6_ASAP7_75t_SL g616 ( 
.A(n_559),
.B(n_311),
.Y(n_616)
);

NOR3xp33_ASAP7_75t_L g617 ( 
.A(n_521),
.B(n_185),
.C(n_176),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_455),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_545),
.A2(n_419),
.B(n_435),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_462),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_465),
.B(n_439),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_456),
.B(n_402),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_508),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_502),
.B(n_402),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_475),
.B(n_419),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_529),
.A2(n_444),
.B1(n_443),
.B2(n_441),
.Y(n_626)
);

O2A1O1Ixp5_ASAP7_75t_L g627 ( 
.A1(n_599),
.A2(n_439),
.B(n_443),
.C(n_441),
.Y(n_627)
);

NOR2xp67_ASAP7_75t_L g628 ( 
.A(n_505),
.B(n_443),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_489),
.A2(n_444),
.B(n_251),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_SL g630 ( 
.A(n_471),
.B(n_348),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_467),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_507),
.B(n_444),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_509),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_477),
.B(n_431),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_541),
.B(n_412),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_462),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_466),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_509),
.Y(n_638)
);

BUFx6f_ASAP7_75t_SL g639 ( 
.A(n_476),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_466),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_544),
.B(n_412),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_476),
.B(n_431),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_483),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_569),
.B(n_422),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_569),
.B(n_422),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_537),
.A2(n_282),
.B1(n_283),
.B2(n_291),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_585),
.B(n_422),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_476),
.B(n_184),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_476),
.B(n_184),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_585),
.B(n_422),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_509),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_540),
.B(n_432),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_500),
.B(n_432),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_477),
.B(n_496),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_495),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_513),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_589),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_496),
.B(n_433),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_518),
.B(n_433),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_483),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_522),
.B(n_405),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_523),
.B(n_434),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_523),
.B(n_434),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_522),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_513),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_549),
.A2(n_567),
.B(n_517),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_537),
.B(n_577),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_572),
.Y(n_668)
);

O2A1O1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_488),
.A2(n_251),
.B(n_179),
.C(n_239),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_526),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_511),
.B(n_425),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_485),
.B(n_186),
.Y(n_672)
);

BUFx5_ASAP7_75t_L g673 ( 
.A(n_583),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_454),
.B(n_425),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_526),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_475),
.B(n_186),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_488),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_L g678 ( 
.A(n_467),
.B(n_187),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_470),
.B(n_427),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_458),
.B(n_427),
.Y(n_680)
);

BUFx6f_ASAP7_75t_SL g681 ( 
.A(n_554),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_501),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_458),
.B(n_427),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_501),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_490),
.B(n_427),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_478),
.B(n_427),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_528),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_513),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_499),
.B(n_427),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_503),
.B(n_427),
.Y(n_690)
);

BUFx6f_ASAP7_75t_SL g691 ( 
.A(n_524),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_475),
.B(n_187),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_490),
.B(n_427),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_506),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_SL g695 ( 
.A(n_528),
.B(n_405),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_506),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g697 ( 
.A(n_563),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_524),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_490),
.B(n_436),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_504),
.B(n_475),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_578),
.B(n_436),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_467),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_576),
.B(n_436),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_512),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_576),
.B(n_436),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_579),
.B(n_580),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_512),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_583),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_479),
.B(n_233),
.Y(n_709)
);

NAND2x1p5_ASAP7_75t_L g710 ( 
.A(n_587),
.B(n_436),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_479),
.B(n_233),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_515),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_494),
.A2(n_293),
.B1(n_297),
.B2(n_300),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_533),
.A2(n_288),
.B1(n_277),
.B2(n_308),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_579),
.B(n_436),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_580),
.B(n_436),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_587),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_516),
.B(n_530),
.Y(n_718)
);

NOR2x1p5_ASAP7_75t_L g719 ( 
.A(n_600),
.B(n_293),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_586),
.B(n_436),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_514),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_479),
.B(n_277),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_515),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_514),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_558),
.B(n_190),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_586),
.B(n_281),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_467),
.B(n_281),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_529),
.A2(n_279),
.B1(n_228),
.B2(n_230),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_479),
.B(n_288),
.Y(n_729)
);

INVxp33_ASAP7_75t_L g730 ( 
.A(n_550),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_519),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_519),
.Y(n_732)
);

NOR3xp33_ASAP7_75t_L g733 ( 
.A(n_571),
.B(n_247),
.C(n_240),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_467),
.B(n_289),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_515),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_588),
.B(n_289),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_534),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_560),
.B(n_192),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_588),
.B(n_292),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_533),
.A2(n_205),
.B1(n_204),
.B2(n_199),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_602),
.B(n_271),
.C(n_258),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_590),
.B(n_292),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_587),
.B(n_298),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_593),
.B(n_298),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_527),
.B(n_299),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_527),
.B(n_299),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_534),
.Y(n_747)
);

BUFx6f_ASAP7_75t_SL g748 ( 
.A(n_593),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_534),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_538),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_538),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_527),
.B(n_306),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_536),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_543),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_536),
.B(n_437),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_598),
.A2(n_306),
.B1(n_308),
.B2(n_244),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_542),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_480),
.B(n_481),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_527),
.B(n_193),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_457),
.A2(n_242),
.B(n_304),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_480),
.B(n_195),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_529),
.A2(n_464),
.B1(n_473),
.B2(n_472),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_527),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_529),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_599),
.B(n_437),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_480),
.B(n_481),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_481),
.B(n_198),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_591),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_527),
.B(n_211),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_542),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_668),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_661),
.B(n_595),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_612),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_618),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_610),
.B(n_484),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_613),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_610),
.B(n_484),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_614),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_611),
.B(n_279),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_670),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_615),
.B(n_484),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_615),
.B(n_621),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_728),
.A2(n_548),
.B1(n_557),
.B2(n_568),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_623),
.Y(n_784)
);

OR2x2_ASAP7_75t_SL g785 ( 
.A(n_718),
.B(n_235),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_728),
.A2(n_546),
.B1(n_547),
.B2(n_548),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_604),
.B(n_497),
.Y(n_787)
);

AO22x1_ASAP7_75t_L g788 ( 
.A1(n_655),
.A2(n_657),
.B1(n_698),
.B2(n_730),
.Y(n_788)
);

OAI22xp33_ASAP7_75t_L g789 ( 
.A1(n_667),
.A2(n_259),
.B1(n_219),
.B2(n_274),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_R g790 ( 
.A(n_681),
.B(n_553),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_670),
.Y(n_791)
);

AND3x2_ASAP7_75t_SL g792 ( 
.A(n_616),
.B(n_555),
.C(n_552),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_708),
.Y(n_793)
);

OAI22xp33_ASAP7_75t_L g794 ( 
.A1(n_659),
.A2(n_248),
.B1(n_267),
.B2(n_263),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_764),
.A2(n_547),
.B1(n_557),
.B2(n_556),
.Y(n_795)
);

INVx5_ASAP7_75t_L g796 ( 
.A(n_631),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_633),
.Y(n_797)
);

NOR2x1p5_ASAP7_75t_L g798 ( 
.A(n_607),
.B(n_265),
.Y(n_798)
);

NOR2x1_ASAP7_75t_R g799 ( 
.A(n_664),
.B(n_188),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_621),
.B(n_486),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_675),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_638),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_606),
.B(n_486),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_632),
.B(n_553),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_SL g805 ( 
.A(n_681),
.B(n_553),
.Y(n_805)
);

OR2x6_ASAP7_75t_L g806 ( 
.A(n_687),
.B(n_552),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_765),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_606),
.A2(n_498),
.B1(n_493),
.B2(n_487),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_605),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_651),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_697),
.B(n_595),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_603),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_642),
.A2(n_457),
.B1(n_459),
.B2(n_461),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_603),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_708),
.Y(n_815)
);

NOR2x2_ASAP7_75t_L g816 ( 
.A(n_695),
.B(n_459),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_697),
.B(n_755),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_622),
.B(n_624),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_604),
.B(n_497),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_719),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_753),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_653),
.B(n_487),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_717),
.Y(n_823)
);

OR2x6_ASAP7_75t_L g824 ( 
.A(n_634),
.B(n_555),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_620),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_634),
.B(n_553),
.Y(n_826)
);

INVx5_ASAP7_75t_L g827 ( 
.A(n_631),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_636),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_604),
.B(n_497),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_654),
.Y(n_830)
);

AND3x1_ASAP7_75t_L g831 ( 
.A(n_617),
.B(n_591),
.C(n_594),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_604),
.B(n_497),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_717),
.Y(n_833)
);

O2A1O1Ixp5_ASAP7_75t_L g834 ( 
.A1(n_666),
.A2(n_491),
.B(n_520),
.C(n_532),
.Y(n_834)
);

INVx4_ASAP7_75t_L g835 ( 
.A(n_631),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_631),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_672),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_642),
.A2(n_493),
.B1(n_498),
.B2(n_487),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_637),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_652),
.B(n_493),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_764),
.A2(n_556),
.B1(n_546),
.B2(n_568),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_628),
.B(n_635),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_640),
.A2(n_498),
.B1(n_469),
.B2(n_473),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_658),
.B(n_662),
.Y(n_844)
);

NAND3xp33_ASAP7_75t_SL g845 ( 
.A(n_733),
.B(n_232),
.C(n_214),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_626),
.A2(n_535),
.B1(n_532),
.B2(n_520),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_761),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_641),
.B(n_461),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_604),
.B(n_497),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_643),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_646),
.B(n_597),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_604),
.B(n_497),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_663),
.B(n_464),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_660),
.B(n_677),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_682),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_684),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_673),
.B(n_531),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_694),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_673),
.B(n_531),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_762),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_696),
.B(n_704),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_702),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_707),
.B(n_468),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_656),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_691),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_673),
.B(n_702),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_721),
.A2(n_724),
.B1(n_732),
.B2(n_731),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_673),
.B(n_531),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_750),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_626),
.B(n_468),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_751),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_630),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_702),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_639),
.B(n_469),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_644),
.B(n_472),
.Y(n_875)
);

OR2x2_ASAP7_75t_SL g876 ( 
.A(n_691),
.B(n_241),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_767),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_645),
.B(n_535),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_647),
.B(n_597),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_757),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_665),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_650),
.B(n_591),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_725),
.B(n_592),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_725),
.B(n_592),
.Y(n_884)
);

OR2x6_ASAP7_75t_L g885 ( 
.A(n_702),
.B(n_592),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_688),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_763),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_770),
.Y(n_888)
);

INVxp67_ASAP7_75t_SL g889 ( 
.A(n_673),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_738),
.B(n_594),
.Y(n_890)
);

OR2x2_ASAP7_75t_SL g891 ( 
.A(n_741),
.B(n_250),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_673),
.B(n_531),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_648),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_712),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_639),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_723),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_748),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_713),
.B(n_594),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_738),
.B(n_460),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_754),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_735),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_R g902 ( 
.A(n_678),
.B(n_553),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_609),
.B(n_460),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_768),
.B(n_460),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_737),
.Y(n_905)
);

OR2x6_ASAP7_75t_L g906 ( 
.A(n_700),
.B(n_575),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_671),
.Y(n_907)
);

INVx8_ASAP7_75t_L g908 ( 
.A(n_748),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_768),
.B(n_460),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_747),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_671),
.B(n_714),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_726),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_758),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_733),
.B(n_617),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_649),
.A2(n_575),
.B1(n_463),
.B2(n_510),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_608),
.B(n_531),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_706),
.B(n_463),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_743),
.B(n_463),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_766),
.A2(n_562),
.B(n_482),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_627),
.A2(n_566),
.B(n_551),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_701),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_736),
.B(n_463),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_763),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_749),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_743),
.A2(n_553),
.B1(n_596),
.B2(n_575),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_710),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_701),
.A2(n_596),
.B1(n_575),
.B2(n_584),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_703),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_710),
.B(n_531),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_705),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_756),
.A2(n_596),
.B1(n_551),
.B2(n_584),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_739),
.B(n_482),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_740),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_769),
.B(n_596),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_742),
.B(n_482),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_680),
.Y(n_936)
);

BUFx4f_ASAP7_75t_L g937 ( 
.A(n_669),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_715),
.Y(n_938)
);

AND3x1_ASAP7_75t_L g939 ( 
.A(n_744),
.B(n_539),
.C(n_562),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_716),
.B(n_482),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_720),
.Y(n_941)
);

CKINVDCx11_ASAP7_75t_R g942 ( 
.A(n_627),
.Y(n_942)
);

NOR2x1p5_ASAP7_75t_L g943 ( 
.A(n_683),
.B(n_492),
.Y(n_943)
);

O2A1O1Ixp5_ASAP7_75t_L g944 ( 
.A1(n_629),
.A2(n_619),
.B(n_686),
.C(n_679),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_769),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_685),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_693),
.Y(n_947)
);

AND2x2_ASAP7_75t_SL g948 ( 
.A(n_727),
.B(n_253),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_674),
.B(n_679),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_674),
.B(n_492),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_686),
.Y(n_951)
);

BUFx12f_ASAP7_75t_L g952 ( 
.A(n_760),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_699),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_745),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_676),
.A2(n_596),
.B1(n_573),
.B2(n_584),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_676),
.A2(n_596),
.B1(n_570),
.B2(n_566),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_773),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_771),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_782),
.B(n_689),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_836),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_889),
.A2(n_625),
.B(n_734),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_912),
.B(n_692),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_818),
.B(n_844),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_911),
.A2(n_690),
.B1(n_689),
.B2(n_709),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_780),
.B(n_791),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_801),
.B(n_692),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_791),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_933),
.A2(n_690),
.B(n_709),
.C(n_722),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_807),
.B(n_826),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_854),
.A2(n_711),
.B1(n_729),
.B2(n_625),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_907),
.A2(n_745),
.B(n_746),
.C(n_573),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_907),
.A2(n_746),
.B(n_551),
.C(n_573),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_951),
.A2(n_570),
.B(n_564),
.C(n_566),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_889),
.A2(n_759),
.B(n_752),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_881),
.Y(n_975)
);

O2A1O1Ixp5_ASAP7_75t_L g976 ( 
.A1(n_944),
.A2(n_491),
.B(n_564),
.C(n_581),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_826),
.B(n_565),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_822),
.A2(n_803),
.B(n_777),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_908),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_774),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_861),
.A2(n_539),
.B1(n_492),
.B2(n_525),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_809),
.B(n_510),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_775),
.A2(n_800),
.B(n_781),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_835),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_881),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_817),
.B(n_510),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_886),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_840),
.A2(n_561),
.B(n_510),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_951),
.A2(n_564),
.B(n_581),
.C(n_570),
.Y(n_989)
);

OA22x2_ASAP7_75t_L g990 ( 
.A1(n_809),
.A2(n_290),
.B1(n_261),
.B2(n_275),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_825),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_917),
.A2(n_562),
.B(n_525),
.Y(n_992)
);

AND2x6_ASAP7_75t_SL g993 ( 
.A(n_914),
.B(n_284),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_807),
.Y(n_994)
);

NOR3xp33_ASAP7_75t_SL g995 ( 
.A(n_845),
.B(n_213),
.C(n_210),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_865),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_908),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_816),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_897),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_895),
.Y(n_1000)
);

OAI21xp33_ASAP7_75t_SL g1001 ( 
.A1(n_948),
.A2(n_581),
.B(n_539),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_828),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_824),
.Y(n_1003)
);

NOR3xp33_ASAP7_75t_L g1004 ( 
.A(n_789),
.B(n_788),
.C(n_914),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_824),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_804),
.B(n_565),
.Y(n_1006)
);

OAI22x1_ASAP7_75t_L g1007 ( 
.A1(n_872),
.A2(n_209),
.B1(n_208),
.B2(n_197),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_830),
.B(n_525),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_804),
.B(n_565),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_847),
.B(n_525),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_779),
.B(n_561),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_787),
.A2(n_562),
.B(n_561),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_772),
.Y(n_1013)
);

AOI21x1_ASAP7_75t_L g1014 ( 
.A1(n_916),
.A2(n_601),
.B(n_582),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_948),
.B(n_937),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_787),
.A2(n_561),
.B(n_582),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_860),
.A2(n_601),
.B1(n_582),
.B2(n_565),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_839),
.B(n_850),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_789),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_855),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_921),
.A2(n_867),
.B1(n_856),
.B2(n_858),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_913),
.B(n_601),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_921),
.A2(n_601),
.B1(n_582),
.B2(n_565),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_869),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_937),
.B(n_601),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_886),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_944),
.A2(n_243),
.B(n_276),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_871),
.A2(n_582),
.B1(n_238),
.B2(n_273),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_SL g1029 ( 
.A(n_872),
.B(n_229),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_880),
.Y(n_1030)
);

OAI21xp33_ASAP7_75t_SL g1031 ( 
.A1(n_888),
.A2(n_4),
.B(n_5),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_900),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_794),
.B(n_7),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_837),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_851),
.A2(n_227),
.B1(n_268),
.B2(n_262),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_819),
.A2(n_226),
.B(n_256),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_877),
.B(n_10),
.Y(n_1037)
);

NAND2x1_ASAP7_75t_L g1038 ( 
.A(n_835),
.B(n_303),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_796),
.B(n_255),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_796),
.B(n_254),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_785),
.B(n_10),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_836),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_790),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_SL g1044 ( 
.A1(n_920),
.A2(n_11),
.B(n_19),
.C(n_20),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_SL g1045 ( 
.A1(n_874),
.A2(n_11),
.B(n_20),
.C(n_21),
.Y(n_1045)
);

NAND2x1p5_ASAP7_75t_L g1046 ( 
.A(n_796),
.B(n_303),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_873),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_790),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_873),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_824),
.B(n_21),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_776),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_778),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_848),
.A2(n_224),
.B(n_223),
.C(n_218),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_842),
.B(n_22),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_806),
.B(n_23),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_794),
.B(n_811),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_806),
.A2(n_189),
.B1(n_303),
.B2(n_30),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_813),
.A2(n_303),
.B1(n_27),
.B2(n_31),
.Y(n_1058)
);

AOI221xp5_ASAP7_75t_L g1059 ( 
.A1(n_820),
.A2(n_303),
.B1(n_31),
.B2(n_32),
.C(n_34),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_796),
.B(n_26),
.Y(n_1060)
);

AO21x1_ASAP7_75t_L g1061 ( 
.A1(n_949),
.A2(n_102),
.B(n_141),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_795),
.B(n_32),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_R g1063 ( 
.A(n_805),
.B(n_150),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_795),
.B(n_841),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_784),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_806),
.B(n_36),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_827),
.B(n_39),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_926),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_798),
.B(n_39),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_797),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_827),
.B(n_41),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_833),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_926),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_834),
.A2(n_848),
.B(n_838),
.Y(n_1074)
);

NOR2x1_ASAP7_75t_L g1075 ( 
.A(n_874),
.B(n_812),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_819),
.A2(n_107),
.B(n_49),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_924),
.Y(n_1077)
);

CKINVDCx6p67_ASAP7_75t_R g1078 ( 
.A(n_827),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_834),
.A2(n_117),
.B(n_54),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_893),
.B(n_42),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_793),
.B(n_59),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_821),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_793),
.B(n_63),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_841),
.B(n_928),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_876),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_831),
.B(n_73),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_883),
.A2(n_94),
.B(n_97),
.C(n_120),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_802),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_930),
.B(n_124),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_829),
.A2(n_127),
.B(n_129),
.Y(n_1090)
);

XOR2x2_ASAP7_75t_L g1091 ( 
.A(n_792),
.B(n_130),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_899),
.A2(n_137),
.B(n_140),
.C(n_884),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_SL g1093 ( 
.A1(n_918),
.A2(n_922),
.B(n_935),
.C(n_932),
.Y(n_1093)
);

NAND3xp33_ASAP7_75t_SL g1094 ( 
.A(n_890),
.B(n_898),
.C(n_783),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_891),
.B(n_870),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_853),
.A2(n_863),
.B1(n_814),
.B2(n_812),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_942),
.A2(n_941),
.B1(n_938),
.B2(n_783),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_815),
.B(n_823),
.Y(n_1098)
);

NAND3xp33_ASAP7_75t_SL g1099 ( 
.A(n_786),
.B(n_915),
.C(n_799),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_810),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_942),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_864),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_996),
.Y(n_1103)
);

AO22x2_ASAP7_75t_L g1104 ( 
.A1(n_1101),
.A2(n_792),
.B1(n_954),
.B2(n_953),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_978),
.A2(n_859),
.B(n_852),
.Y(n_1105)
);

NAND3xp33_ASAP7_75t_L g1106 ( 
.A(n_1004),
.B(n_939),
.C(n_918),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_963),
.A2(n_829),
.B(n_849),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1014),
.A2(n_859),
.B(n_892),
.Y(n_1108)
);

AO21x2_ASAP7_75t_L g1109 ( 
.A1(n_1074),
.A2(n_916),
.B(n_849),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_967),
.B(n_786),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1013),
.B(n_901),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_1078),
.Y(n_1112)
);

AOI21x1_ASAP7_75t_SL g1113 ( 
.A1(n_1033),
.A2(n_903),
.B(n_940),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_964),
.A2(n_950),
.B(n_808),
.Y(n_1114)
);

AO31x2_ASAP7_75t_L g1115 ( 
.A1(n_983),
.A2(n_946),
.A3(n_843),
.B(n_947),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_960),
.Y(n_1116)
);

OAI21xp33_ASAP7_75t_L g1117 ( 
.A1(n_1004),
.A2(n_875),
.B(n_882),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_965),
.B(n_896),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_958),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_965),
.B(n_894),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_994),
.B(n_905),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_976),
.A2(n_832),
.B(n_857),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_1082),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1054),
.A2(n_931),
.B(n_945),
.C(n_943),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_976),
.A2(n_892),
.B(n_868),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_959),
.A2(n_919),
.B(n_878),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1054),
.A2(n_931),
.B(n_815),
.C(n_823),
.Y(n_1127)
);

AOI221xp5_ASAP7_75t_SL g1128 ( 
.A1(n_1019),
.A2(n_909),
.B1(n_904),
.B2(n_879),
.C(n_846),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_969),
.B(n_827),
.Y(n_1129)
);

CKINVDCx20_ASAP7_75t_R g1130 ( 
.A(n_1000),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_961),
.A2(n_832),
.B(n_868),
.Y(n_1131)
);

OAI21xp33_ASAP7_75t_L g1132 ( 
.A1(n_1056),
.A2(n_1062),
.B(n_1057),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_968),
.A2(n_929),
.B(n_955),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_962),
.B(n_910),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1064),
.A2(n_846),
.B1(n_814),
.B2(n_927),
.Y(n_1135)
);

NAND2xp33_ASAP7_75t_R g1136 ( 
.A(n_1063),
.B(n_902),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1079),
.A2(n_852),
.B(n_857),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_962),
.B(n_1095),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_994),
.B(n_833),
.Y(n_1139)
);

INVx4_ASAP7_75t_SL g1140 ( 
.A(n_960),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_1041),
.B(n_906),
.C(n_955),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_957),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_1034),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_960),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_969),
.B(n_998),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1005),
.B(n_885),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1016),
.A2(n_866),
.B(n_929),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_999),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1021),
.A2(n_927),
.B1(n_885),
.B2(n_956),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1012),
.A2(n_866),
.B(n_936),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1018),
.B(n_936),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1001),
.A2(n_956),
.B(n_906),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_960),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1041),
.A2(n_1015),
.B(n_1037),
.C(n_1099),
.Y(n_1154)
);

AOI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1025),
.A2(n_906),
.B(n_885),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1093),
.A2(n_836),
.B(n_862),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1093),
.A2(n_1023),
.B(n_970),
.Y(n_1157)
);

AOI221x1_ASAP7_75t_L g1158 ( 
.A1(n_1058),
.A2(n_862),
.B1(n_934),
.B2(n_923),
.C(n_887),
.Y(n_1158)
);

OA21x2_ASAP7_75t_L g1159 ( 
.A1(n_971),
.A2(n_972),
.B(n_1027),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_986),
.B(n_952),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_992),
.A2(n_925),
.B(n_902),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_973),
.A2(n_925),
.B(n_934),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_980),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1097),
.A2(n_862),
.B1(n_1050),
.B2(n_1017),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1097),
.A2(n_986),
.B1(n_1011),
.B2(n_1017),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_988),
.A2(n_974),
.B(n_1096),
.Y(n_1166)
);

AOI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1084),
.A2(n_1089),
.B(n_1061),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1050),
.B(n_1055),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_991),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1092),
.A2(n_1022),
.B(n_1094),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_981),
.A2(n_1081),
.B(n_1083),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1046),
.A2(n_1076),
.B(n_1090),
.Y(n_1172)
);

OAI22x1_ASAP7_75t_L g1173 ( 
.A1(n_993),
.A2(n_1037),
.B1(n_1066),
.B2(n_1005),
.Y(n_1173)
);

OR2x6_ASAP7_75t_L g1174 ( 
.A(n_1043),
.B(n_1048),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1045),
.A2(n_1044),
.B(n_966),
.C(n_1031),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1002),
.B(n_1030),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_989),
.A2(n_975),
.A3(n_1026),
.B(n_987),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1042),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_SL g1179 ( 
.A1(n_1085),
.A2(n_1007),
.B1(n_1024),
.B2(n_1020),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1046),
.A2(n_1038),
.B(n_1075),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1029),
.B(n_982),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1081),
.A2(n_1083),
.B(n_1006),
.Y(n_1182)
);

NOR4xp25_ASAP7_75t_L g1183 ( 
.A(n_1059),
.B(n_1087),
.C(n_1071),
.D(n_1067),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1003),
.B(n_1032),
.Y(n_1184)
);

NOR2xp67_ASAP7_75t_L g1185 ( 
.A(n_979),
.B(n_997),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1053),
.A2(n_1086),
.B(n_1098),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1042),
.Y(n_1187)
);

INVxp67_ASAP7_75t_SL g1188 ( 
.A(n_1068),
.Y(n_1188)
);

AOI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1036),
.A2(n_1028),
.B(n_1039),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1098),
.A2(n_1010),
.B(n_1008),
.Y(n_1190)
);

AOI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1040),
.A2(n_1073),
.B(n_1068),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_985),
.A2(n_1077),
.A3(n_1100),
.B(n_1065),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1072),
.B(n_1063),
.Y(n_1193)
);

AO32x2_ASAP7_75t_L g1194 ( 
.A1(n_1035),
.A2(n_990),
.A3(n_1091),
.B1(n_1073),
.B2(n_995),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1042),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1009),
.A2(n_977),
.B(n_1008),
.Y(n_1196)
);

OR2x2_ASAP7_75t_L g1197 ( 
.A(n_1102),
.B(n_1051),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1010),
.A2(n_1072),
.B(n_1060),
.Y(n_1198)
);

NAND2xp33_ASAP7_75t_L g1199 ( 
.A(n_995),
.B(n_1042),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1080),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_984),
.A2(n_1047),
.B(n_1049),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1047),
.A2(n_1049),
.B(n_984),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1069),
.Y(n_1203)
);

OAI21xp33_ASAP7_75t_L g1204 ( 
.A1(n_990),
.A2(n_1052),
.B(n_1070),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1088),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1014),
.A2(n_976),
.B(n_944),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_957),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_975),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_963),
.B(n_1013),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_975),
.Y(n_1210)
);

OR2x6_ASAP7_75t_L g1211 ( 
.A(n_1050),
.B(n_908),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_969),
.Y(n_1212)
);

AO32x2_ASAP7_75t_L g1213 ( 
.A1(n_1021),
.A2(n_1058),
.A3(n_964),
.B1(n_1096),
.B2(n_970),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_978),
.A2(n_963),
.B(n_889),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_957),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_963),
.B(n_1013),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_958),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_957),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1054),
.A2(n_1004),
.B(n_963),
.C(n_667),
.Y(n_1219)
);

AOI221x1_ASAP7_75t_L g1220 ( 
.A1(n_1004),
.A2(n_1058),
.B1(n_1041),
.B2(n_1027),
.C(n_1099),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1014),
.A2(n_976),
.B(n_944),
.Y(n_1221)
);

AOI21xp33_ASAP7_75t_L g1222 ( 
.A1(n_1035),
.A2(n_789),
.B(n_948),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1014),
.A2(n_976),
.B(n_944),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1054),
.A2(n_1004),
.B(n_963),
.C(n_667),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1015),
.B(n_485),
.Y(n_1225)
);

INVx1_ASAP7_75t_SL g1226 ( 
.A(n_967),
.Y(n_1226)
);

AOI211x1_ASAP7_75t_L g1227 ( 
.A1(n_1033),
.A2(n_789),
.B(n_794),
.C(n_1015),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_975),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_SL g1229 ( 
.A1(n_1041),
.A2(n_914),
.B1(n_1101),
.B2(n_990),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1014),
.A2(n_976),
.B(n_944),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_978),
.A2(n_983),
.A3(n_971),
.B(n_964),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1014),
.A2(n_976),
.B(n_944),
.Y(n_1232)
);

OA21x2_ASAP7_75t_L g1233 ( 
.A1(n_1074),
.A2(n_944),
.B(n_976),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1054),
.A2(n_1004),
.B(n_963),
.C(n_667),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_957),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_978),
.A2(n_963),
.B(n_889),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_963),
.B(n_1013),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_SL g1238 ( 
.A1(n_963),
.A2(n_889),
.B(n_959),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_963),
.B(n_1013),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_957),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1014),
.A2(n_976),
.B(n_944),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1054),
.A2(n_1004),
.B(n_963),
.C(n_667),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_963),
.B(n_1013),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1054),
.A2(n_1004),
.B(n_963),
.C(n_667),
.Y(n_1244)
);

AOI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1014),
.A2(n_978),
.B(n_961),
.Y(n_1245)
);

O2A1O1Ixp5_ASAP7_75t_L g1246 ( 
.A1(n_1027),
.A2(n_1015),
.B(n_1074),
.C(n_1025),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_975),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1103),
.Y(n_1248)
);

AO21x2_ASAP7_75t_L g1249 ( 
.A1(n_1167),
.A2(n_1157),
.B(n_1170),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_SL g1250 ( 
.A(n_1130),
.B(n_1225),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1138),
.B(n_1226),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1109),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1168),
.B(n_1120),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1119),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1220),
.A2(n_1105),
.A3(n_1158),
.B(n_1236),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1176),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_1123),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_SL g1258 ( 
.A1(n_1179),
.A2(n_1173),
.B1(n_1211),
.B2(n_1227),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1245),
.A2(n_1166),
.B(n_1206),
.Y(n_1259)
);

OAI22x1_ASAP7_75t_L g1260 ( 
.A1(n_1203),
.A2(n_1229),
.B1(n_1141),
.B2(n_1200),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1221),
.A2(n_1241),
.B(n_1223),
.Y(n_1261)
);

AOI221x1_ASAP7_75t_L g1262 ( 
.A1(n_1222),
.A2(n_1242),
.B1(n_1234),
.B2(n_1244),
.C(n_1224),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1132),
.A2(n_1164),
.B1(n_1179),
.B2(n_1104),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1154),
.B(n_1219),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1132),
.A2(n_1171),
.B(n_1186),
.C(n_1182),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1164),
.A2(n_1104),
.B1(n_1110),
.B2(n_1141),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1160),
.B(n_1181),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1211),
.B(n_1121),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1238),
.A2(n_1214),
.B(n_1114),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1184),
.B(n_1209),
.Y(n_1270)
);

AO21x2_ASAP7_75t_L g1271 ( 
.A1(n_1152),
.A2(n_1186),
.B(n_1133),
.Y(n_1271)
);

OAI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1211),
.A2(n_1136),
.B1(n_1149),
.B2(n_1165),
.Y(n_1272)
);

INVxp67_ASAP7_75t_L g1273 ( 
.A(n_1216),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1230),
.A2(n_1232),
.B(n_1137),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1177),
.Y(n_1275)
);

OAI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1135),
.A2(n_1151),
.B1(n_1243),
.B2(n_1239),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1142),
.Y(n_1277)
);

INVx4_ASAP7_75t_L g1278 ( 
.A(n_1140),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1163),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1217),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1237),
.A2(n_1204),
.B1(n_1135),
.B2(n_1134),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1131),
.A2(n_1108),
.B(n_1113),
.Y(n_1282)
);

OAI222xp33_ASAP7_75t_L g1283 ( 
.A1(n_1229),
.A2(n_1194),
.B1(n_1111),
.B2(n_1145),
.C1(n_1197),
.C2(n_1118),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1169),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1188),
.B(n_1207),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_1122),
.A2(n_1125),
.B(n_1246),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1177),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1204),
.A2(n_1143),
.B1(n_1194),
.B2(n_1117),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_1148),
.Y(n_1289)
);

NAND2x1_ASAP7_75t_L g1290 ( 
.A(n_1116),
.B(n_1178),
.Y(n_1290)
);

AOI21xp33_ASAP7_75t_SL g1291 ( 
.A1(n_1112),
.A2(n_1174),
.B(n_1193),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1177),
.Y(n_1292)
);

OA21x2_ASAP7_75t_L g1293 ( 
.A1(n_1114),
.A2(n_1147),
.B(n_1126),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1194),
.A2(n_1106),
.B1(n_1162),
.B2(n_1159),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1107),
.A2(n_1124),
.A3(n_1127),
.B(n_1156),
.Y(n_1295)
);

OA21x2_ASAP7_75t_L g1296 ( 
.A1(n_1117),
.A2(n_1106),
.B(n_1128),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1172),
.A2(n_1150),
.B(n_1161),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1162),
.A2(n_1191),
.B(n_1155),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1128),
.A2(n_1175),
.B(n_1190),
.C(n_1196),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1140),
.B(n_1146),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1180),
.A2(n_1202),
.B(n_1159),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1189),
.A2(n_1198),
.B(n_1201),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_SL g1303 ( 
.A1(n_1139),
.A2(n_1153),
.B(n_1144),
.C(n_1116),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1233),
.A2(n_1153),
.B(n_1144),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1215),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1140),
.B(n_1146),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1212),
.B(n_1218),
.Y(n_1307)
);

AOI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1235),
.A2(n_1240),
.B(n_1185),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1205),
.A2(n_1247),
.B1(n_1228),
.B2(n_1210),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1208),
.A2(n_1112),
.B(n_1231),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1174),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1212),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1212),
.B(n_1192),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1199),
.B(n_1187),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1231),
.A2(n_1115),
.B(n_1109),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1213),
.A2(n_1183),
.B1(n_1187),
.B2(n_1195),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1231),
.A2(n_1115),
.B(n_1213),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1213),
.A2(n_1183),
.B1(n_1187),
.B2(n_1195),
.Y(n_1318)
);

CKINVDCx9p33_ASAP7_75t_R g1319 ( 
.A(n_1195),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1115),
.A2(n_1220),
.A3(n_1157),
.B(n_1170),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1192),
.Y(n_1321)
);

INVxp67_ASAP7_75t_L g1322 ( 
.A(n_1192),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_SL g1323 ( 
.A1(n_1190),
.A2(n_1186),
.B(n_1182),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1209),
.B(n_1216),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1245),
.A2(n_1166),
.B(n_1206),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1132),
.A2(n_529),
.B1(n_728),
.B2(n_1004),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1245),
.A2(n_1166),
.B(n_1206),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1245),
.A2(n_1166),
.B(n_1206),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1219),
.A2(n_1244),
.B(n_1242),
.C(n_1224),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1177),
.Y(n_1330)
);

AO21x2_ASAP7_75t_L g1331 ( 
.A1(n_1167),
.A2(n_1157),
.B(n_1170),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1119),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1168),
.B(n_791),
.Y(n_1333)
);

CKINVDCx12_ASAP7_75t_R g1334 ( 
.A(n_1211),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1132),
.A2(n_529),
.B1(n_728),
.B2(n_1004),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1119),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1245),
.A2(n_1166),
.B(n_1206),
.Y(n_1337)
);

O2A1O1Ixp33_ASAP7_75t_SL g1338 ( 
.A1(n_1219),
.A2(n_1224),
.B(n_1242),
.C(n_1234),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1119),
.Y(n_1339)
);

OA21x2_ASAP7_75t_L g1340 ( 
.A1(n_1157),
.A2(n_1221),
.B(n_1206),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_1211),
.B(n_1164),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1103),
.Y(n_1342)
);

NAND2xp33_ASAP7_75t_L g1343 ( 
.A(n_1171),
.B(n_782),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1103),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1245),
.A2(n_1166),
.B(n_1206),
.Y(n_1345)
);

OAI221xp5_ASAP7_75t_SL g1346 ( 
.A1(n_1154),
.A2(n_1041),
.B1(n_504),
.B2(n_1004),
.C(n_516),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1219),
.A2(n_1234),
.B(n_1242),
.C(n_1224),
.Y(n_1347)
);

OA21x2_ASAP7_75t_L g1348 ( 
.A1(n_1157),
.A2(n_1221),
.B(n_1206),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1177),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1219),
.A2(n_1234),
.B(n_1224),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1219),
.A2(n_1234),
.B(n_1224),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1132),
.A2(n_529),
.B1(n_728),
.B2(n_1004),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1177),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1132),
.A2(n_529),
.B1(n_728),
.B2(n_1004),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1245),
.A2(n_1166),
.B(n_1206),
.Y(n_1355)
);

BUFx8_ASAP7_75t_L g1356 ( 
.A(n_1123),
.Y(n_1356)
);

BUFx2_ASAP7_75t_SL g1357 ( 
.A(n_1103),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_R g1358 ( 
.A(n_1136),
.B(n_655),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1119),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1176),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1245),
.A2(n_1166),
.B(n_1206),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1119),
.Y(n_1362)
);

AOI221x1_ASAP7_75t_L g1363 ( 
.A1(n_1222),
.A2(n_1004),
.B1(n_1219),
.B2(n_1234),
.C(n_1224),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1154),
.B(n_1015),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1154),
.A2(n_1004),
.B1(n_559),
.B2(n_695),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1140),
.B(n_1146),
.Y(n_1366)
);

NAND2x1p5_ASAP7_75t_L g1367 ( 
.A(n_1193),
.B(n_1129),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1168),
.B(n_791),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1132),
.A2(n_529),
.B1(n_728),
.B2(n_1004),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1132),
.A2(n_529),
.B1(n_728),
.B2(n_1004),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1229),
.A2(n_1104),
.B1(n_1179),
.B2(n_1101),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1219),
.A2(n_1234),
.B(n_1224),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1358),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1341),
.B(n_1300),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1253),
.B(n_1268),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1252),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1329),
.A2(n_1264),
.B(n_1347),
.Y(n_1377)
);

O2A1O1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1346),
.A2(n_1329),
.B(n_1264),
.C(n_1338),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1270),
.B(n_1256),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1343),
.A2(n_1265),
.B(n_1338),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1327),
.A2(n_1337),
.B(n_1328),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1333),
.B(n_1368),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1365),
.A2(n_1364),
.B1(n_1350),
.B2(n_1351),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1267),
.B(n_1307),
.Y(n_1384)
);

INVx2_ASAP7_75t_SL g1385 ( 
.A(n_1285),
.Y(n_1385)
);

O2A1O1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1372),
.A2(n_1265),
.B(n_1343),
.C(n_1364),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1267),
.B(n_1254),
.Y(n_1387)
);

AOI21x1_ASAP7_75t_SL g1388 ( 
.A1(n_1356),
.A2(n_1358),
.B(n_1324),
.Y(n_1388)
);

O2A1O1Ixp5_ASAP7_75t_L g1389 ( 
.A1(n_1299),
.A2(n_1272),
.B(n_1276),
.C(n_1314),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1315),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_SL g1391 ( 
.A1(n_1363),
.A2(n_1262),
.B(n_1278),
.Y(n_1391)
);

AOI21x1_ASAP7_75t_SL g1392 ( 
.A1(n_1356),
.A2(n_1250),
.B(n_1357),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1277),
.B(n_1279),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_R g1394 ( 
.A(n_1334),
.B(n_1311),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1339),
.B(n_1311),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1284),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1263),
.A2(n_1354),
.B1(n_1335),
.B2(n_1370),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1293),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1305),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1280),
.B(n_1336),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1304),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1263),
.A2(n_1354),
.B1(n_1352),
.B2(n_1335),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_SL g1403 ( 
.A1(n_1278),
.A2(n_1272),
.B(n_1299),
.Y(n_1403)
);

AO21x2_ASAP7_75t_L g1404 ( 
.A1(n_1249),
.A2(n_1331),
.B(n_1276),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1326),
.A2(n_1352),
.B1(n_1370),
.B2(n_1369),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1326),
.A2(n_1369),
.B1(n_1294),
.B2(n_1371),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1321),
.Y(n_1407)
);

OR2x6_ASAP7_75t_L g1408 ( 
.A(n_1341),
.B(n_1260),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1323),
.A2(n_1291),
.B(n_1283),
.C(n_1296),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1248),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1293),
.Y(n_1411)
);

AOI211xp5_ASAP7_75t_L g1412 ( 
.A1(n_1258),
.A2(n_1314),
.B(n_1257),
.C(n_1303),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1280),
.B(n_1336),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1266),
.A2(n_1289),
.B1(n_1288),
.B2(n_1318),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1271),
.A2(n_1366),
.B(n_1306),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1266),
.A2(n_1289),
.B1(n_1288),
.B2(n_1318),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1345),
.A2(n_1355),
.B(n_1361),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1359),
.B(n_1362),
.Y(n_1418)
);

O2A1O1Ixp5_ASAP7_75t_L g1419 ( 
.A1(n_1290),
.A2(n_1308),
.B(n_1360),
.C(n_1292),
.Y(n_1419)
);

A2O1A1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1316),
.A2(n_1281),
.B(n_1317),
.C(n_1310),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1316),
.A2(n_1302),
.B(n_1297),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1359),
.B(n_1362),
.Y(n_1422)
);

O2A1O1Ixp5_ASAP7_75t_L g1423 ( 
.A1(n_1275),
.A2(n_1292),
.B(n_1287),
.C(n_1353),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1261),
.A2(n_1274),
.B(n_1282),
.Y(n_1424)
);

NOR2xp67_ASAP7_75t_L g1425 ( 
.A(n_1273),
.B(n_1332),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1281),
.A2(n_1367),
.B1(n_1344),
.B2(n_1342),
.Y(n_1426)
);

O2A1O1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1340),
.A2(n_1348),
.B(n_1286),
.C(n_1298),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1313),
.B(n_1320),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1340),
.Y(n_1429)
);

AOI221xp5_ASAP7_75t_L g1430 ( 
.A1(n_1322),
.A2(n_1309),
.B1(n_1353),
.B2(n_1287),
.C(n_1349),
.Y(n_1430)
);

O2A1O1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1348),
.A2(n_1286),
.B(n_1320),
.C(n_1330),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1312),
.B(n_1320),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1295),
.B(n_1255),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1295),
.B(n_1255),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1295),
.B(n_1309),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1301),
.B(n_1251),
.Y(n_1436)
);

CKINVDCx6p67_ASAP7_75t_R g1437 ( 
.A(n_1357),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1253),
.B(n_1268),
.Y(n_1438)
);

CKINVDCx9p33_ASAP7_75t_R g1439 ( 
.A(n_1319),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1343),
.A2(n_1269),
.B(n_1171),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1269),
.A2(n_1325),
.B(n_1259),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1253),
.B(n_1268),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1252),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1251),
.B(n_1270),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1251),
.B(n_1270),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1343),
.A2(n_1269),
.B(n_1171),
.Y(n_1446)
);

INVx2_ASAP7_75t_SL g1447 ( 
.A(n_1285),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1264),
.A2(n_1365),
.B1(n_1346),
.B2(n_1329),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1264),
.A2(n_1365),
.B1(n_1346),
.B2(n_1329),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1329),
.A2(n_1224),
.B(n_1219),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1264),
.A2(n_1365),
.B1(n_1346),
.B2(n_1329),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1264),
.A2(n_1365),
.B1(n_1346),
.B2(n_1329),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1253),
.B(n_1268),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1264),
.A2(n_1365),
.B1(n_1346),
.B2(n_1329),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1285),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1253),
.B(n_1268),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1252),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1377),
.B(n_1383),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_1387),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1396),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1376),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1448),
.B(n_1449),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1433),
.B(n_1434),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1398),
.B(n_1411),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1398),
.B(n_1411),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1437),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1401),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1440),
.A2(n_1446),
.B(n_1421),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1407),
.Y(n_1469)
);

OA21x2_ASAP7_75t_L g1470 ( 
.A1(n_1420),
.A2(n_1380),
.B(n_1429),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1429),
.B(n_1435),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1404),
.B(n_1436),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1424),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1404),
.B(n_1432),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1428),
.B(n_1399),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1420),
.A2(n_1419),
.B(n_1390),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1423),
.A2(n_1389),
.B(n_1430),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1374),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1451),
.B(n_1452),
.Y(n_1479)
);

BUFx12f_ASAP7_75t_L g1480 ( 
.A(n_1373),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1443),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1385),
.B(n_1447),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1431),
.B(n_1441),
.Y(n_1483)
);

NAND4xp25_ASAP7_75t_L g1484 ( 
.A(n_1386),
.B(n_1378),
.C(n_1450),
.D(n_1454),
.Y(n_1484)
);

NAND4xp25_ASAP7_75t_L g1485 ( 
.A(n_1391),
.B(n_1427),
.C(n_1426),
.D(n_1403),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1441),
.B(n_1385),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1409),
.B(n_1412),
.Y(n_1487)
);

AO21x2_ASAP7_75t_L g1488 ( 
.A1(n_1414),
.A2(n_1416),
.B(n_1457),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1393),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1381),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1447),
.B(n_1455),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1417),
.Y(n_1492)
);

INVxp67_ASAP7_75t_L g1493 ( 
.A(n_1384),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1400),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1439),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1471),
.B(n_1486),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1472),
.B(n_1379),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1461),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1471),
.B(n_1382),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1460),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1460),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1461),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1471),
.B(n_1375),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1486),
.B(n_1456),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1473),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1464),
.B(n_1465),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1462),
.A2(n_1406),
.B1(n_1397),
.B2(n_1402),
.Y(n_1507)
);

AOI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1462),
.A2(n_1405),
.B1(n_1415),
.B2(n_1444),
.C(n_1445),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1470),
.B(n_1453),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1464),
.B(n_1442),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1470),
.B(n_1438),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1490),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1470),
.B(n_1422),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1470),
.B(n_1418),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1469),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1470),
.B(n_1463),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1470),
.B(n_1413),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1495),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1499),
.B(n_1459),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1510),
.B(n_1459),
.Y(n_1520)
);

OAI21xp33_ASAP7_75t_SL g1521 ( 
.A1(n_1516),
.A2(n_1485),
.B(n_1458),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1507),
.A2(n_1484),
.B1(n_1479),
.B2(n_1458),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1518),
.B(n_1478),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1515),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1507),
.A2(n_1479),
.B1(n_1495),
.B2(n_1487),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1500),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1510),
.B(n_1482),
.Y(n_1527)
);

OAI33xp33_ASAP7_75t_L g1528 ( 
.A1(n_1497),
.A2(n_1487),
.A3(n_1484),
.B1(n_1491),
.B2(n_1489),
.B3(n_1485),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1510),
.B(n_1482),
.Y(n_1529)
);

OAI211xp5_ASAP7_75t_L g1530 ( 
.A1(n_1508),
.A2(n_1516),
.B(n_1468),
.C(n_1514),
.Y(n_1530)
);

OR2x6_ASAP7_75t_L g1531 ( 
.A(n_1518),
.B(n_1415),
.Y(n_1531)
);

NAND4xp25_ASAP7_75t_SL g1532 ( 
.A(n_1516),
.B(n_1508),
.C(n_1511),
.D(n_1509),
.Y(n_1532)
);

AOI222xp33_ASAP7_75t_L g1533 ( 
.A1(n_1508),
.A2(n_1463),
.B1(n_1474),
.B2(n_1475),
.C1(n_1483),
.C2(n_1472),
.Y(n_1533)
);

AOI221xp5_ASAP7_75t_L g1534 ( 
.A1(n_1516),
.A2(n_1472),
.B1(n_1483),
.B2(n_1488),
.C(n_1474),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1499),
.B(n_1497),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1509),
.A2(n_1488),
.B1(n_1477),
.B2(n_1463),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1518),
.A2(n_1495),
.B1(n_1493),
.B2(n_1494),
.Y(n_1537)
);

INVx4_ASAP7_75t_L g1538 ( 
.A(n_1518),
.Y(n_1538)
);

OAI222xp33_ASAP7_75t_SL g1539 ( 
.A1(n_1502),
.A2(n_1392),
.B1(n_1437),
.B2(n_1466),
.C1(n_1480),
.C2(n_1388),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1500),
.Y(n_1540)
);

BUFx10_ASAP7_75t_L g1541 ( 
.A(n_1498),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1509),
.A2(n_1488),
.B1(n_1408),
.B2(n_1475),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1515),
.Y(n_1543)
);

OAI211xp5_ASAP7_75t_L g1544 ( 
.A1(n_1513),
.A2(n_1468),
.B(n_1481),
.C(n_1467),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1500),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_SL g1546 ( 
.A1(n_1509),
.A2(n_1488),
.B1(n_1476),
.B2(n_1477),
.Y(n_1546)
);

NAND3xp33_ASAP7_75t_L g1547 ( 
.A(n_1502),
.B(n_1474),
.C(n_1476),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1518),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1501),
.Y(n_1549)
);

INVxp67_ASAP7_75t_SL g1550 ( 
.A(n_1505),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1510),
.B(n_1493),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_1499),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_1499),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1497),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1511),
.A2(n_1477),
.B1(n_1408),
.B2(n_1476),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1504),
.Y(n_1556)
);

OA21x2_ASAP7_75t_L g1557 ( 
.A1(n_1512),
.A2(n_1492),
.B(n_1490),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1526),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1531),
.B(n_1513),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1557),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1540),
.Y(n_1561)
);

INVx3_ASAP7_75t_L g1562 ( 
.A(n_1538),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1545),
.Y(n_1563)
);

NOR2x1p5_ASAP7_75t_L g1564 ( 
.A(n_1538),
.B(n_1480),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1556),
.B(n_1496),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1549),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1557),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1521),
.B(n_1511),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1524),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1551),
.B(n_1511),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1534),
.B(n_1513),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1541),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1543),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1557),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1531),
.B(n_1513),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1527),
.Y(n_1576)
);

INVxp67_ASAP7_75t_SL g1577 ( 
.A(n_1547),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1551),
.B(n_1503),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1529),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1520),
.Y(n_1580)
);

INVx4_ASAP7_75t_L g1581 ( 
.A(n_1548),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1535),
.B(n_1503),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1533),
.B(n_1514),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1541),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1550),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1532),
.B(n_1506),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1550),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1554),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1552),
.B(n_1514),
.Y(n_1589)
);

INVx5_ASAP7_75t_L g1590 ( 
.A(n_1523),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1523),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1563),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1576),
.B(n_1579),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1558),
.Y(n_1594)
);

NAND2x1p5_ASAP7_75t_L g1595 ( 
.A(n_1564),
.B(n_1477),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1568),
.B(n_1590),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1590),
.B(n_1514),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1572),
.B(n_1528),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1577),
.A2(n_1522),
.B(n_1525),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1591),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1590),
.B(n_1517),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1590),
.B(n_1553),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1558),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1590),
.B(n_1564),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1576),
.B(n_1506),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1571),
.A2(n_1528),
.B(n_1530),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1561),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1588),
.B(n_1522),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1588),
.B(n_1536),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1578),
.B(n_1536),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1567),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1561),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1566),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1591),
.B(n_1565),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1566),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1580),
.B(n_1583),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1569),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1580),
.B(n_1546),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1584),
.Y(n_1619)
);

INVxp67_ASAP7_75t_L g1620 ( 
.A(n_1572),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1586),
.B(n_1506),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1591),
.B(n_1496),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1569),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1573),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1567),
.Y(n_1625)
);

OAI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1586),
.A2(n_1546),
.B1(n_1542),
.B2(n_1555),
.C(n_1544),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1567),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1594),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1594),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1599),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_L g1631 ( 
.A(n_1606),
.B(n_1555),
.C(n_1584),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1607),
.Y(n_1632)
);

INVx2_ASAP7_75t_SL g1633 ( 
.A(n_1600),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1616),
.B(n_1593),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1596),
.B(n_1562),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1598),
.B(n_1570),
.Y(n_1636)
);

NAND4xp25_ASAP7_75t_L g1637 ( 
.A(n_1596),
.B(n_1581),
.C(n_1537),
.D(n_1589),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1608),
.A2(n_1559),
.B(n_1575),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1600),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1593),
.B(n_1582),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1607),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1619),
.B(n_1581),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1612),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1614),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1621),
.B(n_1519),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1612),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1613),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1592),
.B(n_1581),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1592),
.B(n_1581),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1614),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_SL g1652 ( 
.A1(n_1626),
.A2(n_1373),
.B(n_1575),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1613),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1615),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1615),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1604),
.B(n_1559),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1621),
.B(n_1573),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1603),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1604),
.B(n_1559),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1617),
.Y(n_1660)
);

OAI21xp33_ASAP7_75t_SL g1661 ( 
.A1(n_1610),
.A2(n_1585),
.B(n_1567),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1605),
.B(n_1585),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1634),
.B(n_1630),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1633),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1633),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1639),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1651),
.B(n_1604),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1651),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1644),
.B(n_1620),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1630),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1636),
.B(n_1609),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1653),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1653),
.Y(n_1673)
);

INVx1_ASAP7_75t_SL g1674 ( 
.A(n_1642),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1661),
.B(n_1410),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1640),
.B(n_1605),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1658),
.B(n_1617),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1628),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1648),
.Y(n_1679)
);

AND3x1_ASAP7_75t_L g1680 ( 
.A(n_1635),
.B(n_1602),
.C(n_1618),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1656),
.B(n_1622),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1656),
.B(n_1622),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1660),
.B(n_1623),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1635),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1649),
.B(n_1410),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1638),
.A2(n_1625),
.B(n_1627),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1629),
.Y(n_1687)
);

NOR2x1_ASAP7_75t_L g1688 ( 
.A(n_1670),
.B(n_1652),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1672),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1684),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1680),
.A2(n_1631),
.B1(n_1652),
.B2(n_1595),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1681),
.B(n_1659),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1671),
.A2(n_1595),
.B1(n_1560),
.B2(n_1574),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1680),
.A2(n_1597),
.B1(n_1601),
.B2(n_1595),
.Y(n_1694)
);

AOI222xp33_ASAP7_75t_L g1695 ( 
.A1(n_1670),
.A2(n_1574),
.B1(n_1560),
.B2(n_1650),
.C1(n_1641),
.C2(n_1655),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1672),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1672),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1663),
.A2(n_1601),
.B1(n_1597),
.B2(n_1662),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1663),
.A2(n_1675),
.B1(n_1637),
.B2(n_1666),
.C(n_1676),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1673),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1673),
.Y(n_1701)
);

OAI32xp33_ASAP7_75t_L g1702 ( 
.A1(n_1666),
.A2(n_1662),
.A3(n_1657),
.B1(n_1632),
.B2(n_1643),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1684),
.B(n_1646),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1676),
.B(n_1645),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1678),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1678),
.Y(n_1706)
);

NAND3xp33_ASAP7_75t_L g1707 ( 
.A(n_1695),
.B(n_1665),
.C(n_1664),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1690),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1704),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1689),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1692),
.B(n_1669),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1696),
.B(n_1668),
.Y(n_1712)
);

NAND2x1p5_ASAP7_75t_L g1713 ( 
.A(n_1688),
.B(n_1669),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1703),
.B(n_1679),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1697),
.B(n_1681),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1702),
.B(n_1679),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1691),
.B(n_1667),
.Y(n_1717)
);

OAI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1691),
.A2(n_1677),
.B1(n_1674),
.B2(n_1683),
.C(n_1650),
.Y(n_1718)
);

XNOR2x1_ASAP7_75t_L g1719 ( 
.A(n_1713),
.B(n_1674),
.Y(n_1719)
);

OAI211xp5_ASAP7_75t_L g1720 ( 
.A1(n_1716),
.A2(n_1699),
.B(n_1706),
.C(n_1705),
.Y(n_1720)
);

AOI211xp5_ASAP7_75t_L g1721 ( 
.A1(n_1718),
.A2(n_1694),
.B(n_1698),
.C(n_1686),
.Y(n_1721)
);

NAND4xp25_ASAP7_75t_L g1722 ( 
.A(n_1707),
.B(n_1667),
.C(n_1700),
.D(n_1701),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1711),
.B(n_1682),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1709),
.A2(n_1693),
.B1(n_1698),
.B2(n_1686),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1714),
.B(n_1682),
.Y(n_1725)
);

AOI211xp5_ASAP7_75t_SL g1726 ( 
.A1(n_1708),
.A2(n_1712),
.B(n_1710),
.C(n_1715),
.Y(n_1726)
);

OAI211xp5_ASAP7_75t_L g1727 ( 
.A1(n_1717),
.A2(n_1687),
.B(n_1677),
.C(n_1683),
.Y(n_1727)
);

OAI21xp5_ASAP7_75t_SL g1728 ( 
.A1(n_1713),
.A2(n_1659),
.B(n_1687),
.Y(n_1728)
);

O2A1O1Ixp5_ASAP7_75t_SL g1729 ( 
.A1(n_1712),
.A2(n_1654),
.B(n_1647),
.C(n_1623),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1719),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1723),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1725),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1726),
.Y(n_1733)
);

AOI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1720),
.A2(n_1685),
.B(n_1611),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1732),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1733),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1733),
.B(n_1722),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1730),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1731),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1730),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1738),
.Y(n_1741)
);

CKINVDCx16_ASAP7_75t_R g1742 ( 
.A(n_1738),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1740),
.Y(n_1743)
);

OA22x2_ASAP7_75t_L g1744 ( 
.A1(n_1736),
.A2(n_1728),
.B1(n_1724),
.B2(n_1727),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1735),
.Y(n_1745)
);

INVxp67_ASAP7_75t_SL g1746 ( 
.A(n_1741),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1742),
.B(n_1739),
.Y(n_1747)
);

NOR4xp75_ASAP7_75t_L g1748 ( 
.A(n_1744),
.B(n_1737),
.C(n_1721),
.D(n_1734),
.Y(n_1748)
);

AND3x1_ASAP7_75t_L g1749 ( 
.A(n_1747),
.B(n_1741),
.C(n_1743),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1749),
.B(n_1746),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1750),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1750),
.Y(n_1752)
);

XNOR2xp5_ASAP7_75t_L g1753 ( 
.A(n_1751),
.B(n_1748),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1752),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1753),
.Y(n_1755)
);

XNOR2xp5_ASAP7_75t_L g1756 ( 
.A(n_1754),
.B(n_1745),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1756),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1757),
.A2(n_1755),
.B(n_1625),
.Y(n_1758)
);

OAI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1758),
.A2(n_1729),
.B(n_1627),
.Y(n_1759)
);

OAI221xp5_ASAP7_75t_R g1760 ( 
.A1(n_1759),
.A2(n_1539),
.B1(n_1597),
.B2(n_1601),
.C(n_1602),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1760),
.A2(n_1480),
.B1(n_1587),
.B2(n_1624),
.Y(n_1761)
);

AOI211xp5_ASAP7_75t_L g1762 ( 
.A1(n_1761),
.A2(n_1394),
.B(n_1425),
.C(n_1395),
.Y(n_1762)
);


endmodule