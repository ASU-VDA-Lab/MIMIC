module fake_jpeg_31056_n_490 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_490);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_490;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_55),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_17),
.B(n_9),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_56),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_17),
.B(n_9),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_63),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_69),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_25),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_72),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_22),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_30),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_73),
.B(n_79),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_78),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_83),
.B(n_93),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_30),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_85),
.B(n_86),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_38),
.B(n_9),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_32),
.B(n_9),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_87),
.B(n_90),
.Y(n_163)
);

BUFx4f_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_32),
.B(n_8),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_24),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_18),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_97),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_30),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_98),
.B(n_100),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_39),
.B(n_8),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_101),
.B(n_16),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_22),
.B(n_8),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_103),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_20),
.B1(n_36),
.B2(n_37),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_107),
.A2(n_118),
.B1(n_122),
.B2(n_129),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_54),
.A2(n_36),
.B1(n_39),
.B2(n_20),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_109),
.A2(n_130),
.B1(n_149),
.B2(n_99),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_58),
.A2(n_20),
.B1(n_40),
.B2(n_19),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_27),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_121),
.B(n_134),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_61),
.A2(n_40),
.B1(n_48),
.B2(n_19),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_75),
.A2(n_27),
.B1(n_48),
.B2(n_43),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_125),
.A2(n_139),
.B1(n_89),
.B2(n_66),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_64),
.A2(n_48),
.B1(n_43),
.B2(n_29),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_68),
.A2(n_29),
.B1(n_28),
.B2(n_24),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_70),
.A2(n_48),
.B1(n_43),
.B2(n_28),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_131),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_51),
.B(n_33),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_65),
.B(n_33),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_136),
.B(n_157),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_74),
.A2(n_42),
.B1(n_33),
.B2(n_43),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_78),
.A2(n_33),
.B1(n_2),
.B2(n_3),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_80),
.A2(n_11),
.B1(n_3),
.B2(n_5),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_152),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_50),
.B(n_11),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_81),
.A2(n_8),
.B1(n_3),
.B2(n_5),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_158),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_59),
.B(n_12),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_12),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_67),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_164),
.B(n_181),
.Y(n_251)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_165),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_116),
.A2(n_94),
.B1(n_92),
.B2(n_91),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_166),
.A2(n_169),
.B1(n_211),
.B2(n_217),
.Y(n_225)
);

BUFx4f_ASAP7_75t_SL g167 ( 
.A(n_120),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_167),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_168),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_L g169 ( 
.A1(n_128),
.A2(n_96),
.B1(n_82),
.B2(n_100),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_172),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_116),
.B(n_85),
.C(n_98),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_173),
.B(n_179),
.C(n_209),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_108),
.Y(n_174)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_174),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_175),
.Y(n_223)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_177),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_73),
.C(n_88),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_180),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_67),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_121),
.B(n_88),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_182),
.B(n_188),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_104),
.B(n_63),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_192),
.Y(n_222)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_106),
.Y(n_184)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_184),
.Y(n_258)
);

O2A1O1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_136),
.A2(n_63),
.B(n_56),
.C(n_84),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_186),
.A2(n_154),
.B(n_142),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_L g187 ( 
.A1(n_114),
.A2(n_56),
.B(n_84),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_187),
.B(n_208),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_145),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_76),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_194),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_69),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_151),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_195),
.B(n_199),
.Y(n_248)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_127),
.Y(n_196)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_196),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_117),
.B(n_69),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_198),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_119),
.B(n_57),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_160),
.B(n_95),
.Y(n_199)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_200),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_153),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_201),
.B(n_202),
.Y(n_257)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_142),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_203),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_204),
.A2(n_143),
.B1(n_112),
.B2(n_123),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_144),
.B(n_62),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_207),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_132),
.B(n_133),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_115),
.B(n_57),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_52),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_132),
.B(n_133),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_215),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_138),
.A2(n_97),
.B1(n_77),
.B2(n_62),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_212),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_214),
.A2(n_147),
.B1(n_135),
.B2(n_124),
.Y(n_260)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_159),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_108),
.A2(n_99),
.B1(n_5),
.B2(n_6),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_174),
.A2(n_108),
.B(n_112),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_218),
.A2(n_209),
.B(n_189),
.Y(n_264)
);

AND2x2_ASAP7_75t_SL g220 ( 
.A(n_191),
.B(n_137),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_220),
.B(n_167),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_137),
.C(n_123),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_179),
.C(n_170),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_166),
.A2(n_125),
.B1(n_146),
.B2(n_148),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_229),
.A2(n_252),
.B1(n_256),
.B2(n_260),
.Y(n_265)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_128),
.B1(n_148),
.B2(n_159),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_231),
.A2(n_239),
.B1(n_249),
.B2(n_209),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_174),
.A2(n_111),
.B(n_156),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_243),
.A2(n_218),
.B(n_242),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_170),
.B(n_111),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_194),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_247),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_173),
.A2(n_113),
.B1(n_141),
.B2(n_140),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_213),
.A2(n_113),
.B1(n_141),
.B2(n_140),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_195),
.A2(n_185),
.B1(n_189),
.B2(n_217),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_261),
.B(n_266),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_264),
.A2(n_288),
.B(n_241),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_206),
.C(n_210),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_188),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_273),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_296),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_269),
.A2(n_282),
.B(n_294),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_221),
.C(n_236),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_277),
.Y(n_310)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_219),
.Y(n_271)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_272),
.A2(n_275),
.B1(n_291),
.B2(n_295),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_222),
.B(n_176),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_219),
.Y(n_274)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_248),
.A2(n_169),
.B1(n_204),
.B2(n_193),
.Y(n_275)
);

INVx4_ASAP7_75t_SL g276 ( 
.A(n_259),
.Y(n_276)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_276),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_207),
.C(n_184),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_254),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_278),
.B(n_280),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_237),
.B(n_171),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_279),
.B(n_245),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_239),
.A2(n_165),
.B1(n_186),
.B2(n_202),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_281),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_243),
.A2(n_215),
.B(n_212),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_290),
.Y(n_317)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_232),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_284),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_228),
.A2(n_167),
.B(n_168),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_285),
.A2(n_227),
.B(n_230),
.Y(n_306)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_232),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_286),
.Y(n_314)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_244),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_287),
.Y(n_321)
);

OAI22x1_ASAP7_75t_L g288 ( 
.A1(n_247),
.A2(n_175),
.B1(n_190),
.B2(n_142),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_244),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_289),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_220),
.B(n_216),
.C(n_196),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_249),
.A2(n_147),
.B1(n_135),
.B2(n_172),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_220),
.B(n_177),
.C(n_201),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_226),
.C(n_227),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_235),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_224),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_242),
.A2(n_203),
.B1(n_126),
.B2(n_180),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_225),
.A2(n_178),
.B1(n_126),
.B2(n_7),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_224),
.B(n_200),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_296),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_297),
.B(n_298),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_282),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_SL g300 ( 
.A(n_288),
.B(n_228),
.C(n_256),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_300),
.A2(n_311),
.B(n_313),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_294),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_301),
.B(n_316),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_302),
.B(n_268),
.Y(n_331)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_276),
.Y(n_303)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_303),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_261),
.C(n_270),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_291),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_307),
.A2(n_324),
.B(n_318),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_262),
.A2(n_264),
.B(n_285),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_262),
.A2(n_226),
.B(n_258),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_279),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_271),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_319),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_275),
.A2(n_225),
.B1(n_229),
.B2(n_252),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_323),
.A2(n_265),
.B1(n_263),
.B2(n_295),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_280),
.A2(n_258),
.B(n_241),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_328),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_329),
.A2(n_353),
.B1(n_326),
.B2(n_321),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_343),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_316),
.B(n_263),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g383 ( 
.A(n_332),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_302),
.B(n_277),
.Y(n_335)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_335),
.Y(n_359)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_305),
.Y(n_336)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_336),
.Y(n_373)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_305),
.Y(n_337)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_337),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_338),
.B(n_346),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_325),
.A2(n_272),
.B1(n_281),
.B2(n_266),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_339),
.A2(n_342),
.B1(n_358),
.B2(n_322),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_340),
.A2(n_345),
.B(n_349),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_297),
.B(n_292),
.Y(n_341)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_341),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_298),
.A2(n_300),
.B1(n_313),
.B2(n_306),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_308),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_309),
.B(n_283),
.C(n_290),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_344),
.B(n_347),
.C(n_317),
.Y(n_367)
);

AO22x1_ASAP7_75t_L g345 ( 
.A1(n_318),
.A2(n_269),
.B1(n_265),
.B2(n_231),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_309),
.B(n_293),
.C(n_289),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_315),
.B(n_287),
.Y(n_348)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_348),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_307),
.A2(n_286),
.B(n_284),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_327),
.Y(n_351)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_327),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_352),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_322),
.A2(n_274),
.B1(n_276),
.B2(n_234),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_315),
.B(n_253),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_357),
.Y(n_369)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_308),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_301),
.A2(n_234),
.B1(n_238),
.B2(n_253),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_360),
.A2(n_362),
.B1(n_363),
.B2(n_353),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_310),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_361),
.B(n_380),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_358),
.A2(n_303),
.B1(n_319),
.B2(n_320),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_346),
.A2(n_323),
.B1(n_317),
.B2(n_310),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_340),
.A2(n_311),
.B(n_324),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_350),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_366),
.B(n_375),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_370),
.C(n_379),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_304),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_368),
.B(n_335),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_347),
.B(n_304),
.C(n_321),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_371),
.A2(n_345),
.B1(n_333),
.B2(n_329),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_332),
.B(n_326),
.Y(n_374)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_374),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_350),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_341),
.B(n_314),
.C(n_312),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_342),
.B(n_299),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_314),
.Y(n_381)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_381),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_334),
.B(n_339),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_385),
.B(n_355),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_356),
.Y(n_388)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_388),
.Y(n_412)
);

FAx1_ASAP7_75t_SL g389 ( 
.A(n_372),
.B(n_354),
.CI(n_355),
.CON(n_389),
.SN(n_389)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_397),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_396),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_364),
.B(n_334),
.Y(n_393)
);

AO21x1_ASAP7_75t_L g414 ( 
.A1(n_393),
.A2(n_378),
.B(n_369),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_361),
.B(n_349),
.C(n_346),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_395),
.B(n_410),
.C(n_363),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_380),
.B(n_356),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_398),
.A2(n_384),
.B1(n_365),
.B2(n_373),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_379),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_399),
.B(n_406),
.Y(n_417)
);

MAJx2_ASAP7_75t_L g400 ( 
.A(n_370),
.B(n_345),
.C(n_331),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_409),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_375),
.B(n_333),
.Y(n_401)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_401),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_359),
.B(n_233),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_404),
.B(n_407),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_405),
.A2(n_384),
.B1(n_382),
.B2(n_359),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_352),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_369),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_374),
.B(n_336),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_408),
.B(n_381),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_368),
.B(n_351),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_367),
.B(n_337),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_403),
.Y(n_411)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_411),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_SL g413 ( 
.A(n_396),
.B(n_372),
.C(n_385),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_426),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_400),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_415),
.B(n_423),
.Y(n_437)
);

A2O1A1Ixp33_ASAP7_75t_SL g420 ( 
.A1(n_390),
.A2(n_378),
.B(n_360),
.C(n_371),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_420),
.A2(n_424),
.B(n_389),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_421),
.A2(n_428),
.B1(n_407),
.B2(n_398),
.Y(n_430)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_422),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_390),
.A2(n_365),
.B(n_382),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_387),
.A2(n_402),
.B(n_393),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_425),
.A2(n_330),
.B1(n_386),
.B2(n_409),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_410),
.B(n_377),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_393),
.A2(n_330),
.B1(n_376),
.B2(n_373),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_439),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_412),
.A2(n_386),
.B1(n_376),
.B2(n_395),
.Y(n_431)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_431),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_432),
.A2(n_434),
.B(n_420),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_424),
.A2(n_389),
.B(n_399),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_433),
.A2(n_423),
.B(n_414),
.Y(n_445)
);

XNOR2x1_ASAP7_75t_L g435 ( 
.A(n_418),
.B(n_392),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_435),
.B(n_436),
.C(n_438),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_394),
.C(n_392),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_427),
.B(n_394),
.C(n_391),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_419),
.B(n_357),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_441),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_416),
.B(n_312),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_442),
.B(n_343),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_445),
.A2(n_246),
.B(n_240),
.Y(n_468)
);

INVxp33_ASAP7_75t_L g447 ( 
.A(n_441),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_439),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_444),
.B(n_421),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_452),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_432),
.A2(n_417),
.B(n_428),
.Y(n_450)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_450),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_434),
.A2(n_411),
.B1(n_420),
.B2(n_429),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_451),
.A2(n_435),
.B1(n_259),
.B2(n_223),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_427),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_453),
.B(n_457),
.Y(n_464)
);

OAI321xp33_ASAP7_75t_L g456 ( 
.A1(n_430),
.A2(n_420),
.A3(n_418),
.B1(n_303),
.B2(n_254),
.C(n_233),
.Y(n_456)
);

NAND3xp33_ASAP7_75t_L g465 ( 
.A(n_456),
.B(n_223),
.C(n_255),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_443),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_458),
.A2(n_255),
.B(n_246),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_451),
.A2(n_433),
.B1(n_437),
.B2(n_440),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_460),
.B(n_462),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_465),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_455),
.B(n_438),
.C(n_436),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_466),
.A2(n_468),
.B1(n_448),
.B2(n_454),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_467),
.B(n_469),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_455),
.B(n_240),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_477),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_462),
.B(n_446),
.C(n_458),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_472),
.B(n_476),
.Y(n_478)
);

AND2x2_ASAP7_75t_SL g475 ( 
.A(n_459),
.B(n_447),
.Y(n_475)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_475),
.Y(n_481)
);

NOR3xp33_ASAP7_75t_SL g476 ( 
.A(n_464),
.B(n_448),
.C(n_190),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_465),
.A2(n_238),
.B1(n_6),
.B2(n_13),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_473),
.B(n_460),
.C(n_463),
.Y(n_479)
);

NAND3xp33_ASAP7_75t_L g485 ( 
.A(n_479),
.B(n_6),
.C(n_13),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_471),
.A2(n_190),
.B(n_6),
.Y(n_482)
);

AOI21x1_ASAP7_75t_L g484 ( 
.A1(n_482),
.A2(n_480),
.B(n_474),
.Y(n_484)
);

AOI321xp33_ASAP7_75t_L g483 ( 
.A1(n_478),
.A2(n_475),
.A3(n_471),
.B1(n_474),
.B2(n_14),
.C(n_15),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_483),
.A2(n_13),
.B(n_15),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_484),
.A2(n_485),
.B(n_481),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_486),
.A2(n_487),
.B(n_16),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_488),
.A2(n_0),
.B1(n_15),
.B2(n_333),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_489),
.B(n_15),
.Y(n_490)
);


endmodule