module fake_jpeg_18663_n_230 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_SL g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_0),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_14),
.Y(n_41)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_19),
.B1(n_20),
.B2(n_29),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_55),
.B1(n_17),
.B2(n_29),
.Y(n_71)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_52),
.Y(n_64)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_26),
.B1(n_31),
.B2(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_56),
.B(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_57),
.B(n_58),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_53),
.A2(n_41),
.B(n_40),
.C(n_38),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_78),
.Y(n_90)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g105 ( 
.A(n_63),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_41),
.B(n_32),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_18),
.B(n_32),
.Y(n_87)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_21),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_69),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_37),
.B1(n_20),
.B2(n_19),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_70),
.A2(n_18),
.B1(n_32),
.B2(n_25),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_76),
.B1(n_81),
.B2(n_83),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_80),
.Y(n_109)
);

NAND2x1_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_37),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_34),
.Y(n_93)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_17),
.B1(n_31),
.B2(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_39),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_28),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_42),
.A2(n_54),
.B1(n_49),
.B2(n_24),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_39),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_85),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_39),
.B1(n_34),
.B2(n_22),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_25),
.Y(n_125)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_95),
.B1(n_107),
.B2(n_79),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_60),
.A2(n_49),
.B1(n_26),
.B2(n_27),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_96),
.Y(n_126)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_18),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_27),
.B1(n_18),
.B2(n_32),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_77),
.B1(n_61),
.B2(n_74),
.Y(n_119)
);

INVx5_ASAP7_75t_SL g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_74),
.Y(n_120)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_59),
.A2(n_27),
.B1(n_32),
.B2(n_18),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_R g110 ( 
.A(n_99),
.B(n_58),
.C(n_73),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_96),
.B(n_93),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_65),
.C(n_57),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_27),
.C(n_30),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_125),
.B(n_132),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_73),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_107),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_118),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_117),
.B(n_122),
.Y(n_135)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_121),
.B1(n_123),
.B2(n_105),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_120),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_61),
.B1(n_66),
.B2(n_63),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_85),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_62),
.B1(n_75),
.B2(n_69),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_97),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_124),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_91),
.B(n_62),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_25),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_95),
.B(n_72),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_130),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_87),
.A2(n_25),
.B(n_23),
.C(n_64),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_98),
.Y(n_133)
);

INVx3_ASAP7_75t_SL g152 ( 
.A(n_133),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_30),
.C(n_2),
.Y(n_168)
);

XNOR2x1_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_93),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_1),
.B(n_2),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_145),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_88),
.B(n_108),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_147),
.B(n_148),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_143),
.B(n_151),
.C(n_4),
.Y(n_173)
);

AOI22x1_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_86),
.B1(n_101),
.B2(n_94),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_86),
.B1(n_105),
.B2(n_94),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_149),
.B1(n_30),
.B2(n_6),
.Y(n_171)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_88),
.A3(n_102),
.B1(n_105),
.B2(n_25),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_89),
.B(n_23),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_89),
.B(n_23),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_92),
.B1(n_64),
.B2(n_3),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_1),
.B(n_2),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_116),
.C(n_121),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_113),
.B1(n_111),
.B2(n_115),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_164),
.B1(n_168),
.B2(n_170),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_153),
.B(n_117),
.Y(n_160)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_146),
.C(n_155),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_111),
.B1(n_130),
.B2(n_131),
.Y(n_164)
);

BUFx12f_ASAP7_75t_SL g165 ( 
.A(n_137),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_148),
.B(n_146),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_118),
.Y(n_166)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_173),
.B(n_151),
.C(n_140),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_171),
.A2(n_172),
.B1(n_156),
.B2(n_154),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_6),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_188),
.B1(n_164),
.B2(n_170),
.Y(n_193)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_177),
.A2(n_158),
.B1(n_173),
.B2(n_149),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_157),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_173),
.B(n_145),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_147),
.C(n_139),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_183),
.B(n_186),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_162),
.B(n_165),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_136),
.C(n_154),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_173),
.A2(n_142),
.B1(n_134),
.B2(n_144),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_200),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_192),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_197),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_183),
.B(n_186),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_196),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_157),
.B(n_162),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_195),
.B(n_175),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_181),
.B(n_172),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_199),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_184),
.B(n_171),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_179),
.C(n_187),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_178),
.C(n_190),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_180),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_10),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_10),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_188),
.C(n_177),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_211),
.C(n_204),
.Y(n_219)
);

OAI21x1_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_7),
.B(n_9),
.Y(n_212)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_7),
.B(n_10),
.Y(n_213)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_203),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_215),
.B(n_206),
.Y(n_217)
);

AO21x1_ASAP7_75t_L g222 ( 
.A1(n_217),
.A2(n_216),
.B(n_214),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_220),
.B(n_210),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_222),
.B(n_224),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_218),
.A2(n_204),
.B(n_12),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_220),
.C(n_221),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_225),
.C(n_12),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_11),
.B1(n_13),
.B2(n_223),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_11),
.Y(n_230)
);


endmodule