module real_jpeg_11103_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_1),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_1),
.A2(n_57),
.B1(n_58),
.B2(n_70),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_1),
.A2(n_16),
.B(n_58),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_2),
.A2(n_57),
.B1(n_58),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_2),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_63),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_63),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_3),
.A2(n_68),
.B1(n_74),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_3),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_3),
.A2(n_57),
.B1(n_58),
.B2(n_91),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_91),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_91),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_4),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_42),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_5),
.A2(n_68),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_5),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_75),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_75),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_75),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_SL g35 ( 
.A1(n_8),
.A2(n_36),
.B(n_38),
.C(n_39),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_8),
.B(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_SL g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_11),
.A2(n_68),
.B1(n_74),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_11),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_11),
.A2(n_57),
.B1(n_58),
.B2(n_108),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_108),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_108),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_15),
.A2(n_68),
.B1(n_74),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_15),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_15),
.A2(n_57),
.B1(n_58),
.B2(n_77),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_15),
.A2(n_36),
.B1(n_37),
.B2(n_77),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_77),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_16),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_16),
.A2(n_68),
.B1(n_74),
.B2(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_16),
.B(n_134),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_16),
.A2(n_36),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_16),
.B(n_36),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_16),
.A2(n_26),
.B1(n_31),
.B2(n_187),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_16),
.A2(n_57),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_16),
.B(n_57),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_17),
.A2(n_36),
.B1(n_37),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_17),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_17),
.A2(n_29),
.B1(n_30),
.B2(n_52),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_119),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_117),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_95),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_21),
.B(n_95),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_81),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_46),
.B1(n_79),
.B2(n_80),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_23),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_34),
.B2(n_45),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B(n_32),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_26),
.A2(n_31),
.B1(n_49),
.B2(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_26),
.A2(n_31),
.B1(n_84),
.B2(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_26),
.A2(n_31),
.B1(n_170),
.B2(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_26),
.A2(n_31),
.B1(n_172),
.B2(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_26),
.A2(n_31),
.B1(n_203),
.B2(n_218),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_27),
.A2(n_28),
.B1(n_116),
.B2(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_27),
.A2(n_28),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_29),
.B(n_40),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_29),
.B(n_192),
.Y(n_191)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_30),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_31),
.B(n_112),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_39),
.B1(n_41),
.B2(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_35),
.A2(n_39),
.B1(n_51),
.B2(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_35),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_35),
.A2(n_39),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_35),
.A2(n_39),
.B1(n_178),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_35),
.A2(n_39),
.B1(n_201),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_35),
.A2(n_39),
.B1(n_137),
.B2(n_208),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_37),
.B1(n_56),
.B2(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_36),
.B(n_61),
.Y(n_215)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_37),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_38),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_39),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_39),
.B(n_112),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_46),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_53),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_50),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_65),
.B1(n_66),
.B2(n_78),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_62),
.B2(n_64),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_55),
.A2(n_60),
.B1(n_62),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_55),
.A2(n_60),
.B1(n_94),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_55),
.A2(n_60),
.B1(n_103),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_55),
.A2(n_60),
.B1(n_130),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_55),
.A2(n_60),
.B1(n_156),
.B2(n_210),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B(n_59),
.C(n_60),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_57),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_56),
.Y(n_61)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_59),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_60),
.B(n_112),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_72),
.B1(n_73),
.B2(n_76),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_67),
.A2(n_72),
.B1(n_73),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_67),
.A2(n_72),
.B1(n_90),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_70),
.B(n_71),
.C(n_72),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_70),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_68),
.A2(n_70),
.B(n_112),
.C(n_113),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_88),
.C(n_92),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_85),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_87),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.C(n_99),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_98),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_99),
.A2(n_100),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_104),
.C(n_109),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_114),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_161),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_143),
.B(n_160),
.Y(n_121)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_122),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_140),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_123),
.B(n_140),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.C(n_127),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_127),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.C(n_135),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_129),
.B1(n_135),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_135),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_144),
.B(n_146),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_152),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_147),
.B(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_150),
.A2(n_152),
.B1(n_153),
.B2(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_150),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_158),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_154),
.A2(n_155),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_157),
.B(n_158),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_159),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_240),
.C(n_241),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_234),
.B(n_239),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_220),
.B(n_233),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_205),
.B(n_219),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_195),
.B(n_204),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_184),
.B(n_194),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_173),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_168),
.B(n_173),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_179),
.B2(n_183),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_174),
.B(n_183),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_177),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_179),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_189),
.B(n_193),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_188),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_196),
.B(n_197),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_198),
.B(n_206),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_200),
.CI(n_202),
.CON(n_198),
.SN(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_206),
.Y(n_221)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.CI(n_212),
.CON(n_206),
.SN(n_206)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_211),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_217),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_221),
.B(n_222),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_227),
.B2(n_228),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_230),
.C(n_231),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_229),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_230),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_235),
.B(n_236),
.Y(n_239)
);


endmodule