module fake_jpeg_8257_n_274 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_34),
.Y(n_38)
);

HAxp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_43),
.CON(n_50),
.SN(n_50)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_45),
.Y(n_47)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_44),
.Y(n_46)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_71),
.Y(n_77)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_52),
.Y(n_75)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_64),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_21),
.B1(n_22),
.B2(n_31),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_62),
.B1(n_33),
.B2(n_39),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_21),
.B1(n_31),
.B2(n_22),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_56),
.A2(n_59),
.B1(n_60),
.B2(n_24),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_31),
.B1(n_20),
.B2(n_22),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_33),
.B(n_17),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_21),
.B1(n_25),
.B2(n_35),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_25),
.B1(n_35),
.B2(n_19),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_69),
.Y(n_83)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_41),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_26),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_32),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_80),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_73),
.A2(n_28),
.B(n_1),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_76),
.B(n_104),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_78),
.A2(n_106),
.B1(n_92),
.B2(n_80),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_36),
.B(n_30),
.C(n_29),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_79),
.A2(n_84),
.B(n_28),
.C(n_1),
.Y(n_125)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_81),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_82),
.A2(n_88),
.B1(n_91),
.B2(n_99),
.Y(n_131)
);

OR2x4_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_23),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_85),
.B(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_90),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_59),
.A2(n_39),
.B1(n_69),
.B2(n_36),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_47),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_60),
.A2(n_39),
.B1(n_41),
.B2(n_29),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_96),
.Y(n_132)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_97),
.Y(n_124)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_39),
.B1(n_30),
.B2(n_32),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_51),
.B(n_32),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_102),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_28),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_27),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_37),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_127),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_109),
.B(n_114),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_64),
.B1(n_24),
.B2(n_27),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_110),
.A2(n_126),
.B1(n_89),
.B2(n_12),
.Y(n_153)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_118),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_79),
.A2(n_26),
.B1(n_17),
.B2(n_28),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_113),
.B1(n_125),
.B2(n_119),
.Y(n_144)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_0),
.B(n_3),
.Y(n_141)
);

CKINVDCx10_ASAP7_75t_R g122 ( 
.A(n_72),
.Y(n_122)
);

INVx3_ASAP7_75t_SL g146 ( 
.A(n_122),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_122),
.B(n_87),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_125),
.B(n_3),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_82),
.A2(n_28),
.B1(n_15),
.B2(n_12),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_0),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_0),
.C(n_3),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_5),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_132),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_145),
.Y(n_172)
);

AO22x1_ASAP7_75t_SL g136 ( 
.A1(n_131),
.A2(n_91),
.B1(n_99),
.B2(n_96),
.Y(n_136)
);

AO22x1_ASAP7_75t_SL g185 ( 
.A1(n_136),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_77),
.B(n_101),
.C(n_81),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_137),
.A2(n_140),
.B(n_161),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_138),
.B(n_142),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_75),
.Y(n_139)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_160),
.B(n_121),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_89),
.Y(n_143)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_144),
.A2(n_162),
.B1(n_9),
.B2(n_11),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_107),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_156),
.Y(n_184)
);

INVx3_ASAP7_75t_SL g148 ( 
.A(n_124),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_124),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_158),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_92),
.B1(n_97),
.B2(n_87),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_151),
.A2(n_109),
.B1(n_128),
.B2(n_117),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_108),
.B(n_102),
.Y(n_154)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_155),
.B(n_157),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_105),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_113),
.B(n_15),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_105),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_130),
.B(n_6),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_168),
.B1(n_171),
.B2(n_181),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_164),
.B(n_141),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_150),
.C(n_152),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_167),
.C(n_153),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_115),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_147),
.A2(n_120),
.B1(n_117),
.B2(n_111),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_144),
.B(n_120),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_180),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_136),
.A2(n_112),
.B1(n_74),
.B2(n_133),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_93),
.B(n_112),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_175),
.A2(n_185),
.B(n_146),
.C(n_137),
.Y(n_199)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_178),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_148),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_149),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_162),
.A2(n_6),
.B(n_7),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_136),
.A2(n_74),
.B1(n_93),
.B2(n_10),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_178),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_190),
.B(n_193),
.Y(n_219)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_192),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_172),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_194),
.A2(n_205),
.B(n_206),
.Y(n_224)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_201),
.Y(n_213)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_199),
.A2(n_204),
.B(n_164),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_134),
.Y(n_200)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_161),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_184),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_202),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_208),
.C(n_155),
.Y(n_222)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_182),
.C(n_166),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_135),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_146),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_181),
.B1(n_171),
.B2(n_183),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_151),
.C(n_146),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_210),
.A2(n_199),
.B(n_190),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_215),
.A2(n_189),
.B(n_209),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_191),
.A2(n_185),
.B1(n_177),
.B2(n_175),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_216),
.A2(n_209),
.B1(n_195),
.B2(n_197),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_191),
.A2(n_163),
.B1(n_177),
.B2(n_142),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_218),
.B1(n_221),
.B2(n_192),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_187),
.B1(n_137),
.B2(n_180),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_199),
.A2(n_157),
.B1(n_160),
.B2(n_155),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_223),
.C(n_213),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_201),
.C(n_208),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_227),
.A2(n_229),
.B(n_238),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_196),
.Y(n_228)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_234),
.B(n_237),
.C(n_238),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_236),
.C(n_239),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_212),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_233),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_232),
.A2(n_217),
.B(n_218),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_219),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_229),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_159),
.C(n_11),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_159),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_220),
.B(n_11),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_240),
.B(n_221),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_241),
.Y(n_252)
);

AOI21x1_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_245),
.B(n_248),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_222),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_249),
.C(n_225),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_227),
.A2(n_224),
.B(n_226),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_247),
.A2(n_226),
.B(n_232),
.Y(n_251)
);

BUFx24_ASAP7_75t_SL g249 ( 
.A(n_228),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_253),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_242),
.B(n_236),
.Y(n_254)
);

NOR2xp67_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_255),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_243),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_231),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_262),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_259),
.A2(n_211),
.B(n_214),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_266),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_263),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_264),
.C(n_257),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

OA21x2_ASAP7_75t_SL g271 ( 
.A1(n_269),
.A2(n_258),
.B(n_212),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_271),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_268),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_245),
.Y(n_274)
);


endmodule