module fake_netlist_5_979_n_106 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_106);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_106;

wire n_91;
wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_96;
wire n_37;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_94;
wire n_38;
wire n_105;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_19;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_99;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_102;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVxp33_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

INVxp33_ASAP7_75t_SL g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_R g40 ( 
.A(n_33),
.B(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_24),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_25),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_33),
.B1(n_22),
.B2(n_24),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2x1p5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_25),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_53),
.A2(n_22),
.B1(n_38),
.B2(n_31),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_54),
.B(n_46),
.Y(n_60)
);

O2A1O1Ixp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_45),
.B(n_41),
.C(n_34),
.Y(n_61)
);

NAND2x1p5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_20),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_62),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_66),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_70),
.Y(n_74)
);

AOI211x1_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_68),
.B(n_19),
.C(n_40),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_71),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_79),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_80),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_90),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_89),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_87),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_92),
.Y(n_96)
);

OAI211xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_34),
.B(n_40),
.C(n_81),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_95),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_98)
);

OR3x1_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_93),
.C(n_94),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_85),
.C(n_55),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_96),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_102),
.Y(n_103)
);

NAND5xp2_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_100),
.C(n_69),
.D(n_85),
.E(n_17),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

AOI221xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_85),
.B1(n_55),
.B2(n_13),
.C(n_10),
.Y(n_106)
);


endmodule