module fake_netlist_6_1038_n_2934 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_625, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_628, n_557, n_349, n_233, n_617, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_327, n_369, n_597, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_621, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_612, n_633, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_110, n_151, n_412, n_640, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_528, n_391, n_457, n_364, n_637, n_295, n_385, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2934);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_625;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_233;
input n_617;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_612;
input n_633;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_637;
input n_295;
input n_385;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2934;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_2405;
wire n_1930;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_1371;
wire n_1285;
wire n_873;
wire n_2886;
wire n_1985;
wire n_2838;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_822;
wire n_693;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_1591;
wire n_772;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_2880;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_2843;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_699;
wire n_1986;
wire n_2300;
wire n_2397;
wire n_824;
wire n_686;
wire n_757;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_966;
wire n_2908;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_2922;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_2878;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_690;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2810;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_2916;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_2824;
wire n_697;
wire n_687;
wire n_890;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_840;
wire n_2913;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_794;
wire n_2767;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_1139;
wire n_872;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2643;
wire n_2590;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_765;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2307;
wire n_2069;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_2848;
wire n_919;
wire n_2868;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2896;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_745;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1475;
wire n_1774;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_683;
wire n_811;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_1837;
wire n_964;
wire n_831;
wire n_2218;
wire n_2788;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2301;
wire n_2209;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_2920;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_2863;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2830;
wire n_2781;
wire n_1129;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_1593;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_2841;
wire n_2420;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_2755;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2819;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_2439;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2900;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_2902;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2904;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_2872;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2882;
wire n_2541;
wire n_654;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_776;
wire n_1823;
wire n_2479;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_787;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_2840;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_2671;
wire n_2888;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_1804;
wire n_2923;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_2845;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_1476;
wire n_841;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_2587;
wire n_2931;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_814;
wire n_2746;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_2906;
wire n_1303;
wire n_761;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2858;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2255;
wire n_2112;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_908;
wire n_752;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_2743;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_2600;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_802;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2795;
wire n_2471;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_2879;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_2899;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_516),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_280),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_37),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_405),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_509),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_292),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_528),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_475),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_498),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_199),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_147),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_306),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_192),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_157),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_561),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_259),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_616),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_256),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_182),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_484),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_316),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_378),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_314),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_71),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_158),
.Y(n_665)
);

BUFx10_ASAP7_75t_L g666 ( 
.A(n_330),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_302),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_462),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_143),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_61),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_541),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_71),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_392),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_375),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_521),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_155),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_499),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_526),
.Y(n_678)
);

CKINVDCx14_ASAP7_75t_R g679 ( 
.A(n_485),
.Y(n_679)
);

BUFx2_ASAP7_75t_SL g680 ( 
.A(n_518),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_125),
.Y(n_681)
);

CKINVDCx14_ASAP7_75t_R g682 ( 
.A(n_519),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_382),
.Y(n_683)
);

CKINVDCx14_ASAP7_75t_R g684 ( 
.A(n_68),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_347),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_55),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_573),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_533),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_284),
.Y(n_689)
);

BUFx10_ASAP7_75t_L g690 ( 
.A(n_447),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_64),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_595),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_61),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_380),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_6),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_211),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_95),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_513),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_246),
.Y(n_699)
);

CKINVDCx14_ASAP7_75t_R g700 ( 
.A(n_522),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_214),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_22),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_527),
.Y(n_703)
);

BUFx2_ASAP7_75t_L g704 ( 
.A(n_204),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_483),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_110),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_498),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_274),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_501),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_15),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_626),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_530),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_273),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_73),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_552),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_117),
.Y(n_716)
);

BUFx10_ASAP7_75t_L g717 ( 
.A(n_20),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_555),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_494),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_184),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_110),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_151),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_266),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_397),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_144),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_121),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_277),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_58),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_40),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_281),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_185),
.Y(n_731)
);

INVx1_ASAP7_75t_SL g732 ( 
.A(n_551),
.Y(n_732)
);

BUFx5_ASAP7_75t_L g733 ( 
.A(n_254),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_133),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_146),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_31),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_19),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_501),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_271),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_376),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_318),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_24),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_275),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_398),
.Y(n_744)
);

BUFx10_ASAP7_75t_L g745 ( 
.A(n_109),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_196),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_459),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_540),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_45),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_381),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_441),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_8),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_554),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_11),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_90),
.Y(n_755)
);

BUFx8_ASAP7_75t_SL g756 ( 
.A(n_414),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_451),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_293),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_230),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_149),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_222),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_369),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_521),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_406),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_467),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_12),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_119),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_491),
.Y(n_768)
);

CKINVDCx14_ASAP7_75t_R g769 ( 
.A(n_230),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_405),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_213),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_562),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_559),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_430),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_342),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_16),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_133),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_454),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_270),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_426),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_82),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_136),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_484),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_313),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_459),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_283),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_56),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_204),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_379),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_444),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_154),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_143),
.Y(n_792)
);

CKINVDCx14_ASAP7_75t_R g793 ( 
.A(n_422),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_215),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_514),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_70),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_403),
.Y(n_797)
);

CKINVDCx14_ASAP7_75t_R g798 ( 
.A(n_520),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_366),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_82),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_15),
.Y(n_801)
);

BUFx10_ASAP7_75t_L g802 ( 
.A(n_151),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_190),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_617),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_141),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_463),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_89),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_192),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_533),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_29),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_13),
.Y(n_811)
);

CKINVDCx16_ASAP7_75t_R g812 ( 
.A(n_227),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_512),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_289),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_38),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_618),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_487),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_83),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_352),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_153),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_515),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_37),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_335),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_36),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_394),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_252),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_76),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_59),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_631),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_73),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_606),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_136),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_461),
.Y(n_833)
);

INVx1_ASAP7_75t_SL g834 ( 
.A(n_535),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_97),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_372),
.Y(n_836)
);

BUFx10_ASAP7_75t_L g837 ( 
.A(n_529),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_590),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_612),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_5),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_485),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_64),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_523),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_510),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_450),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_392),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_388),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_57),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_313),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_20),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_563),
.Y(n_851)
);

BUFx10_ASAP7_75t_L g852 ( 
.A(n_123),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_51),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_581),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_300),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_150),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_525),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_42),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_227),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_448),
.Y(n_860)
);

BUFx10_ASAP7_75t_L g861 ( 
.A(n_461),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_304),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_364),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_511),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_477),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_522),
.Y(n_866)
);

BUFx2_ASAP7_75t_SL g867 ( 
.A(n_293),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_281),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_510),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_148),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_75),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_341),
.Y(n_872)
);

BUFx10_ASAP7_75t_L g873 ( 
.A(n_524),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_261),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_508),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_117),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_183),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_94),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_296),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_634),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_517),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_270),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_425),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_543),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_594),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_282),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_112),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_145),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_47),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_613),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_733),
.Y(n_891)
);

INVxp33_ASAP7_75t_L g892 ( 
.A(n_704),
.Y(n_892)
);

INVxp67_ASAP7_75t_SL g893 ( 
.A(n_715),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_756),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_756),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_647),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_733),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_890),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_733),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_679),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_679),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_733),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_733),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_682),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_890),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_682),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_647),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_684),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_684),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_773),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_719),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_733),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_653),
.Y(n_913)
);

INVxp33_ASAP7_75t_L g914 ( 
.A(n_778),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_733),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_699),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_699),
.Y(n_917)
);

NOR2xp67_ASAP7_75t_L g918 ( 
.A(n_699),
.B(n_0),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_648),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_700),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_648),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_709),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_772),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_709),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_700),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_710),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_644),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_710),
.Y(n_928)
);

INVxp67_ASAP7_75t_SL g929 ( 
.A(n_838),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_773),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_723),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_653),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_723),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_737),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_737),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_762),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_762),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_799),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_799),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_824),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_769),
.B(n_1),
.Y(n_941)
);

BUFx10_ASAP7_75t_L g942 ( 
.A(n_644),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_824),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_829),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_850),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_644),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_850),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_812),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_769),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_644),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_765),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_765),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_655),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_793),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_765),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_765),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_830),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_830),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_830),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_793),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_666),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_798),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_830),
.Y(n_963)
);

BUFx3_ASAP7_75t_L g964 ( 
.A(n_831),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_888),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_888),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_676),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_888),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_798),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_888),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_643),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_839),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_666),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_676),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_649),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_674),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_641),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_650),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_686),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_651),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_656),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_642),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_661),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_667),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_686),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_672),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_645),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_673),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_674),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_683),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_851),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_678),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_683),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_646),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_953),
.B(n_657),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_894),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_950),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_952),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_948),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_898),
.B(n_697),
.Y(n_1000)
);

CKINVDCx16_ASAP7_75t_R g1001 ( 
.A(n_895),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_956),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_894),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_957),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_927),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_905),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_896),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_927),
.Y(n_1008)
);

CKINVDCx20_ASAP7_75t_R g1009 ( 
.A(n_896),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_982),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_946),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_946),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_982),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_900),
.B(n_732),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_898),
.B(n_851),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_907),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_951),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_951),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_959),
.Y(n_1019)
);

INVxp67_ASAP7_75t_SL g1020 ( 
.A(n_905),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_963),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_895),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_965),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_966),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_955),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_968),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_970),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_987),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_987),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_955),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_958),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_958),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_994),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_994),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_893),
.B(n_929),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_900),
.B(n_718),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_910),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_961),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_901),
.B(n_804),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_976),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_977),
.Y(n_1041)
);

INVxp67_ASAP7_75t_SL g1042 ( 
.A(n_905),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_910),
.Y(n_1043)
);

XOR2xp5_ASAP7_75t_L g1044 ( 
.A(n_907),
.B(n_913),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_901),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_913),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_954),
.B(n_697),
.Y(n_1047)
);

INVxp33_ASAP7_75t_L g1048 ( 
.A(n_892),
.Y(n_1048)
);

INVxp67_ASAP7_75t_SL g1049 ( 
.A(n_905),
.Y(n_1049)
);

CKINVDCx11_ASAP7_75t_R g1050 ( 
.A(n_932),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_976),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_904),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_989),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_932),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_904),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_906),
.B(n_880),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_910),
.Y(n_1057)
);

CKINVDCx16_ASAP7_75t_R g1058 ( 
.A(n_967),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_989),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_990),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_910),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_997),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_995),
.B(n_906),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1014),
.A2(n_941),
.B1(n_908),
.B2(n_920),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_1015),
.A2(n_897),
.B(n_891),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1020),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_1006),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1042),
.B(n_908),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1049),
.B(n_909),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_1025),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1006),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1000),
.B(n_917),
.Y(n_1072)
);

OAI22x1_ASAP7_75t_R g1073 ( 
.A1(n_1001),
.A2(n_974),
.B1(n_979),
.B2(n_967),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1037),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_999),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1000),
.B(n_916),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_SL g1077 ( 
.A1(n_1058),
.A2(n_695),
.B1(n_758),
.B2(n_740),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_998),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1025),
.Y(n_1079)
);

INVxp33_ASAP7_75t_SL g1080 ( 
.A(n_1038),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_1002),
.B(n_916),
.Y(n_1081)
);

OA21x2_ASAP7_75t_L g1082 ( 
.A1(n_1030),
.A2(n_902),
.B(n_899),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1004),
.B(n_918),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_1043),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1031),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_1019),
.B(n_990),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_1057),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1056),
.B(n_993),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1021),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_1061),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1032),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1047),
.A2(n_909),
.B1(n_925),
.B2(n_920),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1023),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_1041),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_1048),
.Y(n_1095)
);

BUFx8_ASAP7_75t_L g1096 ( 
.A(n_1055),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_SL g1097 ( 
.A(n_1052),
.B(n_816),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1040),
.B(n_993),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_1047),
.A2(n_949),
.B1(n_960),
.B2(n_925),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_1005),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_1024),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1005),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1040),
.B(n_923),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_1026),
.Y(n_1104)
);

OA21x2_ASAP7_75t_L g1105 ( 
.A1(n_1008),
.A2(n_912),
.B(n_903),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1036),
.B(n_962),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1027),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1008),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1011),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1051),
.B(n_923),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1039),
.B(n_949),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_1055),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1011),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_1050),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1051),
.B(n_944),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_SL g1116 ( 
.A1(n_1007),
.A2(n_695),
.B1(n_758),
.B2(n_740),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_1012),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1012),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_1017),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1017),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1018),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1018),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1053),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_1053),
.B(n_971),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1059),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1059),
.B(n_944),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1060),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1035),
.A2(n_915),
.B(n_880),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1060),
.B(n_962),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1045),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1044),
.A2(n_921),
.B(n_919),
.Y(n_1131)
);

OAI22x1_ASAP7_75t_R g1132 ( 
.A1(n_1009),
.A2(n_979),
.B1(n_985),
.B2(n_974),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1052),
.Y(n_1133)
);

CKINVDCx14_ASAP7_75t_R g1134 ( 
.A(n_1016),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1010),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1010),
.B(n_975),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1013),
.A2(n_969),
.B1(n_960),
.B2(n_911),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1013),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_1028),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1028),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_1046),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_1029),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1029),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1033),
.B(n_969),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1033),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1034),
.B(n_973),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1034),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_996),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_996),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1003),
.B(n_930),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_1095),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1114),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_1114),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_R g1154 ( 
.A(n_1134),
.B(n_1003),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_1067),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1100),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_1141),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_1067),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_1080),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1080),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1100),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1075),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1063),
.B(n_1106),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1075),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1062),
.Y(n_1165)
);

INVx4_ASAP7_75t_L g1166 ( 
.A(n_1067),
.Y(n_1166)
);

INVxp67_ASAP7_75t_L g1167 ( 
.A(n_1097),
.Y(n_1167)
);

INVxp33_ASAP7_75t_L g1168 ( 
.A(n_1132),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1102),
.Y(n_1169)
);

INVxp67_ASAP7_75t_L g1170 ( 
.A(n_1094),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1139),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_1139),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1139),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1081),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1094),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_1141),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1102),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_R g1178 ( 
.A(n_1148),
.B(n_1054),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_R g1179 ( 
.A(n_1148),
.B(n_985),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_1112),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1136),
.B(n_816),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1088),
.B(n_930),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1062),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1067),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_R g1185 ( 
.A(n_1148),
.B(n_1022),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1078),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_1139),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_1139),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_1096),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1081),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1111),
.B(n_914),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1078),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_1096),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_R g1194 ( 
.A(n_1149),
.B(n_671),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1089),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1089),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1093),
.Y(n_1197)
);

INVx2_ASAP7_75t_SL g1198 ( 
.A(n_1088),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1108),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1133),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1133),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_1136),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1093),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1081),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1124),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1136),
.Y(n_1206)
);

INVxp67_ASAP7_75t_SL g1207 ( 
.A(n_1117),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1108),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1118),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_1133),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1133),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1133),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1118),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1096),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1124),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1124),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1145),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1070),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1142),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1142),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_R g1221 ( 
.A(n_1149),
.B(n_687),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1065),
.A2(n_980),
.B(n_978),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_1073),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_R g1224 ( 
.A(n_1135),
.B(n_692),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1070),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1120),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1120),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1103),
.Y(n_1228)
);

CKINVDCx6p67_ASAP7_75t_R g1229 ( 
.A(n_1142),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_R g1230 ( 
.A(n_1135),
.B(n_1138),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1142),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1142),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_1144),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1137),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1103),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1064),
.Y(n_1236)
);

CKINVDCx20_ASAP7_75t_R g1237 ( 
.A(n_1077),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1110),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1131),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_R g1240 ( 
.A(n_1138),
.B(n_1140),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1121),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1121),
.Y(n_1242)
);

BUFx10_ASAP7_75t_L g1243 ( 
.A(n_1140),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1067),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_R g1245 ( 
.A(n_1143),
.B(n_711),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1143),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1086),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1147),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1110),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1147),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1150),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1092),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1099),
.B(n_1044),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1109),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1116),
.Y(n_1255)
);

NAND2xp33_ASAP7_75t_SL g1256 ( 
.A(n_1146),
.B(n_1130),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1115),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1129),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_1068),
.Y(n_1259)
);

BUFx10_ASAP7_75t_L g1260 ( 
.A(n_1083),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_1069),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1076),
.B(n_973),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1107),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_1072),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1115),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1126),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1086),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1076),
.B(n_922),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1066),
.B(n_930),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1083),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1086),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_R g1272 ( 
.A(n_1071),
.B(n_748),
.Y(n_1272)
);

NAND2xp33_ASAP7_75t_R g1273 ( 
.A(n_1131),
.B(n_652),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_1072),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1083),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1079),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1126),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_1074),
.Y(n_1278)
);

NOR2xp67_ASAP7_75t_L g1279 ( 
.A(n_1125),
.B(n_924),
.Y(n_1279)
);

CKINVDCx20_ASAP7_75t_R g1280 ( 
.A(n_1123),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1123),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1127),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1101),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1101),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1127),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1101),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1098),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1098),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1163),
.B(n_1101),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1205),
.Y(n_1290)
);

INVx4_ASAP7_75t_L g1291 ( 
.A(n_1171),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1254),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1254),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1191),
.B(n_926),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1155),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1205),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1163),
.B(n_1101),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1162),
.Y(n_1298)
);

AND2x2_ASAP7_75t_SL g1299 ( 
.A(n_1253),
.B(n_701),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1198),
.B(n_1251),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1247),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1191),
.B(n_1104),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1156),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1258),
.B(n_1104),
.Y(n_1304)
);

AND2x6_ASAP7_75t_L g1305 ( 
.A(n_1262),
.B(n_1109),
.Y(n_1305)
);

AND2x6_ASAP7_75t_L g1306 ( 
.A(n_1215),
.B(n_1113),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1156),
.Y(n_1307)
);

OR2x6_ASAP7_75t_L g1308 ( 
.A(n_1206),
.B(n_680),
.Y(n_1308)
);

AND2x6_ASAP7_75t_L g1309 ( 
.A(n_1216),
.B(n_1113),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_1175),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1247),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1267),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1267),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1155),
.Y(n_1314)
);

INVx4_ASAP7_75t_L g1315 ( 
.A(n_1172),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1182),
.B(n_1281),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1271),
.Y(n_1317)
);

AND2x6_ASAP7_75t_L g1318 ( 
.A(n_1228),
.B(n_1119),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1151),
.Y(n_1319)
);

INVx4_ASAP7_75t_L g1320 ( 
.A(n_1173),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1271),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1170),
.B(n_928),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1161),
.Y(n_1323)
);

AND2x6_ASAP7_75t_L g1324 ( 
.A(n_1235),
.B(n_1119),
.Y(n_1324)
);

NAND2xp33_ASAP7_75t_L g1325 ( 
.A(n_1187),
.B(n_1104),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1169),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1174),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1157),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1174),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1188),
.B(n_1104),
.Y(n_1330)
);

INVx1_ASAP7_75t_SL g1331 ( 
.A(n_1264),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1285),
.B(n_1105),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1239),
.A2(n_1104),
.B1(n_1084),
.B2(n_1090),
.Y(n_1333)
);

INVx4_ASAP7_75t_L g1334 ( 
.A(n_1200),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1180),
.B(n_1164),
.Y(n_1335)
);

AND2x6_ASAP7_75t_L g1336 ( 
.A(n_1238),
.B(n_1119),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1287),
.B(n_1105),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1277),
.B(n_1085),
.Y(n_1338)
);

INVx6_ASAP7_75t_L g1339 ( 
.A(n_1260),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1202),
.A2(n_1257),
.B1(n_1265),
.B2(n_1249),
.Y(n_1340)
);

INVx4_ASAP7_75t_L g1341 ( 
.A(n_1201),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1288),
.A2(n_1105),
.B1(n_1082),
.B2(n_726),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1165),
.B(n_1105),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1183),
.B(n_1082),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1246),
.B(n_760),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1190),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1274),
.Y(n_1347)
);

AND2x6_ASAP7_75t_L g1348 ( 
.A(n_1266),
.B(n_1085),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1169),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1177),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1186),
.B(n_1082),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1176),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1177),
.A2(n_1082),
.B1(n_726),
.B2(n_712),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1204),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1199),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1199),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1236),
.A2(n_760),
.B1(n_788),
.B2(n_766),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1210),
.B(n_1091),
.Y(n_1358)
);

OR2x2_ASAP7_75t_SL g1359 ( 
.A(n_1237),
.B(n_701),
.Y(n_1359)
);

XOR2xp5_ASAP7_75t_R g1360 ( 
.A(n_1154),
.B(n_0),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1208),
.A2(n_795),
.B1(n_815),
.B2(n_712),
.Y(n_1361)
);

INVx4_ASAP7_75t_L g1362 ( 
.A(n_1211),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1167),
.B(n_1084),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_SL g1364 ( 
.A(n_1212),
.B(n_1091),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1192),
.B(n_1084),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1208),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1209),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1280),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1155),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1209),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1268),
.B(n_931),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1204),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1213),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1195),
.B(n_1090),
.Y(n_1374)
);

NAND2xp33_ASAP7_75t_L g1375 ( 
.A(n_1283),
.B(n_1087),
.Y(n_1375)
);

BUFx10_ASAP7_75t_L g1376 ( 
.A(n_1152),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1244),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1213),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_L g1379 ( 
.A(n_1196),
.B(n_1090),
.C(n_1117),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1226),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1226),
.Y(n_1381)
);

INVx4_ASAP7_75t_L g1382 ( 
.A(n_1284),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1227),
.A2(n_815),
.B1(n_820),
.B2(n_795),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1263),
.B(n_933),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1278),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1227),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1241),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1181),
.B(n_934),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_1282),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1179),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1241),
.A2(n_876),
.B1(n_820),
.B2(n_698),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1286),
.B(n_1087),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1242),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1242),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1244),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1248),
.B(n_766),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1218),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1250),
.B(n_788),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1197),
.B(n_1079),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1203),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1225),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1243),
.B(n_935),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1276),
.A2(n_876),
.B1(n_702),
.B2(n_703),
.Y(n_1403)
);

INVx6_ASAP7_75t_L g1404 ( 
.A(n_1260),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1207),
.B(n_1065),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_SL g1406 ( 
.A(n_1230),
.B(n_1087),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1179),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1269),
.B(n_1128),
.Y(n_1408)
);

AND2x2_ASAP7_75t_SL g1409 ( 
.A(n_1168),
.B(n_691),
.Y(n_1409)
);

BUFx10_ASAP7_75t_L g1410 ( 
.A(n_1153),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1222),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1158),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1243),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1158),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1279),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1259),
.B(n_789),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1158),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1230),
.B(n_1087),
.Y(n_1418)
);

BUFx10_ASAP7_75t_L g1419 ( 
.A(n_1159),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1160),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1158),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1184),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1219),
.B(n_1128),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1270),
.B(n_981),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1178),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1240),
.B(n_1087),
.Y(n_1426)
);

INVxp67_ASAP7_75t_SL g1427 ( 
.A(n_1184),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1217),
.B(n_789),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1240),
.B(n_753),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1184),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1220),
.B(n_1117),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1185),
.B(n_945),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1184),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1166),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1231),
.B(n_1117),
.Y(n_1435)
);

INVx4_ASAP7_75t_L g1436 ( 
.A(n_1229),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1166),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1275),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1232),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1194),
.B(n_854),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1252),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1261),
.B(n_1117),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1255),
.A2(n_706),
.B1(n_720),
.B2(n_716),
.Y(n_1443)
);

BUFx8_ASAP7_75t_SL g1444 ( 
.A(n_1223),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1185),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1233),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1234),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1194),
.B(n_884),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1178),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1272),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1221),
.B(n_1122),
.Y(n_1451)
);

BUFx10_ASAP7_75t_L g1452 ( 
.A(n_1214),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1221),
.B(n_885),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1256),
.B(n_821),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1189),
.B(n_983),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1272),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1224),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1224),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1273),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1245),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1245),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1273),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1154),
.Y(n_1463)
);

INVx4_ASAP7_75t_SL g1464 ( 
.A(n_1193),
.Y(n_1464)
);

AND2x6_ASAP7_75t_L g1465 ( 
.A(n_1262),
.B(n_1122),
.Y(n_1465)
);

NAND2xp33_ASAP7_75t_L g1466 ( 
.A(n_1171),
.B(n_1122),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1175),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1154),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1205),
.Y(n_1469)
);

AND2x2_ASAP7_75t_SL g1470 ( 
.A(n_1253),
.B(n_722),
.Y(n_1470)
);

NAND2xp33_ASAP7_75t_L g1471 ( 
.A(n_1171),
.B(n_1122),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1163),
.B(n_1122),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1163),
.B(n_821),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_SL g1474 ( 
.A(n_1251),
.B(n_964),
.Y(n_1474)
);

BUFx4f_ASAP7_75t_L g1475 ( 
.A(n_1206),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1254),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1254),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1191),
.B(n_936),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1254),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1254),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1163),
.B(n_855),
.Y(n_1481)
);

AO22x2_ASAP7_75t_L g1482 ( 
.A1(n_1181),
.A2(n_867),
.B1(n_796),
.B2(n_832),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1163),
.B(n_930),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1191),
.B(n_940),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1277),
.B(n_984),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1163),
.B(n_855),
.Y(n_1486)
);

NAND2xp33_ASAP7_75t_SL g1487 ( 
.A(n_1171),
.B(n_654),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1456),
.B(n_964),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1289),
.B(n_972),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1297),
.B(n_991),
.Y(n_1490)
);

INVx8_ASAP7_75t_L g1491 ( 
.A(n_1306),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1476),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1477),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1456),
.B(n_972),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1297),
.B(n_991),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1456),
.B(n_937),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1460),
.B(n_938),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1473),
.B(n_693),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1480),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1472),
.B(n_787),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1473),
.A2(n_988),
.B1(n_992),
.B2(n_986),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1472),
.B(n_783),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1460),
.B(n_939),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1481),
.B(n_792),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1316),
.B(n_819),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1292),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1316),
.B(n_834),
.Y(n_1507)
);

NAND3xp33_ASAP7_75t_L g1508 ( 
.A(n_1481),
.B(n_1486),
.C(n_1396),
.Y(n_1508)
);

CKINVDCx20_ASAP7_75t_R g1509 ( 
.A(n_1468),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1486),
.B(n_658),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_1384),
.Y(n_1511)
);

INVx2_ASAP7_75t_SL g1512 ( 
.A(n_1319),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1293),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1331),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1479),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1294),
.B(n_1478),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1302),
.B(n_659),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1303),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1459),
.A2(n_947),
.B1(n_943),
.B2(n_662),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1443),
.A2(n_725),
.B1(n_729),
.B2(n_724),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1445),
.B(n_660),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1445),
.B(n_663),
.Y(n_1522)
);

NAND3xp33_ASAP7_75t_L g1523 ( 
.A(n_1345),
.B(n_665),
.C(n_664),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1400),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1302),
.B(n_668),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1484),
.B(n_669),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1432),
.B(n_666),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1378),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1300),
.B(n_670),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1304),
.B(n_675),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1483),
.B(n_677),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1307),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1380),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1483),
.B(n_681),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1300),
.B(n_685),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1450),
.B(n_688),
.Y(n_1536)
);

AND3x1_ASAP7_75t_L g1537 ( 
.A(n_1398),
.B(n_734),
.C(n_730),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1457),
.B(n_689),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1462),
.A2(n_694),
.B1(n_705),
.B2(n_696),
.Y(n_1539)
);

BUFx6f_ASAP7_75t_SL g1540 ( 
.A(n_1376),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_SL g1541 ( 
.A(n_1376),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1386),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1371),
.B(n_707),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1387),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1363),
.B(n_708),
.Y(n_1545)
);

INVxp67_ASAP7_75t_SL g1546 ( 
.A(n_1427),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1467),
.Y(n_1547)
);

AND2x2_ASAP7_75t_SL g1548 ( 
.A(n_1470),
.B(n_735),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1410),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1363),
.B(n_739),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1337),
.B(n_741),
.Y(n_1551)
);

NAND2xp33_ASAP7_75t_L g1552 ( 
.A(n_1305),
.B(n_881),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1310),
.B(n_713),
.Y(n_1553)
);

NOR2xp67_ASAP7_75t_L g1554 ( 
.A(n_1291),
.B(n_537),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1299),
.B(n_690),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1305),
.B(n_714),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1305),
.B(n_721),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1410),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1377),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1393),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1402),
.B(n_690),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1331),
.B(n_727),
.Y(n_1562)
);

AOI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1441),
.A2(n_1461),
.B1(n_1458),
.B2(n_1442),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1323),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1310),
.B(n_728),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_SL g1566 ( 
.A(n_1291),
.B(n_690),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1441),
.B(n_731),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1485),
.B(n_1447),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1446),
.B(n_736),
.Y(n_1569)
);

OAI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1442),
.A2(n_738),
.B1(n_746),
.B2(n_743),
.Y(n_1570)
);

INVx2_ASAP7_75t_SL g1571 ( 
.A(n_1335),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1337),
.B(n_742),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1326),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1349),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1382),
.B(n_749),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1382),
.B(n_750),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1454),
.B(n_752),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1428),
.B(n_754),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1305),
.B(n_744),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1350),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1347),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1394),
.Y(n_1582)
);

NAND2xp33_ASAP7_75t_SL g1583 ( 
.A(n_1447),
.B(n_755),
.Y(n_1583)
);

NOR3xp33_ASAP7_75t_L g1584 ( 
.A(n_1416),
.B(n_761),
.C(n_759),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1338),
.B(n_763),
.Y(n_1585)
);

INVxp67_ASAP7_75t_L g1586 ( 
.A(n_1347),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1358),
.A2(n_1364),
.B1(n_1338),
.B2(n_1415),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1399),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1355),
.Y(n_1589)
);

NOR3xp33_ASAP7_75t_L g1590 ( 
.A(n_1416),
.B(n_771),
.C(n_764),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1385),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1315),
.B(n_774),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1399),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1340),
.B(n_775),
.Y(n_1594)
);

BUFx5_ASAP7_75t_L g1595 ( 
.A(n_1318),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1321),
.B(n_776),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_L g1597 ( 
.A(n_1295),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_L g1598 ( 
.A(n_1295),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1321),
.B(n_1327),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1356),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1327),
.B(n_780),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1366),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1329),
.B(n_781),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1329),
.B(n_784),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1315),
.B(n_785),
.Y(n_1605)
);

A2O1A1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1301),
.A2(n_751),
.B(n_757),
.C(n_747),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1367),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1370),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1320),
.B(n_786),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1372),
.B(n_790),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1373),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1485),
.B(n_717),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1381),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1320),
.B(n_797),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1334),
.B(n_801),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1328),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1372),
.B(n_803),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_L g1618 ( 
.A(n_1465),
.B(n_1318),
.Y(n_1618)
);

INVxp33_ASAP7_75t_L g1619 ( 
.A(n_1298),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1290),
.B(n_806),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1334),
.B(n_807),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1290),
.B(n_808),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1341),
.B(n_810),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1474),
.A2(n_814),
.B1(n_817),
.B2(n_811),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1352),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_1420),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1341),
.B(n_1362),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1397),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1401),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1362),
.B(n_818),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1482),
.A2(n_1312),
.B1(n_1313),
.B2(n_1311),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1317),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1447),
.B(n_823),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1424),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1368),
.B(n_826),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1296),
.B(n_827),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1296),
.B(n_833),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1346),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1475),
.B(n_717),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1469),
.B(n_835),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1368),
.B(n_840),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1389),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1475),
.B(n_841),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1439),
.B(n_842),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1469),
.B(n_843),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1424),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1482),
.B(n_844),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1482),
.B(n_845),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1389),
.B(n_1407),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1354),
.Y(n_1650)
);

NOR2xp67_ASAP7_75t_L g1651 ( 
.A(n_1436),
.B(n_538),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1444),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1377),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1322),
.B(n_846),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1395),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1407),
.B(n_847),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1365),
.B(n_848),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1413),
.B(n_857),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1365),
.B(n_859),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1374),
.B(n_860),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1388),
.B(n_862),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1374),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1487),
.A2(n_864),
.B1(n_868),
.B2(n_863),
.Y(n_1663)
);

INVxp33_ASAP7_75t_L g1664 ( 
.A(n_1449),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1417),
.Y(n_1665)
);

A2O1A1Ixp33_ASAP7_75t_L g1666 ( 
.A1(n_1451),
.A2(n_1379),
.B(n_1325),
.C(n_1330),
.Y(n_1666)
);

BUFx5_ASAP7_75t_L g1667 ( 
.A(n_1318),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1451),
.B(n_869),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1295),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1395),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1427),
.B(n_871),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1314),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1438),
.B(n_874),
.Y(n_1673)
);

BUFx3_ASAP7_75t_L g1674 ( 
.A(n_1419),
.Y(n_1674)
);

NAND2xp33_ASAP7_75t_SL g1675 ( 
.A(n_1436),
.B(n_875),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1465),
.B(n_877),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1343),
.B(n_1351),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1343),
.B(n_767),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1425),
.B(n_878),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1449),
.B(n_882),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1344),
.B(n_768),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1390),
.B(n_883),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1443),
.A2(n_777),
.B1(n_779),
.B2(n_770),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1463),
.B(n_887),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_SL g1685 ( 
.A(n_1314),
.B(n_1369),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1412),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1344),
.B(n_782),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1351),
.B(n_791),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1433),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1429),
.B(n_717),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1332),
.B(n_794),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1314),
.B(n_745),
.Y(n_1692)
);

BUFx2_ASAP7_75t_L g1693 ( 
.A(n_1308),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1524),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1518),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1568),
.B(n_1464),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_SL g1697 ( 
.A(n_1548),
.B(n_1409),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1532),
.Y(n_1698)
);

NAND2x1p5_ASAP7_75t_L g1699 ( 
.A(n_1626),
.B(n_1369),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1528),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1642),
.Y(n_1701)
);

AO22x2_ASAP7_75t_L g1702 ( 
.A1(n_1508),
.A2(n_1357),
.B1(n_1464),
.B2(n_1423),
.Y(n_1702)
);

AO22x2_ASAP7_75t_L g1703 ( 
.A1(n_1647),
.A2(n_1357),
.B1(n_1464),
.B2(n_1423),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1533),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1542),
.Y(n_1705)
);

AO22x2_ASAP7_75t_L g1706 ( 
.A1(n_1648),
.A2(n_1411),
.B1(n_1379),
.B2(n_1360),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1516),
.B(n_1308),
.Y(n_1707)
);

BUFx2_ASAP7_75t_L g1708 ( 
.A(n_1581),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1544),
.Y(n_1709)
);

AO22x2_ASAP7_75t_L g1710 ( 
.A1(n_1555),
.A2(n_1405),
.B1(n_1418),
.B2(n_1406),
.Y(n_1710)
);

OAI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1498),
.A2(n_1308),
.B1(n_1448),
.B2(n_1453),
.C(n_1440),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1527),
.B(n_1419),
.Y(n_1712)
);

AO22x2_ASAP7_75t_L g1713 ( 
.A1(n_1510),
.A2(n_1405),
.B1(n_1426),
.B2(n_1455),
.Y(n_1713)
);

NAND2x1p5_ASAP7_75t_L g1714 ( 
.A(n_1512),
.B(n_1369),
.Y(n_1714)
);

AO22x2_ASAP7_75t_L g1715 ( 
.A1(n_1584),
.A2(n_1455),
.B1(n_1392),
.B2(n_1408),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1504),
.B(n_1465),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1564),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1573),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1561),
.B(n_1511),
.Y(n_1719)
);

OAI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1577),
.A2(n_1403),
.B1(n_1391),
.B2(n_1383),
.C(n_1361),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1571),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1574),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1560),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1616),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1582),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1492),
.Y(n_1726)
);

AO22x2_ASAP7_75t_L g1727 ( 
.A1(n_1590),
.A2(n_1520),
.B1(n_1683),
.B2(n_1514),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1514),
.B(n_1452),
.Y(n_1728)
);

NAND2x1p5_ASAP7_75t_L g1729 ( 
.A(n_1547),
.B(n_1422),
.Y(n_1729)
);

NAND2x1p5_ASAP7_75t_L g1730 ( 
.A(n_1625),
.B(n_1422),
.Y(n_1730)
);

AO22x2_ASAP7_75t_L g1731 ( 
.A1(n_1520),
.A2(n_1408),
.B1(n_800),
.B2(n_809),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1580),
.Y(n_1732)
);

AND2x6_ASAP7_75t_L g1733 ( 
.A(n_1588),
.B(n_1422),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1589),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1493),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1499),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1600),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1608),
.Y(n_1738)
);

AOI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1578),
.A2(n_1465),
.B1(n_1309),
.B2(n_1306),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1611),
.Y(n_1740)
);

BUFx8_ASAP7_75t_L g1741 ( 
.A(n_1540),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1591),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1613),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1563),
.B(n_1452),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1513),
.Y(n_1745)
);

NAND2x1p5_ASAP7_75t_L g1746 ( 
.A(n_1674),
.B(n_1434),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1646),
.B(n_1339),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1515),
.Y(n_1748)
);

OAI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1690),
.A2(n_1403),
.B1(n_1391),
.B2(n_1383),
.C(n_1361),
.Y(n_1749)
);

INVx3_ASAP7_75t_L g1750 ( 
.A(n_1540),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1602),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1607),
.Y(n_1752)
);

AO22x2_ASAP7_75t_L g1753 ( 
.A1(n_1683),
.A2(n_813),
.B1(n_822),
.B2(n_805),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1506),
.Y(n_1754)
);

OA22x2_ASAP7_75t_L g1755 ( 
.A1(n_1587),
.A2(n_1359),
.B1(n_1333),
.B2(n_828),
.Y(n_1755)
);

AO22x2_ASAP7_75t_L g1756 ( 
.A1(n_1523),
.A2(n_836),
.B1(n_849),
.B2(n_825),
.Y(n_1756)
);

AO22x2_ASAP7_75t_L g1757 ( 
.A1(n_1502),
.A2(n_856),
.B1(n_858),
.B2(n_853),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1546),
.A2(n_1435),
.B1(n_1431),
.B2(n_1437),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1628),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1629),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1633),
.A2(n_1309),
.B1(n_1306),
.B2(n_1339),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1632),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1612),
.B(n_1339),
.Y(n_1763)
);

INVxp67_ASAP7_75t_L g1764 ( 
.A(n_1649),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1567),
.A2(n_1309),
.B1(n_1306),
.B2(n_1404),
.Y(n_1765)
);

AO22x2_ASAP7_75t_L g1766 ( 
.A1(n_1502),
.A2(n_866),
.B1(n_870),
.B2(n_865),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1566),
.B(n_1431),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1509),
.Y(n_1768)
);

OAI221xp5_ASAP7_75t_L g1769 ( 
.A1(n_1537),
.A2(n_1404),
.B1(n_1471),
.B2(n_1466),
.C(n_886),
.Y(n_1769)
);

AND2x6_ASAP7_75t_L g1770 ( 
.A(n_1593),
.B(n_1414),
.Y(n_1770)
);

AO22x2_ASAP7_75t_L g1771 ( 
.A1(n_1550),
.A2(n_879),
.B1(n_889),
.B2(n_872),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1638),
.Y(n_1772)
);

AO22x2_ASAP7_75t_L g1773 ( 
.A1(n_1550),
.A2(n_1332),
.B1(n_1430),
.B2(n_1421),
.Y(n_1773)
);

OAI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1543),
.A2(n_1404),
.B1(n_1435),
.B2(n_1375),
.C(n_1353),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1665),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1650),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1689),
.Y(n_1777)
);

CKINVDCx20_ASAP7_75t_R g1778 ( 
.A(n_1652),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1566),
.B(n_1353),
.Y(n_1779)
);

AO22x2_ASAP7_75t_L g1780 ( 
.A1(n_1500),
.A2(n_1348),
.B1(n_802),
.B2(n_837),
.Y(n_1780)
);

AO22x2_ASAP7_75t_L g1781 ( 
.A1(n_1500),
.A2(n_1662),
.B1(n_1579),
.B2(n_1586),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1686),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1505),
.B(n_1348),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1653),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1655),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1634),
.B(n_1309),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1505),
.B(n_1348),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1635),
.A2(n_1348),
.B1(n_1324),
.B2(n_1336),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1641),
.A2(n_1324),
.B1(n_1336),
.B2(n_1318),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1627),
.B(n_1324),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1507),
.B(n_1324),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1559),
.Y(n_1792)
);

OR2x2_ASAP7_75t_SL g1793 ( 
.A(n_1594),
.B(n_745),
.Y(n_1793)
);

NAND2x1p5_ASAP7_75t_L g1794 ( 
.A(n_1597),
.B(n_1336),
.Y(n_1794)
);

NAND2x1p5_ASAP7_75t_L g1795 ( 
.A(n_1597),
.B(n_1336),
.Y(n_1795)
);

AO22x2_ASAP7_75t_L g1796 ( 
.A1(n_1579),
.A2(n_802),
.B1(n_837),
.B2(n_745),
.Y(n_1796)
);

INVx2_ASAP7_75t_SL g1797 ( 
.A(n_1693),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1670),
.Y(n_1798)
);

INVxp67_ASAP7_75t_L g1799 ( 
.A(n_1562),
.Y(n_1799)
);

NAND2x1p5_ASAP7_75t_L g1800 ( 
.A(n_1597),
.B(n_1342),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1639),
.B(n_1342),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1549),
.Y(n_1802)
);

AOI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1592),
.A2(n_837),
.B1(n_852),
.B2(n_802),
.Y(n_1803)
);

AO22x2_ASAP7_75t_L g1804 ( 
.A1(n_1692),
.A2(n_1525),
.B1(n_1517),
.B2(n_1530),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1681),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_1558),
.Y(n_1806)
);

AOI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1615),
.A2(n_861),
.B1(n_873),
.B2(n_852),
.Y(n_1807)
);

AO22x2_ASAP7_75t_L g1808 ( 
.A1(n_1497),
.A2(n_861),
.B1(n_873),
.B2(n_852),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1507),
.B(n_861),
.Y(n_1809)
);

INVxp67_ASAP7_75t_L g1810 ( 
.A(n_1569),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1496),
.B(n_539),
.Y(n_1811)
);

OAI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1661),
.A2(n_873),
.B1(n_3),
.B2(n_1),
.C(n_2),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1687),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1687),
.Y(n_1814)
);

NOR2xp67_ASAP7_75t_L g1815 ( 
.A(n_1682),
.B(n_542),
.Y(n_1815)
);

AO22x2_ASAP7_75t_L g1816 ( 
.A1(n_1503),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1526),
.B(n_4),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1521),
.B(n_5),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1688),
.Y(n_1819)
);

AO22x2_ASAP7_75t_L g1820 ( 
.A1(n_1536),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1820)
);

NAND2x1p5_ASAP7_75t_L g1821 ( 
.A(n_1598),
.B(n_550),
.Y(n_1821)
);

AND2x4_ASAP7_75t_L g1822 ( 
.A(n_1488),
.B(n_544),
.Y(n_1822)
);

INVx3_ASAP7_75t_L g1823 ( 
.A(n_1541),
.Y(n_1823)
);

OAI221xp5_ASAP7_75t_L g1824 ( 
.A1(n_1663),
.A2(n_10),
.B1(n_7),
.B2(n_9),
.C(n_11),
.Y(n_1824)
);

OAI221xp5_ASAP7_75t_L g1825 ( 
.A1(n_1585),
.A2(n_12),
.B1(n_9),
.B2(n_10),
.C(n_13),
.Y(n_1825)
);

NOR2xp67_ASAP7_75t_L g1826 ( 
.A(n_1630),
.B(n_545),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1559),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1688),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1664),
.B(n_942),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1598),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1678),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1678),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1691),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1545),
.B(n_14),
.Y(n_1834)
);

AND2x2_ASAP7_75t_SL g1835 ( 
.A(n_1618),
.B(n_14),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1657),
.B(n_16),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1659),
.B(n_17),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_SL g1838 ( 
.A(n_1522),
.B(n_942),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1599),
.Y(n_1839)
);

AO22x1_ASAP7_75t_L g1840 ( 
.A1(n_1619),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1691),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1551),
.Y(n_1842)
);

AO22x2_ASAP7_75t_L g1843 ( 
.A1(n_1538),
.A2(n_22),
.B1(n_18),
.B2(n_21),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1598),
.Y(n_1844)
);

OR2x6_ASAP7_75t_L g1845 ( 
.A(n_1491),
.B(n_546),
.Y(n_1845)
);

AO22x2_ASAP7_75t_L g1846 ( 
.A1(n_1551),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_1846)
);

AO22x2_ASAP7_75t_L g1847 ( 
.A1(n_1572),
.A2(n_1529),
.B1(n_1535),
.B2(n_1668),
.Y(n_1847)
);

NAND2x1p5_ASAP7_75t_L g1848 ( 
.A(n_1669),
.B(n_556),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1669),
.Y(n_1849)
);

AO22x2_ASAP7_75t_L g1850 ( 
.A1(n_1572),
.A2(n_1494),
.B1(n_1534),
.B2(n_1531),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1680),
.B(n_942),
.Y(n_1851)
);

AOI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1656),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_1852)
);

BUFx6f_ASAP7_75t_SL g1853 ( 
.A(n_1669),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1685),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1660),
.Y(n_1855)
);

BUFx2_ASAP7_75t_L g1856 ( 
.A(n_1672),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1606),
.Y(n_1857)
);

BUFx8_ASAP7_75t_L g1858 ( 
.A(n_1541),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1489),
.B(n_25),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1671),
.Y(n_1860)
);

AO22x2_ASAP7_75t_L g1861 ( 
.A1(n_1490),
.A2(n_1495),
.B1(n_1677),
.B2(n_1679),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1684),
.B(n_26),
.Y(n_1862)
);

AO22x2_ASAP7_75t_L g1863 ( 
.A1(n_1490),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_1863)
);

OAI221xp5_ASAP7_75t_L g1864 ( 
.A1(n_1501),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.C(n_31),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1643),
.B(n_1658),
.Y(n_1865)
);

AO22x2_ASAP7_75t_L g1866 ( 
.A1(n_1495),
.A2(n_33),
.B1(n_30),
.B2(n_32),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1672),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1553),
.B(n_1565),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1672),
.Y(n_1869)
);

NAND2x1p5_ASAP7_75t_L g1870 ( 
.A(n_1554),
.B(n_557),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_1583),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1596),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1601),
.Y(n_1873)
);

NAND2x1p5_ASAP7_75t_L g1874 ( 
.A(n_1651),
.B(n_558),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1675),
.Y(n_1875)
);

INVxp67_ASAP7_75t_L g1876 ( 
.A(n_1654),
.Y(n_1876)
);

OAI221xp5_ASAP7_75t_L g1877 ( 
.A1(n_1624),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.C(n_35),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1677),
.B(n_34),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1603),
.Y(n_1879)
);

AO22x2_ASAP7_75t_L g1880 ( 
.A1(n_1673),
.A2(n_38),
.B1(n_35),
.B2(n_36),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1539),
.B(n_39),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1604),
.Y(n_1882)
);

NAND2x1p5_ASAP7_75t_L g1883 ( 
.A(n_1644),
.B(n_549),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1570),
.B(n_39),
.Y(n_1884)
);

AO22x2_ASAP7_75t_L g1885 ( 
.A1(n_1556),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1885)
);

OAI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1868),
.A2(n_1666),
.B(n_1557),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1830),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1818),
.A2(n_1676),
.B1(n_1552),
.B2(n_1623),
.Y(n_1888)
);

NOR3xp33_ASAP7_75t_L g1889 ( 
.A(n_1711),
.B(n_1812),
.C(n_1697),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1855),
.B(n_1519),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1764),
.B(n_1610),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1776),
.Y(n_1892)
);

INVxp67_ASAP7_75t_L g1893 ( 
.A(n_1701),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1860),
.B(n_1617),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1694),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1801),
.B(n_1620),
.Y(n_1896)
);

BUFx6f_ASAP7_75t_L g1897 ( 
.A(n_1830),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1700),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1799),
.A2(n_1631),
.B1(n_1636),
.B2(n_1622),
.Y(n_1899)
);

OAI321xp33_ASAP7_75t_L g1900 ( 
.A1(n_1824),
.A2(n_1640),
.A3(n_1637),
.B1(n_1645),
.B2(n_1609),
.C(n_1576),
.Y(n_1900)
);

NOR2x1_ASAP7_75t_L g1901 ( 
.A(n_1826),
.B(n_1575),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1809),
.B(n_1605),
.Y(n_1902)
);

O2A1O1Ixp33_ASAP7_75t_L g1903 ( 
.A1(n_1862),
.A2(n_1614),
.B(n_1621),
.C(n_1491),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1704),
.Y(n_1904)
);

OAI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1810),
.A2(n_1876),
.B1(n_1716),
.B2(n_1749),
.Y(n_1905)
);

OAI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1859),
.A2(n_1667),
.B(n_1595),
.Y(n_1906)
);

O2A1O1Ixp33_ASAP7_75t_L g1907 ( 
.A1(n_1877),
.A2(n_44),
.B(n_41),
.C(n_43),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1719),
.B(n_43),
.Y(n_1908)
);

OAI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1720),
.A2(n_1667),
.B1(n_1595),
.B2(n_46),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1695),
.Y(n_1910)
);

A2O1A1Ixp33_ASAP7_75t_L g1911 ( 
.A1(n_1834),
.A2(n_1836),
.B(n_1837),
.C(n_1817),
.Y(n_1911)
);

OAI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1779),
.A2(n_1667),
.B(n_1595),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1744),
.A2(n_1667),
.B1(n_1595),
.B2(n_46),
.Y(n_1913)
);

AOI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1805),
.A2(n_1667),
.B(n_639),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1813),
.B(n_44),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1814),
.A2(n_640),
.B(n_548),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1707),
.B(n_45),
.Y(n_1917)
);

NAND3xp33_ASAP7_75t_L g1918 ( 
.A(n_1852),
.B(n_47),
.C(n_48),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1819),
.B(n_48),
.Y(n_1919)
);

OAI21x1_ASAP7_75t_L g1920 ( 
.A1(n_1791),
.A2(n_553),
.B(n_547),
.Y(n_1920)
);

A2O1A1Ixp33_ASAP7_75t_L g1921 ( 
.A1(n_1872),
.A2(n_51),
.B(n_49),
.C(n_50),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1705),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1721),
.B(n_1873),
.Y(n_1923)
);

INVx5_ASAP7_75t_L g1924 ( 
.A(n_1733),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1698),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1851),
.B(n_1879),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1828),
.B(n_1831),
.Y(n_1927)
);

BUFx2_ASAP7_75t_L g1928 ( 
.A(n_1708),
.Y(n_1928)
);

BUFx3_ASAP7_75t_L g1929 ( 
.A(n_1724),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1832),
.A2(n_629),
.B(n_628),
.Y(n_1930)
);

A2O1A1Ixp33_ASAP7_75t_L g1931 ( 
.A1(n_1882),
.A2(n_52),
.B(n_49),
.C(n_50),
.Y(n_1931)
);

NOR3xp33_ASAP7_75t_L g1932 ( 
.A(n_1838),
.B(n_52),
.C(n_53),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1833),
.B(n_53),
.Y(n_1933)
);

INVx3_ASAP7_75t_L g1934 ( 
.A(n_1794),
.Y(n_1934)
);

BUFx3_ASAP7_75t_L g1935 ( 
.A(n_1708),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1709),
.Y(n_1936)
);

BUFx8_ASAP7_75t_L g1937 ( 
.A(n_1853),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1841),
.A2(n_637),
.B(n_636),
.Y(n_1938)
);

AOI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1842),
.A2(n_638),
.B(n_564),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1878),
.B(n_54),
.Y(n_1940)
);

O2A1O1Ixp33_ASAP7_75t_L g1941 ( 
.A1(n_1864),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_1941)
);

A2O1A1Ixp33_ASAP7_75t_L g1942 ( 
.A1(n_1803),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1727),
.B(n_60),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1742),
.B(n_560),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1727),
.B(n_60),
.Y(n_1945)
);

AOI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1774),
.A2(n_625),
.B(n_624),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1712),
.B(n_62),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1839),
.B(n_62),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1767),
.A2(n_632),
.B(n_630),
.Y(n_1949)
);

AOI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1710),
.A2(n_635),
.B(n_633),
.Y(n_1950)
);

HB1xp67_ASAP7_75t_L g1951 ( 
.A(n_1797),
.Y(n_1951)
);

OAI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1783),
.A2(n_63),
.B(n_65),
.Y(n_1952)
);

AOI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1710),
.A2(n_566),
.B(n_565),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1768),
.B(n_567),
.Y(n_1954)
);

AOI21xp5_ASAP7_75t_L g1955 ( 
.A1(n_1739),
.A2(n_608),
.B(n_607),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1696),
.B(n_568),
.Y(n_1956)
);

AO22x1_ASAP7_75t_L g1957 ( 
.A1(n_1871),
.A2(n_66),
.B1(n_63),
.B2(n_65),
.Y(n_1957)
);

INVx2_ASAP7_75t_SL g1958 ( 
.A(n_1802),
.Y(n_1958)
);

NOR3xp33_ASAP7_75t_L g1959 ( 
.A(n_1825),
.B(n_66),
.C(n_67),
.Y(n_1959)
);

O2A1O1Ixp33_ASAP7_75t_SL g1960 ( 
.A1(n_1884),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1763),
.B(n_69),
.Y(n_1961)
);

BUFx8_ASAP7_75t_SL g1962 ( 
.A(n_1778),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1881),
.B(n_1781),
.Y(n_1963)
);

INVxp67_ASAP7_75t_L g1964 ( 
.A(n_1728),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1781),
.B(n_70),
.Y(n_1965)
);

AOI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1758),
.A2(n_623),
.B(n_622),
.Y(n_1966)
);

INVxp67_ASAP7_75t_L g1967 ( 
.A(n_1747),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1807),
.A2(n_75),
.B1(n_72),
.B2(n_74),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1771),
.B(n_72),
.Y(n_1969)
);

AOI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1850),
.A2(n_601),
.B(n_600),
.Y(n_1970)
);

INVx3_ASAP7_75t_L g1971 ( 
.A(n_1795),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1850),
.A2(n_603),
.B(n_602),
.Y(n_1972)
);

AOI21xp33_ASAP7_75t_L g1973 ( 
.A1(n_1804),
.A2(n_1847),
.B(n_1787),
.Y(n_1973)
);

AO32x1_ASAP7_75t_L g1974 ( 
.A1(n_1857),
.A2(n_77),
.A3(n_74),
.B1(n_76),
.B2(n_78),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1702),
.B(n_77),
.Y(n_1975)
);

OAI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1761),
.A2(n_1788),
.B1(n_1789),
.B2(n_1755),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1723),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1771),
.B(n_78),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1804),
.B(n_79),
.Y(n_1979)
);

AOI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1773),
.A2(n_614),
.B(n_611),
.Y(n_1980)
);

OAI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1769),
.A2(n_79),
.B(n_80),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1725),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_SL g1983 ( 
.A(n_1865),
.B(n_80),
.Y(n_1983)
);

AOI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1773),
.A2(n_621),
.B(n_620),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1815),
.B(n_81),
.Y(n_1985)
);

OAI21xp5_ASAP7_75t_L g1986 ( 
.A1(n_1765),
.A2(n_81),
.B(n_83),
.Y(n_1986)
);

OAI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1702),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1987)
);

BUFx3_ASAP7_75t_L g1988 ( 
.A(n_1699),
.Y(n_1988)
);

AOI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1875),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1989)
);

CKINVDCx20_ASAP7_75t_R g1990 ( 
.A(n_1741),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1835),
.B(n_87),
.Y(n_1991)
);

AOI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1713),
.A2(n_1861),
.B(n_1847),
.Y(n_1992)
);

A2O1A1Ixp33_ASAP7_75t_L g1993 ( 
.A1(n_1811),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1717),
.B(n_88),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1822),
.B(n_90),
.Y(n_1995)
);

INVx3_ASAP7_75t_L g1996 ( 
.A(n_1786),
.Y(n_1996)
);

AOI21xp5_ASAP7_75t_L g1997 ( 
.A1(n_1713),
.A2(n_570),
.B(n_569),
.Y(n_1997)
);

OAI21x1_ASAP7_75t_L g1998 ( 
.A1(n_1800),
.A2(n_1870),
.B(n_1735),
.Y(n_1998)
);

AOI21x1_ASAP7_75t_L g1999 ( 
.A1(n_1861),
.A2(n_572),
.B(n_571),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_SL g2000 ( 
.A(n_1845),
.B(n_91),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1726),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1718),
.B(n_91),
.Y(n_2002)
);

AOI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1715),
.A2(n_627),
.B(n_575),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1715),
.A2(n_1874),
.B(n_1845),
.Y(n_2004)
);

O2A1O1Ixp33_ASAP7_75t_L g2005 ( 
.A1(n_1829),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1790),
.A2(n_576),
.B(n_574),
.Y(n_2006)
);

AOI21xp5_ASAP7_75t_L g2007 ( 
.A1(n_1883),
.A2(n_1731),
.B(n_1736),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1762),
.Y(n_2008)
);

AOI21xp5_ASAP7_75t_L g2009 ( 
.A1(n_1731),
.A2(n_578),
.B(n_577),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1722),
.B(n_92),
.Y(n_2010)
);

INVx4_ASAP7_75t_L g2011 ( 
.A(n_1806),
.Y(n_2011)
);

AOI21x1_ASAP7_75t_L g2012 ( 
.A1(n_1780),
.A2(n_580),
.B(n_579),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1703),
.B(n_93),
.Y(n_2013)
);

BUFx4f_ASAP7_75t_L g2014 ( 
.A(n_1750),
.Y(n_2014)
);

AOI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_1775),
.A2(n_583),
.B(n_582),
.Y(n_2015)
);

NAND3xp33_ASAP7_75t_L g2016 ( 
.A(n_1840),
.B(n_95),
.C(n_96),
.Y(n_2016)
);

BUFx2_ASAP7_75t_L g2017 ( 
.A(n_1856),
.Y(n_2017)
);

AOI21xp5_ASAP7_75t_L g2018 ( 
.A1(n_1777),
.A2(n_619),
.B(n_585),
.Y(n_2018)
);

AOI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_1854),
.A2(n_615),
.B(n_586),
.Y(n_2019)
);

CKINVDCx20_ASAP7_75t_R g2020 ( 
.A(n_1858),
.Y(n_2020)
);

NOR2x1_ASAP7_75t_L g2021 ( 
.A(n_1823),
.B(n_1759),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1703),
.B(n_96),
.Y(n_2022)
);

AOI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1737),
.A2(n_587),
.B(n_584),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1772),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1756),
.B(n_1757),
.Y(n_2025)
);

AOI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_1756),
.A2(n_1706),
.B1(n_1753),
.B2(n_1808),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1732),
.B(n_97),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1734),
.B(n_1751),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1760),
.Y(n_2029)
);

AND2x4_ASAP7_75t_L g2030 ( 
.A(n_1844),
.B(n_588),
.Y(n_2030)
);

AOI21xp5_ASAP7_75t_L g2031 ( 
.A1(n_1738),
.A2(n_591),
.B(n_589),
.Y(n_2031)
);

OAI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1752),
.A2(n_98),
.B(n_99),
.Y(n_2032)
);

AOI21xp5_ASAP7_75t_L g2033 ( 
.A1(n_1740),
.A2(n_593),
.B(n_592),
.Y(n_2033)
);

NAND2xp33_ASAP7_75t_L g2034 ( 
.A(n_1733),
.B(n_98),
.Y(n_2034)
);

INVxp67_ASAP7_75t_L g2035 ( 
.A(n_1784),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1754),
.B(n_99),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1743),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1757),
.B(n_100),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1766),
.B(n_100),
.Y(n_2039)
);

OAI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_1782),
.A2(n_597),
.B(n_596),
.Y(n_2040)
);

HB1xp67_ASAP7_75t_L g2041 ( 
.A(n_1849),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1745),
.Y(n_2042)
);

AOI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_1748),
.A2(n_610),
.B(n_599),
.Y(n_2043)
);

AOI21xp5_ASAP7_75t_L g2044 ( 
.A1(n_1821),
.A2(n_609),
.B(n_604),
.Y(n_2044)
);

AOI21xp5_ASAP7_75t_L g2045 ( 
.A1(n_1848),
.A2(n_605),
.B(n_598),
.Y(n_2045)
);

AOI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_1792),
.A2(n_536),
.B(n_101),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1766),
.B(n_101),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1785),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_1746),
.B(n_102),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1753),
.B(n_1798),
.Y(n_2050)
);

O2A1O1Ixp33_ASAP7_75t_L g2051 ( 
.A1(n_1827),
.A2(n_104),
.B(n_102),
.C(n_103),
.Y(n_2051)
);

AOI21xp5_ASAP7_75t_L g2052 ( 
.A1(n_1780),
.A2(n_536),
.B(n_103),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1706),
.B(n_104),
.Y(n_2053)
);

BUFx12f_ASAP7_75t_L g2054 ( 
.A(n_1730),
.Y(n_2054)
);

BUFx2_ASAP7_75t_L g2055 ( 
.A(n_1867),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1886),
.A2(n_1846),
.B(n_1816),
.Y(n_2056)
);

AOI21xp5_ASAP7_75t_L g2057 ( 
.A1(n_1946),
.A2(n_1846),
.B(n_1816),
.Y(n_2057)
);

AOI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_2034),
.A2(n_1866),
.B(n_1863),
.Y(n_2058)
);

AOI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_1906),
.A2(n_1866),
.B(n_1863),
.Y(n_2059)
);

O2A1O1Ixp33_ASAP7_75t_L g2060 ( 
.A1(n_1911),
.A2(n_1942),
.B(n_1907),
.C(n_1889),
.Y(n_2060)
);

BUFx5_ASAP7_75t_L g2061 ( 
.A(n_2029),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_R g2062 ( 
.A(n_1937),
.B(n_1869),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1895),
.Y(n_2063)
);

BUFx6f_ASAP7_75t_L g2064 ( 
.A(n_1929),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1926),
.B(n_1729),
.Y(n_2065)
);

NOR2xp33_ASAP7_75t_L g2066 ( 
.A(n_1967),
.B(n_1793),
.Y(n_2066)
);

CKINVDCx20_ASAP7_75t_R g2067 ( 
.A(n_1962),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1892),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1910),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1898),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_1902),
.B(n_1793),
.Y(n_2071)
);

BUFx2_ASAP7_75t_L g2072 ( 
.A(n_1935),
.Y(n_2072)
);

A2O1A1Ixp33_ASAP7_75t_SL g2073 ( 
.A1(n_1959),
.A2(n_1885),
.B(n_1808),
.C(n_1796),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1927),
.B(n_1880),
.Y(n_2074)
);

O2A1O1Ixp33_ASAP7_75t_SL g2075 ( 
.A1(n_1993),
.A2(n_1880),
.B(n_1885),
.C(n_1820),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1904),
.Y(n_2076)
);

INVx2_ASAP7_75t_SL g2077 ( 
.A(n_2014),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_L g2078 ( 
.A(n_1964),
.B(n_1714),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_SL g2079 ( 
.A(n_1888),
.B(n_1796),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1925),
.Y(n_2080)
);

BUFx2_ASAP7_75t_L g2081 ( 
.A(n_1928),
.Y(n_2081)
);

BUFx2_ASAP7_75t_L g2082 ( 
.A(n_2017),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_1903),
.B(n_1770),
.Y(n_2083)
);

NAND3xp33_ASAP7_75t_SL g2084 ( 
.A(n_2000),
.B(n_1843),
.C(n_1820),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_SL g2085 ( 
.A1(n_2026),
.A2(n_1843),
.B1(n_1770),
.B2(n_1733),
.Y(n_2085)
);

BUFx3_ASAP7_75t_L g2086 ( 
.A(n_1937),
.Y(n_2086)
);

HB1xp67_ASAP7_75t_L g2087 ( 
.A(n_1893),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1922),
.Y(n_2088)
);

BUFx3_ASAP7_75t_L g2089 ( 
.A(n_2014),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_R g2090 ( 
.A(n_1990),
.B(n_1770),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_SL g2091 ( 
.A(n_1894),
.B(n_105),
.Y(n_2091)
);

AOI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_1966),
.A2(n_2040),
.B(n_1981),
.Y(n_2092)
);

O2A1O1Ixp33_ASAP7_75t_L g2093 ( 
.A1(n_1941),
.A2(n_107),
.B(n_105),
.C(n_106),
.Y(n_2093)
);

INVx3_ASAP7_75t_L g2094 ( 
.A(n_1924),
.Y(n_2094)
);

CKINVDCx14_ASAP7_75t_R g2095 ( 
.A(n_2020),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1905),
.B(n_1890),
.Y(n_2096)
);

BUFx6f_ASAP7_75t_L g2097 ( 
.A(n_1887),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1891),
.B(n_1923),
.Y(n_2098)
);

AOI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_2040),
.A2(n_1900),
.B(n_1896),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1940),
.B(n_535),
.Y(n_2100)
);

BUFx6f_ASAP7_75t_L g2101 ( 
.A(n_1887),
.Y(n_2101)
);

BUFx2_ASAP7_75t_L g2102 ( 
.A(n_2055),
.Y(n_2102)
);

OAI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_1918),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_1996),
.B(n_108),
.Y(n_2104)
);

INVxp67_ASAP7_75t_SL g2105 ( 
.A(n_2035),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_1917),
.B(n_1908),
.Y(n_2106)
);

AOI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_1900),
.A2(n_109),
.B(n_111),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1963),
.B(n_111),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1936),
.Y(n_2109)
);

OAI22xp5_ASAP7_75t_L g2110 ( 
.A1(n_1918),
.A2(n_1991),
.B1(n_2016),
.B2(n_1989),
.Y(n_2110)
);

AOI21xp5_ASAP7_75t_L g2111 ( 
.A1(n_1912),
.A2(n_112),
.B(n_113),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1915),
.B(n_113),
.Y(n_2112)
);

BUFx2_ASAP7_75t_L g2113 ( 
.A(n_1951),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1977),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1919),
.B(n_534),
.Y(n_2115)
);

A2O1A1Ixp33_ASAP7_75t_L g2116 ( 
.A1(n_1986),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_2116)
);

INVx5_ASAP7_75t_L g2117 ( 
.A(n_1924),
.Y(n_2117)
);

A2O1A1Ixp33_ASAP7_75t_SL g2118 ( 
.A1(n_2032),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_2118)
);

CKINVDCx5p33_ASAP7_75t_R g2119 ( 
.A(n_1958),
.Y(n_2119)
);

NOR2xp33_ASAP7_75t_L g2120 ( 
.A(n_2011),
.B(n_118),
.Y(n_2120)
);

NOR2xp67_ASAP7_75t_SL g2121 ( 
.A(n_2016),
.B(n_118),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1982),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1933),
.B(n_534),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2037),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2001),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_SL g2126 ( 
.A(n_2011),
.B(n_119),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_SL g2127 ( 
.A(n_1901),
.B(n_120),
.Y(n_2127)
);

AOI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_1914),
.A2(n_120),
.B(n_121),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2028),
.B(n_532),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1899),
.B(n_532),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2025),
.B(n_122),
.Y(n_2131)
);

AOI21xp5_ASAP7_75t_L g2132 ( 
.A1(n_1909),
.A2(n_122),
.B(n_123),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_1975),
.B(n_124),
.Y(n_2133)
);

OAI22xp5_ASAP7_75t_L g2134 ( 
.A1(n_1995),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_L g2135 ( 
.A(n_1983),
.B(n_126),
.Y(n_2135)
);

INVx5_ASAP7_75t_L g2136 ( 
.A(n_1924),
.Y(n_2136)
);

OAI22xp5_ASAP7_75t_SL g2137 ( 
.A1(n_2053),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_2137)
);

OAI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_2021),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_2138)
);

NAND3xp33_ASAP7_75t_L g2139 ( 
.A(n_1932),
.B(n_1968),
.C(n_1952),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2042),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1943),
.B(n_130),
.Y(n_2141)
);

OR2x6_ASAP7_75t_SL g2142 ( 
.A(n_1987),
.B(n_130),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_SL g2143 ( 
.A(n_2000),
.B(n_131),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2008),
.Y(n_2144)
);

NOR3xp33_ASAP7_75t_SL g2145 ( 
.A(n_2052),
.B(n_1979),
.C(n_1945),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2024),
.Y(n_2146)
);

INVx3_ASAP7_75t_L g2147 ( 
.A(n_1934),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_SL g2148 ( 
.A(n_1985),
.B(n_131),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2048),
.Y(n_2149)
);

OAI22xp5_ASAP7_75t_SL g2150 ( 
.A1(n_2039),
.A2(n_135),
.B1(n_132),
.B2(n_134),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1965),
.Y(n_2151)
);

HB1xp67_ASAP7_75t_L g2152 ( 
.A(n_2041),
.Y(n_2152)
);

BUFx2_ASAP7_75t_SL g2153 ( 
.A(n_1988),
.Y(n_2153)
);

O2A1O1Ixp33_ASAP7_75t_L g2154 ( 
.A1(n_1921),
.A2(n_135),
.B(n_132),
.C(n_134),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1948),
.B(n_531),
.Y(n_2155)
);

O2A1O1Ixp33_ASAP7_75t_L g2156 ( 
.A1(n_1931),
.A2(n_139),
.B(n_137),
.C(n_138),
.Y(n_2156)
);

OAI22xp5_ASAP7_75t_L g2157 ( 
.A1(n_2050),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2038),
.B(n_140),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2013),
.B(n_140),
.Y(n_2159)
);

OAI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_1947),
.A2(n_144),
.B1(n_141),
.B2(n_142),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2022),
.B(n_531),
.Y(n_2161)
);

BUFx2_ASAP7_75t_L g2162 ( 
.A(n_1887),
.Y(n_2162)
);

INVxp67_ASAP7_75t_SL g2163 ( 
.A(n_1998),
.Y(n_2163)
);

NOR3xp33_ASAP7_75t_L g2164 ( 
.A(n_1957),
.B(n_2005),
.C(n_2047),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_2054),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2061),
.Y(n_2166)
);

INVx2_ASAP7_75t_SL g2167 ( 
.A(n_2064),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2124),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2140),
.Y(n_2169)
);

AND2x4_ASAP7_75t_L g2170 ( 
.A(n_2081),
.B(n_2004),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2061),
.Y(n_2171)
);

AOI21xp33_ASAP7_75t_L g2172 ( 
.A1(n_2060),
.A2(n_1973),
.B(n_1913),
.Y(n_2172)
);

OAI22x1_ASAP7_75t_L g2173 ( 
.A1(n_2079),
.A2(n_1969),
.B1(n_1978),
.B2(n_2012),
.Y(n_2173)
);

BUFx2_ASAP7_75t_L g2174 ( 
.A(n_2102),
.Y(n_2174)
);

INVx3_ASAP7_75t_L g2175 ( 
.A(n_2147),
.Y(n_2175)
);

AOI22xp33_ASAP7_75t_L g2176 ( 
.A1(n_2139),
.A2(n_1976),
.B1(n_2049),
.B2(n_1954),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2063),
.Y(n_2177)
);

BUFx8_ASAP7_75t_L g2178 ( 
.A(n_2086),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2070),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_2067),
.Y(n_2180)
);

BUFx12f_ASAP7_75t_L g2181 ( 
.A(n_2165),
.Y(n_2181)
);

INVx1_ASAP7_75t_SL g2182 ( 
.A(n_2072),
.Y(n_2182)
);

AOI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_2139),
.A2(n_2007),
.B1(n_2046),
.B2(n_2009),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2076),
.Y(n_2184)
);

BUFx6f_ASAP7_75t_L g2185 ( 
.A(n_2064),
.Y(n_2185)
);

BUFx6f_ASAP7_75t_L g2186 ( 
.A(n_2064),
.Y(n_2186)
);

BUFx6f_ASAP7_75t_L g2187 ( 
.A(n_2097),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2088),
.Y(n_2188)
);

INVx5_ASAP7_75t_L g2189 ( 
.A(n_2117),
.Y(n_2189)
);

HB1xp67_ASAP7_75t_L g2190 ( 
.A(n_2152),
.Y(n_2190)
);

BUFx3_ASAP7_75t_L g2191 ( 
.A(n_2082),
.Y(n_2191)
);

AOI22xp5_ASAP7_75t_L g2192 ( 
.A1(n_2110),
.A2(n_1956),
.B1(n_1944),
.B2(n_1996),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_2097),
.Y(n_2193)
);

BUFx6f_ASAP7_75t_L g2194 ( 
.A(n_2097),
.Y(n_2194)
);

AOI21xp5_ASAP7_75t_L g2195 ( 
.A1(n_2092),
.A2(n_2099),
.B(n_2083),
.Y(n_2195)
);

AOI21xp5_ASAP7_75t_L g2196 ( 
.A1(n_2096),
.A2(n_1974),
.B(n_1955),
.Y(n_2196)
);

INVxp67_ASAP7_75t_SL g2197 ( 
.A(n_2105),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2106),
.B(n_1992),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2109),
.Y(n_2199)
);

INVx3_ASAP7_75t_SL g2200 ( 
.A(n_2119),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2114),
.Y(n_2201)
);

INVx1_ASAP7_75t_SL g2202 ( 
.A(n_2098),
.Y(n_2202)
);

INVx4_ASAP7_75t_L g2203 ( 
.A(n_2117),
.Y(n_2203)
);

OR2x6_ASAP7_75t_L g2204 ( 
.A(n_2058),
.B(n_2003),
.Y(n_2204)
);

AND2x6_ASAP7_75t_L g2205 ( 
.A(n_2094),
.B(n_2030),
.Y(n_2205)
);

BUFx6f_ASAP7_75t_L g2206 ( 
.A(n_2101),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2061),
.Y(n_2207)
);

BUFx4f_ASAP7_75t_L g2208 ( 
.A(n_2101),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2061),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_L g2210 ( 
.A(n_2071),
.B(n_2066),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2151),
.B(n_2036),
.Y(n_2211)
);

BUFx6f_ASAP7_75t_L g2212 ( 
.A(n_2101),
.Y(n_2212)
);

AOI22xp33_ASAP7_75t_L g2213 ( 
.A1(n_2164),
.A2(n_1961),
.B1(n_1956),
.B2(n_2030),
.Y(n_2213)
);

BUFx6f_ASAP7_75t_L g2214 ( 
.A(n_2089),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2133),
.B(n_1897),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2144),
.Y(n_2216)
);

INVx2_ASAP7_75t_SL g2217 ( 
.A(n_2113),
.Y(n_2217)
);

INVx2_ASAP7_75t_SL g2218 ( 
.A(n_2062),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2122),
.B(n_1897),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2061),
.Y(n_2220)
);

INVx3_ASAP7_75t_SL g2221 ( 
.A(n_2077),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2125),
.Y(n_2222)
);

BUFx12f_ASAP7_75t_L g2223 ( 
.A(n_2104),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2146),
.Y(n_2224)
);

CKINVDCx11_ASAP7_75t_R g2225 ( 
.A(n_2142),
.Y(n_2225)
);

INVx1_ASAP7_75t_SL g2226 ( 
.A(n_2153),
.Y(n_2226)
);

OR2x6_ASAP7_75t_L g2227 ( 
.A(n_2056),
.B(n_1950),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2074),
.B(n_1994),
.Y(n_2228)
);

OAI222xp33_ASAP7_75t_L g2229 ( 
.A1(n_2121),
.A2(n_2051),
.B1(n_1970),
.B2(n_1972),
.C1(n_1953),
.C2(n_1997),
.Y(n_2229)
);

OR2x2_ASAP7_75t_L g2230 ( 
.A(n_2149),
.B(n_2002),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2163),
.Y(n_2231)
);

OAI221xp5_ASAP7_75t_L g2232 ( 
.A1(n_2073),
.A2(n_1960),
.B1(n_1949),
.B2(n_2019),
.C(n_2018),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2197),
.B(n_2059),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2202),
.B(n_2087),
.Y(n_2234)
);

OR2x6_ASAP7_75t_L g2235 ( 
.A(n_2195),
.B(n_2204),
.Y(n_2235)
);

AOI21xp5_ASAP7_75t_L g2236 ( 
.A1(n_2196),
.A2(n_2116),
.B(n_2118),
.Y(n_2236)
);

A2O1A1Ixp33_ASAP7_75t_L g2237 ( 
.A1(n_2176),
.A2(n_2093),
.B(n_2156),
.C(n_2154),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2222),
.Y(n_2238)
);

BUFx6f_ASAP7_75t_L g2239 ( 
.A(n_2185),
.Y(n_2239)
);

OR2x6_ASAP7_75t_SL g2240 ( 
.A(n_2180),
.B(n_2131),
.Y(n_2240)
);

INVx5_ASAP7_75t_L g2241 ( 
.A(n_2204),
.Y(n_2241)
);

AOI21xp5_ASAP7_75t_L g2242 ( 
.A1(n_2232),
.A2(n_2057),
.B(n_2128),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2190),
.B(n_2108),
.Y(n_2243)
);

OR2x2_ASAP7_75t_L g2244 ( 
.A(n_2222),
.B(n_2141),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2168),
.Y(n_2245)
);

BUFx2_ASAP7_75t_L g2246 ( 
.A(n_2174),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2224),
.Y(n_2247)
);

OR2x2_ASAP7_75t_SL g2248 ( 
.A(n_2228),
.B(n_2084),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2169),
.B(n_2145),
.Y(n_2249)
);

OAI22xp5_ASAP7_75t_L g2250 ( 
.A1(n_2213),
.A2(n_2085),
.B1(n_2137),
.B2(n_2143),
.Y(n_2250)
);

AOI21xp5_ASAP7_75t_L g2251 ( 
.A1(n_2229),
.A2(n_2111),
.B(n_2075),
.Y(n_2251)
);

BUFx3_ASAP7_75t_L g2252 ( 
.A(n_2178),
.Y(n_2252)
);

AOI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_2192),
.A2(n_2103),
.B1(n_2126),
.B2(n_2150),
.Y(n_2253)
);

OAI22xp5_ASAP7_75t_L g2254 ( 
.A1(n_2183),
.A2(n_2085),
.B1(n_2137),
.B2(n_2150),
.Y(n_2254)
);

AOI22xp5_ASAP7_75t_L g2255 ( 
.A1(n_2210),
.A2(n_2130),
.B1(n_2135),
.B2(n_2157),
.Y(n_2255)
);

INVx4_ASAP7_75t_L g2256 ( 
.A(n_2185),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_2185),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2216),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2198),
.B(n_2120),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2224),
.Y(n_2260)
);

INVx1_ASAP7_75t_SL g2261 ( 
.A(n_2226),
.Y(n_2261)
);

NAND2x1p5_ASAP7_75t_L g2262 ( 
.A(n_2189),
.B(n_2117),
.Y(n_2262)
);

AOI22xp5_ASAP7_75t_L g2263 ( 
.A1(n_2227),
.A2(n_2160),
.B1(n_2134),
.B2(n_2127),
.Y(n_2263)
);

AOI21xp5_ASAP7_75t_L g2264 ( 
.A1(n_2172),
.A2(n_2136),
.B(n_1984),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2191),
.B(n_2162),
.Y(n_2265)
);

CKINVDCx5p33_ASAP7_75t_R g2266 ( 
.A(n_2200),
.Y(n_2266)
);

OAI22xp5_ASAP7_75t_L g2267 ( 
.A1(n_2227),
.A2(n_2107),
.B1(n_2132),
.B2(n_2138),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2177),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2179),
.Y(n_2269)
);

AND2x4_ASAP7_75t_L g2270 ( 
.A(n_2170),
.B(n_2136),
.Y(n_2270)
);

OR2x6_ASAP7_75t_L g2271 ( 
.A(n_2203),
.B(n_1980),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_2186),
.Y(n_2272)
);

AOI22xp33_ASAP7_75t_L g2273 ( 
.A1(n_2254),
.A2(n_2225),
.B1(n_2173),
.B2(n_2170),
.Y(n_2273)
);

BUFx8_ASAP7_75t_L g2274 ( 
.A(n_2252),
.Y(n_2274)
);

INVx2_ASAP7_75t_SL g2275 ( 
.A(n_2246),
.Y(n_2275)
);

BUFx8_ASAP7_75t_L g2276 ( 
.A(n_2239),
.Y(n_2276)
);

INVx6_ASAP7_75t_L g2277 ( 
.A(n_2241),
.Y(n_2277)
);

INVx2_ASAP7_75t_SL g2278 ( 
.A(n_2268),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2238),
.Y(n_2279)
);

CKINVDCx11_ASAP7_75t_R g2280 ( 
.A(n_2240),
.Y(n_2280)
);

NAND2x1p5_ASAP7_75t_L g2281 ( 
.A(n_2241),
.B(n_2189),
.Y(n_2281)
);

AOI22xp33_ASAP7_75t_L g2282 ( 
.A1(n_2267),
.A2(n_2223),
.B1(n_2205),
.B2(n_2148),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2247),
.Y(n_2283)
);

INVx3_ASAP7_75t_L g2284 ( 
.A(n_2270),
.Y(n_2284)
);

AOI22xp33_ASAP7_75t_L g2285 ( 
.A1(n_2251),
.A2(n_2205),
.B1(n_2091),
.B2(n_2158),
.Y(n_2285)
);

BUFx12f_ASAP7_75t_L g2286 ( 
.A(n_2266),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_2261),
.Y(n_2287)
);

AOI22xp33_ASAP7_75t_L g2288 ( 
.A1(n_2250),
.A2(n_2205),
.B1(n_2159),
.B2(n_2161),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_2239),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2260),
.Y(n_2290)
);

CKINVDCx20_ASAP7_75t_R g2291 ( 
.A(n_2265),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2269),
.Y(n_2292)
);

BUFx12f_ASAP7_75t_L g2293 ( 
.A(n_2248),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_2245),
.Y(n_2294)
);

CKINVDCx5p33_ASAP7_75t_R g2295 ( 
.A(n_2239),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2233),
.B(n_2217),
.Y(n_2296)
);

BUFx2_ASAP7_75t_SL g2297 ( 
.A(n_2241),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2258),
.Y(n_2298)
);

INVx2_ASAP7_75t_SL g2299 ( 
.A(n_2275),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2279),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2279),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2283),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2283),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2284),
.B(n_2235),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2290),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2278),
.Y(n_2306)
);

AOI22xp33_ASAP7_75t_L g2307 ( 
.A1(n_2293),
.A2(n_2242),
.B1(n_2236),
.B2(n_2235),
.Y(n_2307)
);

BUFx6f_ASAP7_75t_L g2308 ( 
.A(n_2286),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2302),
.Y(n_2309)
);

HB1xp67_ASAP7_75t_L g2310 ( 
.A(n_2306),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2302),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2306),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2300),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2301),
.Y(n_2314)
);

AO21x2_ASAP7_75t_L g2315 ( 
.A1(n_2304),
.A2(n_2264),
.B(n_1999),
.Y(n_2315)
);

OR2x2_ASAP7_75t_L g2316 ( 
.A(n_2313),
.B(n_2275),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2314),
.B(n_2303),
.Y(n_2317)
);

OAI211xp5_ASAP7_75t_L g2318 ( 
.A1(n_2310),
.A2(n_2280),
.B(n_2253),
.C(n_2288),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2312),
.B(n_2304),
.Y(n_2319)
);

AO21x2_ASAP7_75t_L g2320 ( 
.A1(n_2309),
.A2(n_2305),
.B(n_2293),
.Y(n_2320)
);

AO32x1_ASAP7_75t_L g2321 ( 
.A1(n_2312),
.A2(n_2299),
.A3(n_2256),
.B1(n_2203),
.B2(n_2167),
.Y(n_2321)
);

NOR2x1_ASAP7_75t_SL g2322 ( 
.A(n_2314),
.B(n_2297),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2311),
.B(n_2284),
.Y(n_2323)
);

OAI22xp5_ASAP7_75t_SL g2324 ( 
.A1(n_2309),
.A2(n_2307),
.B1(n_2308),
.B2(n_2273),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2315),
.B(n_2284),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2319),
.B(n_2299),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2322),
.B(n_2308),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2320),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2317),
.Y(n_2329)
);

INVxp67_ASAP7_75t_L g2330 ( 
.A(n_2320),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2321),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2318),
.B(n_2259),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2317),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_2323),
.B(n_2308),
.Y(n_2334)
);

INVx3_ASAP7_75t_L g2335 ( 
.A(n_2316),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2318),
.B(n_2308),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2329),
.B(n_2333),
.Y(n_2337)
);

OR2x2_ASAP7_75t_L g2338 ( 
.A(n_2335),
.B(n_2324),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2334),
.B(n_2308),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2334),
.Y(n_2340)
);

NOR3xp33_ASAP7_75t_L g2341 ( 
.A(n_2336),
.B(n_2100),
.C(n_2237),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2335),
.B(n_2325),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2326),
.B(n_2095),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2326),
.B(n_2286),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2335),
.B(n_2287),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2343),
.Y(n_2346)
);

HB1xp67_ASAP7_75t_L g2347 ( 
.A(n_2340),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2341),
.B(n_2332),
.Y(n_2348)
);

INVx2_ASAP7_75t_SL g2349 ( 
.A(n_2339),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2349),
.B(n_2344),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2346),
.B(n_2327),
.Y(n_2351)
);

HB1xp67_ASAP7_75t_L g2352 ( 
.A(n_2347),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2348),
.B(n_2338),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2352),
.Y(n_2354)
);

AND2x4_ASAP7_75t_L g2355 ( 
.A(n_2351),
.B(n_2345),
.Y(n_2355)
);

OR2x6_ASAP7_75t_L g2356 ( 
.A(n_2350),
.B(n_2181),
.Y(n_2356)
);

OR2x2_ASAP7_75t_L g2357 ( 
.A(n_2353),
.B(n_2342),
.Y(n_2357)
);

OR2x2_ASAP7_75t_L g2358 ( 
.A(n_2352),
.B(n_2337),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2352),
.Y(n_2359)
);

OR2x2_ASAP7_75t_L g2360 ( 
.A(n_2354),
.B(n_2359),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2358),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2357),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2355),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2356),
.B(n_2337),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2354),
.B(n_2330),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2355),
.B(n_2327),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2355),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2355),
.B(n_2328),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2355),
.B(n_2328),
.Y(n_2369)
);

INVxp67_ASAP7_75t_SL g2370 ( 
.A(n_2366),
.Y(n_2370)
);

INVx1_ASAP7_75t_SL g2371 ( 
.A(n_2360),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2363),
.B(n_2331),
.Y(n_2372)
);

INVx3_ASAP7_75t_L g2373 ( 
.A(n_2367),
.Y(n_2373)
);

XNOR2xp5_ASAP7_75t_L g2374 ( 
.A(n_2362),
.B(n_2218),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2361),
.B(n_2331),
.Y(n_2375)
);

XOR2x2_ASAP7_75t_L g2376 ( 
.A(n_2364),
.B(n_2178),
.Y(n_2376)
);

XOR2x2_ASAP7_75t_L g2377 ( 
.A(n_2364),
.B(n_2368),
.Y(n_2377)
);

INVx2_ASAP7_75t_SL g2378 ( 
.A(n_2369),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2365),
.Y(n_2379)
);

XOR2x2_ASAP7_75t_L g2380 ( 
.A(n_2365),
.B(n_2221),
.Y(n_2380)
);

NOR2xp33_ASAP7_75t_L g2381 ( 
.A(n_2363),
.B(n_2274),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2366),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2370),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2376),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2377),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2373),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2373),
.Y(n_2387)
);

NAND3x1_ASAP7_75t_L g2388 ( 
.A(n_2372),
.B(n_2274),
.C(n_2115),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2375),
.Y(n_2389)
);

OAI22xp5_ASAP7_75t_L g2390 ( 
.A1(n_2371),
.A2(n_2287),
.B1(n_2255),
.B2(n_2123),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2382),
.Y(n_2391)
);

AOI22xp33_ASAP7_75t_L g2392 ( 
.A1(n_2381),
.A2(n_2297),
.B1(n_2315),
.B2(n_2274),
.Y(n_2392)
);

HB1xp67_ASAP7_75t_L g2393 ( 
.A(n_2374),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2378),
.B(n_2234),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2380),
.B(n_2291),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2379),
.Y(n_2396)
);

OAI22xp5_ASAP7_75t_L g2397 ( 
.A1(n_2379),
.A2(n_2277),
.B1(n_2285),
.B2(n_2289),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2389),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2383),
.Y(n_2399)
);

OAI22xp5_ASAP7_75t_L g2400 ( 
.A1(n_2385),
.A2(n_2277),
.B1(n_2295),
.B2(n_2289),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2386),
.Y(n_2401)
);

NOR2xp33_ASAP7_75t_L g2402 ( 
.A(n_2387),
.B(n_2214),
.Y(n_2402)
);

INVxp67_ASAP7_75t_L g2403 ( 
.A(n_2393),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_SL g2404 ( 
.A(n_2390),
.B(n_2214),
.Y(n_2404)
);

HB1xp67_ASAP7_75t_L g2405 ( 
.A(n_2396),
.Y(n_2405)
);

OAI22xp5_ASAP7_75t_L g2406 ( 
.A1(n_2391),
.A2(n_2277),
.B1(n_2295),
.B2(n_2182),
.Y(n_2406)
);

INVx3_ASAP7_75t_L g2407 ( 
.A(n_2388),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2394),
.Y(n_2408)
);

INVxp67_ASAP7_75t_SL g2409 ( 
.A(n_2384),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2390),
.Y(n_2410)
);

INVx1_ASAP7_75t_SL g2411 ( 
.A(n_2395),
.Y(n_2411)
);

INVxp67_ASAP7_75t_SL g2412 ( 
.A(n_2405),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2409),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2398),
.Y(n_2414)
);

OAI222xp33_ASAP7_75t_L g2415 ( 
.A1(n_2400),
.A2(n_2392),
.B1(n_2397),
.B2(n_2112),
.C1(n_2155),
.C2(n_2321),
.Y(n_2415)
);

OR2x2_ASAP7_75t_L g2416 ( 
.A(n_2410),
.B(n_2243),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2402),
.B(n_2407),
.Y(n_2417)
);

AO21x1_ASAP7_75t_L g2418 ( 
.A1(n_2401),
.A2(n_2321),
.B(n_2129),
.Y(n_2418)
);

AOI21xp33_ASAP7_75t_L g2419 ( 
.A1(n_2403),
.A2(n_2027),
.B(n_2010),
.Y(n_2419)
);

AOI22xp5_ASAP7_75t_L g2420 ( 
.A1(n_2411),
.A2(n_2214),
.B1(n_2277),
.B2(n_2186),
.Y(n_2420)
);

OAI21xp5_ASAP7_75t_L g2421 ( 
.A1(n_2399),
.A2(n_2211),
.B(n_2104),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2407),
.B(n_2315),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2404),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2406),
.B(n_2215),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2408),
.B(n_2249),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_SL g2426 ( 
.A(n_2407),
.B(n_2186),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2409),
.B(n_2296),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2409),
.B(n_2244),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2405),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2407),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2405),
.Y(n_2431)
);

NAND4xp25_ASAP7_75t_L g2432 ( 
.A(n_2400),
.B(n_2282),
.C(n_2263),
.D(n_2078),
.Y(n_2432)
);

AOI22xp33_ASAP7_75t_L g2433 ( 
.A1(n_2409),
.A2(n_2276),
.B1(n_2256),
.B2(n_2272),
.Y(n_2433)
);

INVx3_ASAP7_75t_L g2434 ( 
.A(n_2430),
.Y(n_2434)
);

NOR2x1_ASAP7_75t_L g2435 ( 
.A(n_2429),
.B(n_142),
.Y(n_2435)
);

INVxp67_ASAP7_75t_L g2436 ( 
.A(n_2412),
.Y(n_2436)
);

NOR2xp33_ASAP7_75t_L g2437 ( 
.A(n_2431),
.B(n_145),
.Y(n_2437)
);

OR2x2_ASAP7_75t_L g2438 ( 
.A(n_2413),
.B(n_146),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2417),
.Y(n_2439)
);

OR2x2_ASAP7_75t_L g2440 ( 
.A(n_2426),
.B(n_147),
.Y(n_2440)
);

AOI22xp5_ASAP7_75t_L g2441 ( 
.A1(n_2414),
.A2(n_1897),
.B1(n_2281),
.B2(n_2278),
.Y(n_2441)
);

NOR2xp33_ASAP7_75t_L g2442 ( 
.A(n_2416),
.B(n_148),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2427),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2420),
.B(n_2423),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2428),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2433),
.B(n_149),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2424),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2421),
.B(n_150),
.Y(n_2448)
);

NOR2xp33_ASAP7_75t_L g2449 ( 
.A(n_2425),
.B(n_152),
.Y(n_2449)
);

HB1xp67_ASAP7_75t_L g2450 ( 
.A(n_2422),
.Y(n_2450)
);

AND2x2_ASAP7_75t_L g2451 ( 
.A(n_2419),
.B(n_2281),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2432),
.B(n_152),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2418),
.B(n_153),
.Y(n_2453)
);

OR2x2_ASAP7_75t_L g2454 ( 
.A(n_2415),
.B(n_154),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2413),
.B(n_2281),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2412),
.Y(n_2456)
);

NOR2xp33_ASAP7_75t_L g2457 ( 
.A(n_2430),
.B(n_155),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2412),
.B(n_156),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2412),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2412),
.B(n_156),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2412),
.B(n_157),
.Y(n_2461)
);

NAND2xp33_ASAP7_75t_L g2462 ( 
.A(n_2430),
.B(n_2090),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_2413),
.B(n_2292),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2413),
.B(n_2292),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2412),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2412),
.Y(n_2466)
);

NAND2x1p5_ASAP7_75t_L g2467 ( 
.A(n_2429),
.B(n_2136),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2412),
.B(n_158),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2412),
.B(n_159),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2413),
.B(n_2294),
.Y(n_2470)
);

OA22x2_ASAP7_75t_L g2471 ( 
.A1(n_2456),
.A2(n_2459),
.B1(n_2466),
.B2(n_2465),
.Y(n_2471)
);

AOI22xp5_ASAP7_75t_L g2472 ( 
.A1(n_2462),
.A2(n_2276),
.B1(n_2272),
.B2(n_2257),
.Y(n_2472)
);

AOI22xp5_ASAP7_75t_L g2473 ( 
.A1(n_2436),
.A2(n_2276),
.B1(n_2272),
.B2(n_2257),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2438),
.Y(n_2474)
);

AND4x1_ASAP7_75t_L g2475 ( 
.A(n_2435),
.B(n_161),
.C(n_159),
.D(n_160),
.Y(n_2475)
);

OAI22xp5_ASAP7_75t_L g2476 ( 
.A1(n_2434),
.A2(n_2271),
.B1(n_2257),
.B2(n_2208),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2458),
.Y(n_2477)
);

AOI22xp33_ASAP7_75t_L g2478 ( 
.A1(n_2434),
.A2(n_2276),
.B1(n_2271),
.B2(n_2193),
.Y(n_2478)
);

OAI22xp5_ASAP7_75t_L g2479 ( 
.A1(n_2439),
.A2(n_2208),
.B1(n_2262),
.B2(n_2230),
.Y(n_2479)
);

INVx2_ASAP7_75t_SL g2480 ( 
.A(n_2440),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2460),
.Y(n_2481)
);

BUFx6f_ASAP7_75t_L g2482 ( 
.A(n_2461),
.Y(n_2482)
);

AO221x1_ASAP7_75t_L g2483 ( 
.A1(n_2447),
.A2(n_2194),
.B1(n_2206),
.B2(n_2193),
.C(n_2187),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2468),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2469),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2455),
.Y(n_2486)
);

BUFx3_ASAP7_75t_L g2487 ( 
.A(n_2444),
.Y(n_2487)
);

AOI22xp5_ASAP7_75t_L g2488 ( 
.A1(n_2445),
.A2(n_2193),
.B1(n_2194),
.B2(n_2187),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2437),
.Y(n_2489)
);

HB1xp67_ASAP7_75t_SL g2490 ( 
.A(n_2443),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2454),
.Y(n_2491)
);

AOI221xp5_ASAP7_75t_L g2492 ( 
.A1(n_2442),
.A2(n_2446),
.B1(n_2453),
.B2(n_2452),
.C(n_2448),
.Y(n_2492)
);

OAI322xp33_ASAP7_75t_L g2493 ( 
.A1(n_2467),
.A2(n_2015),
.A3(n_2043),
.B1(n_2031),
.B2(n_2033),
.C1(n_2023),
.C2(n_1939),
.Y(n_2493)
);

AOI22xp5_ASAP7_75t_L g2494 ( 
.A1(n_2451),
.A2(n_2194),
.B1(n_2206),
.B2(n_2187),
.Y(n_2494)
);

INVxp67_ASAP7_75t_L g2495 ( 
.A(n_2457),
.Y(n_2495)
);

AOI22x1_ASAP7_75t_L g2496 ( 
.A1(n_2450),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_2496)
);

NAND4xp25_ASAP7_75t_SL g2497 ( 
.A(n_2470),
.B(n_2044),
.C(n_2045),
.D(n_2006),
.Y(n_2497)
);

AOI221xp5_ASAP7_75t_L g2498 ( 
.A1(n_2449),
.A2(n_1938),
.B1(n_1930),
.B2(n_1916),
.C(n_164),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2463),
.Y(n_2499)
);

AND4x1_ASAP7_75t_L g2500 ( 
.A(n_2464),
.B(n_164),
.C(n_162),
.D(n_163),
.Y(n_2500)
);

AOI31xp33_ASAP7_75t_L g2501 ( 
.A1(n_2441),
.A2(n_166),
.A3(n_163),
.B(n_165),
.Y(n_2501)
);

AO22x2_ASAP7_75t_L g2502 ( 
.A1(n_2441),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2438),
.Y(n_2503)
);

OAI22x1_ASAP7_75t_SL g2504 ( 
.A1(n_2456),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_2504)
);

AND4x1_ASAP7_75t_L g2505 ( 
.A(n_2435),
.B(n_170),
.C(n_168),
.D(n_169),
.Y(n_2505)
);

AOI22x1_ASAP7_75t_L g2506 ( 
.A1(n_2456),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_2506)
);

OAI22xp5_ASAP7_75t_L g2507 ( 
.A1(n_2436),
.A2(n_2290),
.B1(n_2189),
.B2(n_2212),
.Y(n_2507)
);

OAI322xp33_ASAP7_75t_L g2508 ( 
.A1(n_2436),
.A2(n_176),
.A3(n_175),
.B1(n_173),
.B2(n_171),
.C1(n_172),
.C2(n_174),
.Y(n_2508)
);

NOR3xp33_ASAP7_75t_L g2509 ( 
.A(n_2486),
.B(n_2491),
.C(n_2492),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_2500),
.B(n_2475),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2505),
.Y(n_2511)
);

AOI22xp5_ASAP7_75t_L g2512 ( 
.A1(n_2473),
.A2(n_2212),
.B1(n_2206),
.B2(n_2270),
.Y(n_2512)
);

OAI22xp5_ASAP7_75t_L g2513 ( 
.A1(n_2478),
.A2(n_2212),
.B1(n_2298),
.B2(n_2294),
.Y(n_2513)
);

NOR3xp33_ASAP7_75t_L g2514 ( 
.A(n_2503),
.B(n_173),
.C(n_174),
.Y(n_2514)
);

AOI31xp33_ASAP7_75t_L g2515 ( 
.A1(n_2499),
.A2(n_177),
.A3(n_175),
.B(n_176),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2487),
.B(n_2298),
.Y(n_2516)
);

OA211x2_ASAP7_75t_L g2517 ( 
.A1(n_2495),
.A2(n_179),
.B(n_177),
.C(n_178),
.Y(n_2517)
);

OAI21xp33_ASAP7_75t_L g2518 ( 
.A1(n_2471),
.A2(n_2219),
.B(n_2065),
.Y(n_2518)
);

AOI21xp5_ASAP7_75t_L g2519 ( 
.A1(n_2474),
.A2(n_178),
.B(n_179),
.Y(n_2519)
);

NAND4xp25_ASAP7_75t_L g2520 ( 
.A(n_2489),
.B(n_2477),
.C(n_2484),
.D(n_2481),
.Y(n_2520)
);

AOI21xp5_ASAP7_75t_L g2521 ( 
.A1(n_2501),
.A2(n_2480),
.B(n_2485),
.Y(n_2521)
);

NOR3x1_ASAP7_75t_L g2522 ( 
.A(n_2483),
.B(n_180),
.C(n_181),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2506),
.B(n_180),
.Y(n_2523)
);

OAI21x1_ASAP7_75t_L g2524 ( 
.A1(n_2496),
.A2(n_1920),
.B(n_2094),
.Y(n_2524)
);

AOI211x1_ASAP7_75t_SL g2525 ( 
.A1(n_2507),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_2525)
);

NOR3xp33_ASAP7_75t_L g2526 ( 
.A(n_2508),
.B(n_184),
.C(n_185),
.Y(n_2526)
);

AOI21xp5_ASAP7_75t_L g2527 ( 
.A1(n_2502),
.A2(n_186),
.B(n_187),
.Y(n_2527)
);

AOI21xp5_ASAP7_75t_L g2528 ( 
.A1(n_2502),
.A2(n_186),
.B(n_187),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2504),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_SL g2530 ( 
.A(n_2482),
.B(n_188),
.Y(n_2530)
);

NAND3xp33_ASAP7_75t_SL g2531 ( 
.A(n_2490),
.B(n_188),
.C(n_189),
.Y(n_2531)
);

OAI211xp5_ASAP7_75t_L g2532 ( 
.A1(n_2482),
.A2(n_191),
.B(n_189),
.C(n_190),
.Y(n_2532)
);

AOI21xp5_ASAP7_75t_L g2533 ( 
.A1(n_2479),
.A2(n_191),
.B(n_193),
.Y(n_2533)
);

NOR3xp33_ASAP7_75t_L g2534 ( 
.A(n_2476),
.B(n_193),
.C(n_194),
.Y(n_2534)
);

NOR3x1_ASAP7_75t_L g2535 ( 
.A(n_2488),
.B(n_194),
.C(n_195),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2472),
.B(n_195),
.Y(n_2536)
);

AOI21xp5_ASAP7_75t_L g2537 ( 
.A1(n_2494),
.A2(n_196),
.B(n_197),
.Y(n_2537)
);

OAI21x1_ASAP7_75t_SL g2538 ( 
.A1(n_2498),
.A2(n_197),
.B(n_198),
.Y(n_2538)
);

OAI21xp5_ASAP7_75t_L g2539 ( 
.A1(n_2497),
.A2(n_198),
.B(n_199),
.Y(n_2539)
);

AOI22xp5_ASAP7_75t_L g2540 ( 
.A1(n_2493),
.A2(n_2147),
.B1(n_2205),
.B2(n_2175),
.Y(n_2540)
);

NOR3x1_ASAP7_75t_L g2541 ( 
.A(n_2480),
.B(n_200),
.C(n_201),
.Y(n_2541)
);

HB1xp67_ASAP7_75t_L g2542 ( 
.A(n_2475),
.Y(n_2542)
);

NAND3xp33_ASAP7_75t_L g2543 ( 
.A(n_2475),
.B(n_200),
.C(n_201),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2475),
.Y(n_2544)
);

OAI21xp5_ASAP7_75t_L g2545 ( 
.A1(n_2471),
.A2(n_202),
.B(n_203),
.Y(n_2545)
);

NOR2xp33_ASAP7_75t_L g2546 ( 
.A(n_2475),
.B(n_202),
.Y(n_2546)
);

INVxp67_ASAP7_75t_L g2547 ( 
.A(n_2504),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2500),
.B(n_203),
.Y(n_2548)
);

NAND4xp25_ASAP7_75t_L g2549 ( 
.A(n_2487),
.B(n_207),
.C(n_205),
.D(n_206),
.Y(n_2549)
);

XNOR2x1_ASAP7_75t_SL g2550 ( 
.A(n_2480),
.B(n_205),
.Y(n_2550)
);

AOI21xp5_ASAP7_75t_L g2551 ( 
.A1(n_2471),
.A2(n_206),
.B(n_207),
.Y(n_2551)
);

NOR3xp33_ASAP7_75t_L g2552 ( 
.A(n_2486),
.B(n_208),
.C(n_209),
.Y(n_2552)
);

AOI21xp33_ASAP7_75t_L g2553 ( 
.A1(n_2471),
.A2(n_208),
.B(n_209),
.Y(n_2553)
);

AOI21xp5_ASAP7_75t_L g2554 ( 
.A1(n_2471),
.A2(n_210),
.B(n_211),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2475),
.Y(n_2555)
);

NOR3xp33_ASAP7_75t_L g2556 ( 
.A(n_2486),
.B(n_210),
.C(n_212),
.Y(n_2556)
);

XNOR2x1_ASAP7_75t_L g2557 ( 
.A(n_2471),
.B(n_212),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2475),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2506),
.Y(n_2559)
);

AOI22xp33_ASAP7_75t_SL g2560 ( 
.A1(n_2487),
.A2(n_2175),
.B1(n_1971),
.B2(n_1934),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2475),
.Y(n_2561)
);

NOR2xp33_ASAP7_75t_L g2562 ( 
.A(n_2475),
.B(n_213),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2475),
.Y(n_2563)
);

AOI22xp5_ASAP7_75t_L g2564 ( 
.A1(n_2473),
.A2(n_2231),
.B1(n_1971),
.B2(n_2188),
.Y(n_2564)
);

NOR3x1_ASAP7_75t_L g2565 ( 
.A(n_2480),
.B(n_214),
.C(n_215),
.Y(n_2565)
);

AOI211x1_ASAP7_75t_L g2566 ( 
.A1(n_2501),
.A2(n_218),
.B(n_216),
.C(n_217),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2500),
.B(n_216),
.Y(n_2567)
);

AOI21xp5_ASAP7_75t_L g2568 ( 
.A1(n_2471),
.A2(n_217),
.B(n_218),
.Y(n_2568)
);

OAI211xp5_ASAP7_75t_SL g2569 ( 
.A1(n_2492),
.A2(n_221),
.B(n_219),
.C(n_220),
.Y(n_2569)
);

NOR3xp33_ASAP7_75t_L g2570 ( 
.A(n_2486),
.B(n_219),
.C(n_220),
.Y(n_2570)
);

OAI21xp33_ASAP7_75t_L g2571 ( 
.A1(n_2487),
.A2(n_2231),
.B(n_2199),
.Y(n_2571)
);

AOI22xp5_ASAP7_75t_L g2572 ( 
.A1(n_2473),
.A2(n_2201),
.B1(n_2184),
.B2(n_2171),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2550),
.Y(n_2573)
);

NOR3xp33_ASAP7_75t_L g2574 ( 
.A(n_2520),
.B(n_221),
.C(n_222),
.Y(n_2574)
);

NAND4xp25_ASAP7_75t_L g2575 ( 
.A(n_2509),
.B(n_225),
.C(n_223),
.D(n_224),
.Y(n_2575)
);

HB1xp67_ASAP7_75t_L g2576 ( 
.A(n_2517),
.Y(n_2576)
);

NOR3xp33_ASAP7_75t_L g2577 ( 
.A(n_2547),
.B(n_2553),
.C(n_2531),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2551),
.B(n_223),
.Y(n_2578)
);

NOR3xp33_ASAP7_75t_L g2579 ( 
.A(n_2545),
.B(n_224),
.C(n_225),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_L g2580 ( 
.A(n_2529),
.B(n_226),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_L g2581 ( 
.A(n_2543),
.B(n_226),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2557),
.Y(n_2582)
);

AOI22xp5_ASAP7_75t_L g2583 ( 
.A1(n_2546),
.A2(n_2171),
.B1(n_2207),
.B2(n_2166),
.Y(n_2583)
);

NOR2xp33_ASAP7_75t_L g2584 ( 
.A(n_2548),
.B(n_228),
.Y(n_2584)
);

AOI211xp5_ASAP7_75t_L g2585 ( 
.A1(n_2569),
.A2(n_2554),
.B(n_2568),
.C(n_2562),
.Y(n_2585)
);

NOR3x1_ASAP7_75t_L g2586 ( 
.A(n_2567),
.B(n_228),
.C(n_229),
.Y(n_2586)
);

NOR3xp33_ASAP7_75t_SL g2587 ( 
.A(n_2521),
.B(n_229),
.C(n_231),
.Y(n_2587)
);

NAND4xp75_ASAP7_75t_L g2588 ( 
.A(n_2535),
.B(n_233),
.C(n_231),
.D(n_232),
.Y(n_2588)
);

NOR2xp33_ASAP7_75t_L g2589 ( 
.A(n_2549),
.B(n_232),
.Y(n_2589)
);

NOR2x1_ASAP7_75t_L g2590 ( 
.A(n_2532),
.B(n_233),
.Y(n_2590)
);

AND3x1_ASAP7_75t_L g2591 ( 
.A(n_2534),
.B(n_234),
.C(n_235),
.Y(n_2591)
);

AOI22xp5_ASAP7_75t_SL g2592 ( 
.A1(n_2510),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_2592)
);

INVx1_ASAP7_75t_SL g2593 ( 
.A(n_2523),
.Y(n_2593)
);

XNOR2x2_ASAP7_75t_L g2594 ( 
.A(n_2566),
.B(n_236),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2541),
.Y(n_2595)
);

OA211x2_ASAP7_75t_L g2596 ( 
.A1(n_2530),
.A2(n_2536),
.B(n_2539),
.C(n_2518),
.Y(n_2596)
);

NOR2xp33_ASAP7_75t_L g2597 ( 
.A(n_2511),
.B(n_237),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2527),
.B(n_2528),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2515),
.B(n_237),
.Y(n_2599)
);

NAND4xp75_ASAP7_75t_L g2600 ( 
.A(n_2522),
.B(n_240),
.C(n_238),
.D(n_239),
.Y(n_2600)
);

NOR2x1_ASAP7_75t_L g2601 ( 
.A(n_2544),
.B(n_238),
.Y(n_2601)
);

NAND3xp33_ASAP7_75t_SL g2602 ( 
.A(n_2525),
.B(n_239),
.C(n_240),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2565),
.Y(n_2603)
);

XNOR2xp5_ASAP7_75t_L g2604 ( 
.A(n_2542),
.B(n_241),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_2555),
.B(n_241),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2514),
.B(n_242),
.Y(n_2606)
);

AND3x2_ASAP7_75t_L g2607 ( 
.A(n_2552),
.B(n_242),
.C(n_243),
.Y(n_2607)
);

NOR2xp67_ASAP7_75t_L g2608 ( 
.A(n_2558),
.B(n_243),
.Y(n_2608)
);

NAND5xp2_ASAP7_75t_L g2609 ( 
.A(n_2526),
.B(n_246),
.C(n_244),
.D(n_245),
.E(n_247),
.Y(n_2609)
);

NOR3xp33_ASAP7_75t_L g2610 ( 
.A(n_2561),
.B(n_244),
.C(n_245),
.Y(n_2610)
);

OAI211xp5_ASAP7_75t_SL g2611 ( 
.A1(n_2563),
.A2(n_249),
.B(n_247),
.C(n_248),
.Y(n_2611)
);

AOI21xp5_ASAP7_75t_L g2612 ( 
.A1(n_2519),
.A2(n_248),
.B(n_249),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2556),
.B(n_250),
.Y(n_2613)
);

AND2x4_ASAP7_75t_L g2614 ( 
.A(n_2559),
.B(n_250),
.Y(n_2614)
);

NOR2x1_ASAP7_75t_L g2615 ( 
.A(n_2537),
.B(n_2533),
.Y(n_2615)
);

NOR3xp33_ASAP7_75t_L g2616 ( 
.A(n_2570),
.B(n_251),
.C(n_252),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2516),
.B(n_251),
.Y(n_2617)
);

OAI22xp5_ASAP7_75t_L g2618 ( 
.A1(n_2512),
.A2(n_2207),
.B1(n_2209),
.B2(n_2166),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2560),
.B(n_253),
.Y(n_2619)
);

NAND3xp33_ASAP7_75t_L g2620 ( 
.A(n_2564),
.B(n_253),
.C(n_254),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2538),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2572),
.Y(n_2622)
);

NOR4xp25_ASAP7_75t_L g2623 ( 
.A(n_2571),
.B(n_257),
.C(n_255),
.D(n_256),
.Y(n_2623)
);

NOR2xp33_ASAP7_75t_L g2624 ( 
.A(n_2540),
.B(n_255),
.Y(n_2624)
);

AOI22xp5_ASAP7_75t_L g2625 ( 
.A1(n_2513),
.A2(n_2220),
.B1(n_2209),
.B2(n_2068),
.Y(n_2625)
);

NAND3xp33_ASAP7_75t_L g2626 ( 
.A(n_2524),
.B(n_257),
.C(n_258),
.Y(n_2626)
);

NOR3xp33_ASAP7_75t_L g2627 ( 
.A(n_2520),
.B(n_258),
.C(n_259),
.Y(n_2627)
);

NOR2x1_ASAP7_75t_L g2628 ( 
.A(n_2531),
.B(n_260),
.Y(n_2628)
);

NOR3xp33_ASAP7_75t_L g2629 ( 
.A(n_2520),
.B(n_260),
.C(n_261),
.Y(n_2629)
);

NOR4xp25_ASAP7_75t_L g2630 ( 
.A(n_2547),
.B(n_264),
.C(n_262),
.D(n_263),
.Y(n_2630)
);

NOR3xp33_ASAP7_75t_L g2631 ( 
.A(n_2520),
.B(n_262),
.C(n_263),
.Y(n_2631)
);

NOR2x1_ASAP7_75t_L g2632 ( 
.A(n_2531),
.B(n_264),
.Y(n_2632)
);

NAND5xp2_ASAP7_75t_L g2633 ( 
.A(n_2509),
.B(n_267),
.C(n_265),
.D(n_266),
.E(n_268),
.Y(n_2633)
);

NOR3xp33_ASAP7_75t_L g2634 ( 
.A(n_2520),
.B(n_265),
.C(n_267),
.Y(n_2634)
);

O2A1O1Ixp33_ASAP7_75t_L g2635 ( 
.A1(n_2547),
.A2(n_271),
.B(n_268),
.C(n_269),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2550),
.Y(n_2636)
);

OAI211xp5_ASAP7_75t_L g2637 ( 
.A1(n_2553),
.A2(n_273),
.B(n_269),
.C(n_272),
.Y(n_2637)
);

NOR4xp75_ASAP7_75t_L g2638 ( 
.A(n_2545),
.B(n_275),
.C(n_272),
.D(n_274),
.Y(n_2638)
);

NOR2x1p5_ASAP7_75t_L g2639 ( 
.A(n_2510),
.B(n_276),
.Y(n_2639)
);

NOR3xp33_ASAP7_75t_L g2640 ( 
.A(n_2520),
.B(n_276),
.C(n_277),
.Y(n_2640)
);

AOI22xp5_ASAP7_75t_L g2641 ( 
.A1(n_2547),
.A2(n_2220),
.B1(n_2069),
.B2(n_2080),
.Y(n_2641)
);

AO22x2_ASAP7_75t_L g2642 ( 
.A1(n_2557),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_2642)
);

NAND4xp25_ASAP7_75t_L g2643 ( 
.A(n_2509),
.B(n_282),
.C(n_278),
.D(n_279),
.Y(n_2643)
);

AND4x1_ASAP7_75t_L g2644 ( 
.A(n_2509),
.B(n_285),
.C(n_283),
.D(n_284),
.Y(n_2644)
);

O2A1O1Ixp5_ASAP7_75t_L g2645 ( 
.A1(n_2553),
.A2(n_287),
.B(n_285),
.C(n_286),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2550),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2614),
.B(n_286),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2642),
.Y(n_2648)
);

OR2x2_ASAP7_75t_L g2649 ( 
.A(n_2630),
.B(n_287),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2614),
.B(n_288),
.Y(n_2650)
);

NAND3xp33_ASAP7_75t_SL g2651 ( 
.A(n_2638),
.B(n_288),
.C(n_289),
.Y(n_2651)
);

NAND2xp33_ASAP7_75t_SL g2652 ( 
.A(n_2587),
.B(n_290),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2608),
.B(n_290),
.Y(n_2653)
);

AND3x2_ASAP7_75t_L g2654 ( 
.A(n_2576),
.B(n_291),
.C(n_292),
.Y(n_2654)
);

NOR2x1_ASAP7_75t_L g2655 ( 
.A(n_2601),
.B(n_291),
.Y(n_2655)
);

NAND4xp75_ASAP7_75t_L g2656 ( 
.A(n_2586),
.B(n_296),
.C(n_294),
.D(n_295),
.Y(n_2656)
);

NAND4xp25_ASAP7_75t_L g2657 ( 
.A(n_2609),
.B(n_297),
.C(n_294),
.D(n_295),
.Y(n_2657)
);

AND3x2_ASAP7_75t_L g2658 ( 
.A(n_2573),
.B(n_297),
.C(n_298),
.Y(n_2658)
);

NOR2x1_ASAP7_75t_L g2659 ( 
.A(n_2636),
.B(n_298),
.Y(n_2659)
);

NOR2x1_ASAP7_75t_L g2660 ( 
.A(n_2646),
.B(n_299),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2642),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2607),
.B(n_299),
.Y(n_2662)
);

NOR3xp33_ASAP7_75t_L g2663 ( 
.A(n_2584),
.B(n_300),
.C(n_301),
.Y(n_2663)
);

NOR3xp33_ASAP7_75t_L g2664 ( 
.A(n_2577),
.B(n_301),
.C(n_302),
.Y(n_2664)
);

AND3x2_ASAP7_75t_L g2665 ( 
.A(n_2580),
.B(n_303),
.C(n_304),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2617),
.Y(n_2666)
);

OAI211xp5_ASAP7_75t_SL g2667 ( 
.A1(n_2585),
.A2(n_306),
.B(n_303),
.C(n_305),
.Y(n_2667)
);

NOR3x1_ASAP7_75t_L g2668 ( 
.A(n_2600),
.B(n_2588),
.C(n_2637),
.Y(n_2668)
);

AOI221x1_ASAP7_75t_L g2669 ( 
.A1(n_2582),
.A2(n_308),
.B1(n_305),
.B2(n_307),
.C(n_309),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2604),
.Y(n_2670)
);

NOR2x1p5_ASAP7_75t_L g2671 ( 
.A(n_2602),
.B(n_307),
.Y(n_2671)
);

OR2x2_ASAP7_75t_L g2672 ( 
.A(n_2633),
.B(n_308),
.Y(n_2672)
);

NOR3x1_ASAP7_75t_L g2673 ( 
.A(n_2575),
.B(n_309),
.C(n_310),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2639),
.Y(n_2674)
);

NOR4xp25_ASAP7_75t_L g2675 ( 
.A(n_2595),
.B(n_312),
.C(n_310),
.D(n_311),
.Y(n_2675)
);

NAND4xp75_ASAP7_75t_L g2676 ( 
.A(n_2628),
.B(n_314),
.C(n_311),
.D(n_312),
.Y(n_2676)
);

OR2x2_ASAP7_75t_L g2677 ( 
.A(n_2643),
.B(n_315),
.Y(n_2677)
);

NAND3xp33_ASAP7_75t_L g2678 ( 
.A(n_2574),
.B(n_315),
.C(n_316),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2594),
.Y(n_2679)
);

AO22x1_ASAP7_75t_L g2680 ( 
.A1(n_2632),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_2680)
);

NOR3xp33_ASAP7_75t_L g2681 ( 
.A(n_2597),
.B(n_317),
.C(n_319),
.Y(n_2681)
);

NOR2x1_ASAP7_75t_L g2682 ( 
.A(n_2598),
.B(n_320),
.Y(n_2682)
);

NAND3xp33_ASAP7_75t_L g2683 ( 
.A(n_2627),
.B(n_320),
.C(n_321),
.Y(n_2683)
);

AOI211xp5_ASAP7_75t_L g2684 ( 
.A1(n_2581),
.A2(n_2589),
.B(n_2616),
.C(n_2579),
.Y(n_2684)
);

NOR3xp33_ASAP7_75t_L g2685 ( 
.A(n_2605),
.B(n_321),
.C(n_322),
.Y(n_2685)
);

NAND3xp33_ASAP7_75t_L g2686 ( 
.A(n_2629),
.B(n_322),
.C(n_323),
.Y(n_2686)
);

AOI221xp5_ASAP7_75t_L g2687 ( 
.A1(n_2623),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.C(n_326),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2644),
.B(n_324),
.Y(n_2688)
);

NAND4xp25_ASAP7_75t_L g2689 ( 
.A(n_2596),
.B(n_327),
.C(n_325),
.D(n_326),
.Y(n_2689)
);

NAND3xp33_ASAP7_75t_SL g2690 ( 
.A(n_2631),
.B(n_327),
.C(n_328),
.Y(n_2690)
);

OAI221xp5_ASAP7_75t_L g2691 ( 
.A1(n_2634),
.A2(n_328),
.B1(n_329),
.B2(n_330),
.C(n_331),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2599),
.Y(n_2692)
);

NOR3xp33_ASAP7_75t_L g2693 ( 
.A(n_2621),
.B(n_329),
.C(n_331),
.Y(n_2693)
);

NOR3xp33_ASAP7_75t_L g2694 ( 
.A(n_2578),
.B(n_332),
.C(n_333),
.Y(n_2694)
);

NOR2x1_ASAP7_75t_L g2695 ( 
.A(n_2603),
.B(n_2611),
.Y(n_2695)
);

NAND3xp33_ASAP7_75t_L g2696 ( 
.A(n_2640),
.B(n_332),
.C(n_333),
.Y(n_2696)
);

NAND4xp25_ASAP7_75t_L g2697 ( 
.A(n_2645),
.B(n_336),
.C(n_334),
.D(n_335),
.Y(n_2697)
);

NOR3xp33_ASAP7_75t_L g2698 ( 
.A(n_2606),
.B(n_334),
.C(n_336),
.Y(n_2698)
);

NOR2x1_ASAP7_75t_L g2699 ( 
.A(n_2590),
.B(n_337),
.Y(n_2699)
);

OAI22xp33_ASAP7_75t_L g2700 ( 
.A1(n_2613),
.A2(n_2619),
.B1(n_2626),
.B2(n_2620),
.Y(n_2700)
);

NAND4xp25_ASAP7_75t_L g2701 ( 
.A(n_2612),
.B(n_339),
.C(n_337),
.D(n_338),
.Y(n_2701)
);

NOR2x1_ASAP7_75t_L g2702 ( 
.A(n_2635),
.B(n_338),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2591),
.Y(n_2703)
);

NOR4xp25_ASAP7_75t_L g2704 ( 
.A(n_2593),
.B(n_341),
.C(n_339),
.D(n_340),
.Y(n_2704)
);

NOR2x1_ASAP7_75t_L g2705 ( 
.A(n_2615),
.B(n_340),
.Y(n_2705)
);

NOR3xp33_ASAP7_75t_L g2706 ( 
.A(n_2610),
.B(n_2622),
.C(n_2624),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_SL g2707 ( 
.A(n_2592),
.B(n_342),
.Y(n_2707)
);

NOR2x1_ASAP7_75t_L g2708 ( 
.A(n_2618),
.B(n_343),
.Y(n_2708)
);

NOR2xp33_ASAP7_75t_L g2709 ( 
.A(n_2583),
.B(n_343),
.Y(n_2709)
);

AND5x1_ASAP7_75t_L g2710 ( 
.A(n_2641),
.B(n_344),
.C(n_345),
.D(n_346),
.E(n_347),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2625),
.Y(n_2711)
);

NAND3xp33_ASAP7_75t_L g2712 ( 
.A(n_2574),
.B(n_344),
.C(n_345),
.Y(n_2712)
);

AOI221xp5_ASAP7_75t_L g2713 ( 
.A1(n_2652),
.A2(n_346),
.B1(n_348),
.B2(n_349),
.C(n_350),
.Y(n_2713)
);

OAI21xp33_ASAP7_75t_L g2714 ( 
.A1(n_2657),
.A2(n_348),
.B(n_349),
.Y(n_2714)
);

BUFx6f_ASAP7_75t_L g2715 ( 
.A(n_2679),
.Y(n_2715)
);

INVxp33_ASAP7_75t_L g2716 ( 
.A(n_2689),
.Y(n_2716)
);

AOI221xp5_ASAP7_75t_L g2717 ( 
.A1(n_2687),
.A2(n_350),
.B1(n_351),
.B2(n_352),
.C(n_353),
.Y(n_2717)
);

AOI32xp33_ASAP7_75t_L g2718 ( 
.A1(n_2695),
.A2(n_351),
.A3(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_2718)
);

AOI22xp5_ASAP7_75t_L g2719 ( 
.A1(n_2651),
.A2(n_356),
.B1(n_354),
.B2(n_355),
.Y(n_2719)
);

O2A1O1Ixp33_ASAP7_75t_L g2720 ( 
.A1(n_2662),
.A2(n_358),
.B(n_356),
.C(n_357),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2665),
.B(n_357),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2705),
.Y(n_2722)
);

NOR2xp67_ASAP7_75t_L g2723 ( 
.A(n_2697),
.B(n_358),
.Y(n_2723)
);

AOI22xp5_ASAP7_75t_SL g2724 ( 
.A1(n_2680),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.Y(n_2724)
);

AOI22x1_ASAP7_75t_L g2725 ( 
.A1(n_2671),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.Y(n_2725)
);

NAND4xp25_ASAP7_75t_SL g2726 ( 
.A(n_2678),
.B(n_364),
.C(n_362),
.D(n_363),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2659),
.Y(n_2727)
);

AOI22xp5_ASAP7_75t_L g2728 ( 
.A1(n_2703),
.A2(n_365),
.B1(n_362),
.B2(n_363),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2673),
.B(n_365),
.Y(n_2729)
);

INVx4_ASAP7_75t_R g2730 ( 
.A(n_2648),
.Y(n_2730)
);

A2O1A1Ixp33_ASAP7_75t_L g2731 ( 
.A1(n_2709),
.A2(n_368),
.B(n_366),
.C(n_367),
.Y(n_2731)
);

AOI22xp5_ASAP7_75t_L g2732 ( 
.A1(n_2694),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.Y(n_2732)
);

OAI211xp5_ASAP7_75t_L g2733 ( 
.A1(n_2704),
.A2(n_2675),
.B(n_2650),
.C(n_2647),
.Y(n_2733)
);

OAI221xp5_ASAP7_75t_SL g2734 ( 
.A1(n_2649),
.A2(n_370),
.B1(n_371),
.B2(n_372),
.C(n_373),
.Y(n_2734)
);

OAI322xp33_ASAP7_75t_L g2735 ( 
.A1(n_2707),
.A2(n_2661),
.A3(n_2700),
.B1(n_2672),
.B2(n_2670),
.C1(n_2674),
.C2(n_2692),
.Y(n_2735)
);

AOI22xp5_ASAP7_75t_L g2736 ( 
.A1(n_2706),
.A2(n_373),
.B1(n_370),
.B2(n_371),
.Y(n_2736)
);

NOR2xp67_ASAP7_75t_L g2737 ( 
.A(n_2701),
.B(n_374),
.Y(n_2737)
);

OAI21xp5_ASAP7_75t_L g2738 ( 
.A1(n_2683),
.A2(n_374),
.B(n_375),
.Y(n_2738)
);

NAND2xp33_ASAP7_75t_SL g2739 ( 
.A(n_2688),
.B(n_376),
.Y(n_2739)
);

AOI31xp33_ASAP7_75t_L g2740 ( 
.A1(n_2699),
.A2(n_379),
.A3(n_377),
.B(n_378),
.Y(n_2740)
);

OAI21xp5_ASAP7_75t_L g2741 ( 
.A1(n_2686),
.A2(n_377),
.B(n_380),
.Y(n_2741)
);

O2A1O1Ixp33_ASAP7_75t_L g2742 ( 
.A1(n_2653),
.A2(n_383),
.B(n_381),
.C(n_382),
.Y(n_2742)
);

NOR3xp33_ASAP7_75t_L g2743 ( 
.A(n_2666),
.B(n_383),
.C(n_384),
.Y(n_2743)
);

HB1xp67_ASAP7_75t_L g2744 ( 
.A(n_2655),
.Y(n_2744)
);

OA211x2_ASAP7_75t_L g2745 ( 
.A1(n_2690),
.A2(n_384),
.B(n_385),
.C(n_386),
.Y(n_2745)
);

NAND3x1_ASAP7_75t_SL g2746 ( 
.A(n_2682),
.B(n_385),
.C(n_386),
.Y(n_2746)
);

NAND3xp33_ASAP7_75t_L g2747 ( 
.A(n_2664),
.B(n_2698),
.C(n_2693),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2668),
.B(n_387),
.Y(n_2748)
);

A2O1A1O1Ixp25_ASAP7_75t_L g2749 ( 
.A1(n_2711),
.A2(n_2691),
.B(n_2702),
.C(n_2684),
.D(n_2710),
.Y(n_2749)
);

AOI221xp5_ASAP7_75t_L g2750 ( 
.A1(n_2696),
.A2(n_387),
.B1(n_388),
.B2(n_389),
.C(n_390),
.Y(n_2750)
);

OAI21xp5_ASAP7_75t_L g2751 ( 
.A1(n_2712),
.A2(n_389),
.B(n_390),
.Y(n_2751)
);

HB1xp67_ASAP7_75t_L g2752 ( 
.A(n_2660),
.Y(n_2752)
);

OAI31xp33_ASAP7_75t_L g2753 ( 
.A1(n_2667),
.A2(n_391),
.A3(n_393),
.B(n_394),
.Y(n_2753)
);

OAI211xp5_ASAP7_75t_SL g2754 ( 
.A1(n_2677),
.A2(n_391),
.B(n_393),
.C(n_395),
.Y(n_2754)
);

XOR2xp5_ASAP7_75t_L g2755 ( 
.A(n_2656),
.B(n_2676),
.Y(n_2755)
);

AOI22xp33_ASAP7_75t_L g2756 ( 
.A1(n_2708),
.A2(n_395),
.B1(n_396),
.B2(n_397),
.Y(n_2756)
);

OAI221xp5_ASAP7_75t_SL g2757 ( 
.A1(n_2663),
.A2(n_2685),
.B1(n_2681),
.B2(n_2658),
.C(n_2669),
.Y(n_2757)
);

O2A1O1Ixp33_ASAP7_75t_L g2758 ( 
.A1(n_2654),
.A2(n_396),
.B(n_398),
.C(n_399),
.Y(n_2758)
);

INVx1_ASAP7_75t_SL g2759 ( 
.A(n_2649),
.Y(n_2759)
);

XNOR2xp5_ASAP7_75t_L g2760 ( 
.A(n_2657),
.B(n_399),
.Y(n_2760)
);

AOI22xp5_ASAP7_75t_L g2761 ( 
.A1(n_2748),
.A2(n_400),
.B1(n_401),
.B2(n_402),
.Y(n_2761)
);

AOI22xp5_ASAP7_75t_L g2762 ( 
.A1(n_2714),
.A2(n_400),
.B1(n_401),
.B2(n_402),
.Y(n_2762)
);

AOI22xp5_ASAP7_75t_L g2763 ( 
.A1(n_2715),
.A2(n_403),
.B1(n_404),
.B2(n_406),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2740),
.B(n_404),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2746),
.Y(n_2765)
);

CKINVDCx5p33_ASAP7_75t_R g2766 ( 
.A(n_2715),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2721),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2724),
.Y(n_2768)
);

AOI22xp5_ASAP7_75t_L g2769 ( 
.A1(n_2715),
.A2(n_407),
.B1(n_408),
.B2(n_409),
.Y(n_2769)
);

NOR2x1_ASAP7_75t_L g2770 ( 
.A(n_2727),
.B(n_407),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2760),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_SL g2772 ( 
.A(n_2719),
.B(n_408),
.Y(n_2772)
);

NOR2x1_ASAP7_75t_L g2773 ( 
.A(n_2722),
.B(n_409),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2729),
.Y(n_2774)
);

AOI22xp5_ASAP7_75t_L g2775 ( 
.A1(n_2723),
.A2(n_410),
.B1(n_411),
.B2(n_412),
.Y(n_2775)
);

AOI22xp5_ASAP7_75t_L g2776 ( 
.A1(n_2737),
.A2(n_410),
.B1(n_411),
.B2(n_412),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2725),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2745),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2755),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2758),
.Y(n_2780)
);

AOI22xp33_ASAP7_75t_SL g2781 ( 
.A1(n_2759),
.A2(n_2733),
.B1(n_2752),
.B2(n_2744),
.Y(n_2781)
);

AND2x4_ASAP7_75t_L g2782 ( 
.A(n_2738),
.B(n_413),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2730),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2728),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2720),
.Y(n_2785)
);

INVxp67_ASAP7_75t_SL g2786 ( 
.A(n_2742),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2754),
.Y(n_2787)
);

AOI22xp5_ASAP7_75t_L g2788 ( 
.A1(n_2726),
.A2(n_413),
.B1(n_414),
.B2(n_415),
.Y(n_2788)
);

AOI22xp5_ASAP7_75t_L g2789 ( 
.A1(n_2739),
.A2(n_415),
.B1(n_416),
.B2(n_417),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2741),
.Y(n_2790)
);

AO22x2_ASAP7_75t_L g2791 ( 
.A1(n_2747),
.A2(n_416),
.B1(n_417),
.B2(n_418),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2751),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2756),
.B(n_418),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2732),
.Y(n_2794)
);

AOI22xp5_ASAP7_75t_L g2795 ( 
.A1(n_2743),
.A2(n_419),
.B1(n_420),
.B2(n_421),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2731),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2734),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2716),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2735),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2749),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2713),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2736),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2757),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_SL g2804 ( 
.A(n_2783),
.B(n_2753),
.Y(n_2804)
);

NAND2x1_ASAP7_75t_L g2805 ( 
.A(n_2773),
.B(n_2718),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2775),
.B(n_2750),
.Y(n_2806)
);

AOI211xp5_ASAP7_75t_L g2807 ( 
.A1(n_2799),
.A2(n_2717),
.B(n_420),
.C(n_421),
.Y(n_2807)
);

CKINVDCx20_ASAP7_75t_R g2808 ( 
.A(n_2766),
.Y(n_2808)
);

BUFx12f_ASAP7_75t_L g2809 ( 
.A(n_2781),
.Y(n_2809)
);

NAND4xp25_ASAP7_75t_L g2810 ( 
.A(n_2800),
.B(n_419),
.C(n_422),
.D(n_423),
.Y(n_2810)
);

NAND3xp33_ASAP7_75t_L g2811 ( 
.A(n_2770),
.B(n_423),
.C(n_424),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2776),
.B(n_424),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2764),
.Y(n_2813)
);

INVx1_ASAP7_75t_SL g2814 ( 
.A(n_2778),
.Y(n_2814)
);

A2O1A1Ixp33_ASAP7_75t_L g2815 ( 
.A1(n_2788),
.A2(n_425),
.B(n_426),
.C(n_427),
.Y(n_2815)
);

INVxp67_ASAP7_75t_L g2816 ( 
.A(n_2761),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2791),
.Y(n_2817)
);

NOR3xp33_ASAP7_75t_L g2818 ( 
.A(n_2803),
.B(n_427),
.C(n_428),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2762),
.Y(n_2819)
);

NOR2x1p5_ASAP7_75t_L g2820 ( 
.A(n_2793),
.B(n_428),
.Y(n_2820)
);

OR2x2_ASAP7_75t_L g2821 ( 
.A(n_2765),
.B(n_429),
.Y(n_2821)
);

NOR2xp67_ASAP7_75t_L g2822 ( 
.A(n_2789),
.B(n_429),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2782),
.Y(n_2823)
);

NAND4xp75_ASAP7_75t_L g2824 ( 
.A(n_2768),
.B(n_430),
.C(n_431),
.D(n_432),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2791),
.Y(n_2825)
);

AOI211x1_ASAP7_75t_L g2826 ( 
.A1(n_2772),
.A2(n_431),
.B(n_432),
.C(n_433),
.Y(n_2826)
);

NOR4xp75_ASAP7_75t_L g2827 ( 
.A(n_2786),
.B(n_433),
.C(n_434),
.D(n_435),
.Y(n_2827)
);

NOR2x1_ASAP7_75t_L g2828 ( 
.A(n_2780),
.B(n_2777),
.Y(n_2828)
);

NAND2xp33_ASAP7_75t_R g2829 ( 
.A(n_2785),
.B(n_434),
.Y(n_2829)
);

AOI21xp5_ASAP7_75t_SL g2830 ( 
.A1(n_2787),
.A2(n_435),
.B(n_436),
.Y(n_2830)
);

HB1xp67_ASAP7_75t_L g2831 ( 
.A(n_2795),
.Y(n_2831)
);

AND2x4_ASAP7_75t_L g2832 ( 
.A(n_2774),
.B(n_436),
.Y(n_2832)
);

OAI21xp33_ASAP7_75t_L g2833 ( 
.A1(n_2814),
.A2(n_2798),
.B(n_2779),
.Y(n_2833)
);

AOI221xp5_ASAP7_75t_L g2834 ( 
.A1(n_2826),
.A2(n_2797),
.B1(n_2801),
.B2(n_2802),
.C(n_2790),
.Y(n_2834)
);

OAI22xp33_ASAP7_75t_SL g2835 ( 
.A1(n_2805),
.A2(n_2796),
.B1(n_2792),
.B2(n_2767),
.Y(n_2835)
);

AOI22xp5_ASAP7_75t_L g2836 ( 
.A1(n_2809),
.A2(n_2784),
.B1(n_2794),
.B2(n_2771),
.Y(n_2836)
);

NAND4xp75_ASAP7_75t_L g2837 ( 
.A(n_2828),
.B(n_2769),
.C(n_2763),
.D(n_439),
.Y(n_2837)
);

OAI321xp33_ASAP7_75t_L g2838 ( 
.A1(n_2807),
.A2(n_437),
.A3(n_438),
.B1(n_439),
.B2(n_440),
.C(n_441),
.Y(n_2838)
);

AOI21xp5_ASAP7_75t_L g2839 ( 
.A1(n_2804),
.A2(n_437),
.B(n_438),
.Y(n_2839)
);

AOI322xp5_ASAP7_75t_L g2840 ( 
.A1(n_2808),
.A2(n_440),
.A3(n_442),
.B1(n_443),
.B2(n_444),
.C1(n_445),
.C2(n_446),
.Y(n_2840)
);

AND2x4_ASAP7_75t_SL g2841 ( 
.A(n_2823),
.B(n_442),
.Y(n_2841)
);

INVx1_ASAP7_75t_SL g2842 ( 
.A(n_2821),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2820),
.B(n_443),
.Y(n_2843)
);

AO21x1_ASAP7_75t_L g2844 ( 
.A1(n_2829),
.A2(n_445),
.B(n_446),
.Y(n_2844)
);

AND2x2_ASAP7_75t_L g2845 ( 
.A(n_2818),
.B(n_447),
.Y(n_2845)
);

OAI221xp5_ASAP7_75t_L g2846 ( 
.A1(n_2815),
.A2(n_448),
.B1(n_449),
.B2(n_450),
.C(n_451),
.Y(n_2846)
);

NAND3xp33_ASAP7_75t_L g2847 ( 
.A(n_2811),
.B(n_449),
.C(n_452),
.Y(n_2847)
);

AOI31xp33_ASAP7_75t_L g2848 ( 
.A1(n_2817),
.A2(n_452),
.A3(n_453),
.B(n_454),
.Y(n_2848)
);

NOR2xp33_ASAP7_75t_L g2849 ( 
.A(n_2812),
.B(n_453),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2827),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2830),
.B(n_455),
.Y(n_2851)
);

NOR2x1_ASAP7_75t_L g2852 ( 
.A(n_2824),
.B(n_455),
.Y(n_2852)
);

NOR2x1_ASAP7_75t_L g2853 ( 
.A(n_2825),
.B(n_456),
.Y(n_2853)
);

AND2x4_ASAP7_75t_L g2854 ( 
.A(n_2822),
.B(n_456),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2832),
.Y(n_2855)
);

OAI221xp5_ASAP7_75t_L g2856 ( 
.A1(n_2816),
.A2(n_457),
.B1(n_458),
.B2(n_460),
.C(n_462),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2832),
.Y(n_2857)
);

AND2x4_ASAP7_75t_L g2858 ( 
.A(n_2819),
.B(n_457),
.Y(n_2858)
);

OAI21xp5_ASAP7_75t_SL g2859 ( 
.A1(n_2806),
.A2(n_2831),
.B(n_2813),
.Y(n_2859)
);

AOI22xp5_ASAP7_75t_L g2860 ( 
.A1(n_2810),
.A2(n_458),
.B1(n_460),
.B2(n_463),
.Y(n_2860)
);

NAND3xp33_ASAP7_75t_L g2861 ( 
.A(n_2818),
.B(n_464),
.C(n_465),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2827),
.Y(n_2862)
);

INVxp67_ASAP7_75t_L g2863 ( 
.A(n_2829),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2818),
.B(n_464),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2853),
.Y(n_2865)
);

INVx4_ASAP7_75t_L g2866 ( 
.A(n_2855),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2841),
.Y(n_2867)
);

OAI22xp5_ASAP7_75t_L g2868 ( 
.A1(n_2860),
.A2(n_465),
.B1(n_466),
.B2(n_467),
.Y(n_2868)
);

INVx2_ASAP7_75t_SL g2869 ( 
.A(n_2843),
.Y(n_2869)
);

NOR2xp33_ASAP7_75t_L g2870 ( 
.A(n_2851),
.B(n_466),
.Y(n_2870)
);

NOR2x1_ASAP7_75t_L g2871 ( 
.A(n_2857),
.B(n_468),
.Y(n_2871)
);

NOR2x1p5_ASAP7_75t_L g2872 ( 
.A(n_2837),
.B(n_468),
.Y(n_2872)
);

BUFx2_ASAP7_75t_L g2873 ( 
.A(n_2844),
.Y(n_2873)
);

AOI31xp33_ASAP7_75t_L g2874 ( 
.A1(n_2863),
.A2(n_469),
.A3(n_470),
.B(n_471),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2852),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2849),
.Y(n_2876)
);

XNOR2x1_ASAP7_75t_L g2877 ( 
.A(n_2836),
.B(n_469),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2847),
.Y(n_2878)
);

OAI211xp5_ASAP7_75t_L g2879 ( 
.A1(n_2833),
.A2(n_470),
.B(n_471),
.C(n_472),
.Y(n_2879)
);

AOI211xp5_ASAP7_75t_L g2880 ( 
.A1(n_2835),
.A2(n_472),
.B(n_473),
.C(n_474),
.Y(n_2880)
);

OR3x2_ASAP7_75t_L g2881 ( 
.A(n_2850),
.B(n_473),
.C(n_474),
.Y(n_2881)
);

XNOR2x1_ASAP7_75t_L g2882 ( 
.A(n_2854),
.B(n_2862),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2861),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2858),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2881),
.Y(n_2885)
);

AO21x2_ASAP7_75t_L g2886 ( 
.A1(n_2865),
.A2(n_2859),
.B(n_2839),
.Y(n_2886)
);

XOR2x2_ASAP7_75t_L g2887 ( 
.A(n_2877),
.B(n_2834),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2880),
.B(n_2845),
.Y(n_2888)
);

AOI21xp33_ASAP7_75t_L g2889 ( 
.A1(n_2870),
.A2(n_2842),
.B(n_2864),
.Y(n_2889)
);

XNOR2x1_ASAP7_75t_L g2890 ( 
.A(n_2882),
.B(n_2838),
.Y(n_2890)
);

AO22x2_ASAP7_75t_L g2891 ( 
.A1(n_2884),
.A2(n_2858),
.B1(n_2846),
.B2(n_2848),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2871),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2868),
.B(n_2840),
.Y(n_2893)
);

AO21x2_ASAP7_75t_L g2894 ( 
.A1(n_2875),
.A2(n_2856),
.B(n_476),
.Y(n_2894)
);

INVxp67_ASAP7_75t_SL g2895 ( 
.A(n_2872),
.Y(n_2895)
);

INVxp67_ASAP7_75t_L g2896 ( 
.A(n_2873),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2867),
.Y(n_2897)
);

NAND3xp33_ASAP7_75t_L g2898 ( 
.A(n_2866),
.B(n_475),
.C(n_476),
.Y(n_2898)
);

HB1xp67_ASAP7_75t_L g2899 ( 
.A(n_2894),
.Y(n_2899)
);

OAI22xp5_ASAP7_75t_L g2900 ( 
.A1(n_2896),
.A2(n_2878),
.B1(n_2883),
.B2(n_2869),
.Y(n_2900)
);

OA22x2_ASAP7_75t_L g2901 ( 
.A1(n_2892),
.A2(n_2879),
.B1(n_2876),
.B2(n_2874),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2891),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2898),
.Y(n_2903)
);

AO22x2_ASAP7_75t_L g2904 ( 
.A1(n_2890),
.A2(n_477),
.B1(n_478),
.B2(n_479),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2885),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2897),
.Y(n_2906)
);

OAI22x1_ASAP7_75t_L g2907 ( 
.A1(n_2895),
.A2(n_478),
.B1(n_479),
.B2(n_480),
.Y(n_2907)
);

OAI22xp5_ASAP7_75t_L g2908 ( 
.A1(n_2906),
.A2(n_2893),
.B1(n_2888),
.B2(n_2889),
.Y(n_2908)
);

XNOR2x1_ASAP7_75t_L g2909 ( 
.A(n_2900),
.B(n_2887),
.Y(n_2909)
);

XOR2xp5_ASAP7_75t_L g2910 ( 
.A(n_2901),
.B(n_2886),
.Y(n_2910)
);

NAND4xp25_ASAP7_75t_L g2911 ( 
.A(n_2902),
.B(n_480),
.C(n_481),
.D(n_482),
.Y(n_2911)
);

AOI22xp5_ASAP7_75t_L g2912 ( 
.A1(n_2905),
.A2(n_481),
.B1(n_482),
.B2(n_483),
.Y(n_2912)
);

OAI221xp5_ASAP7_75t_L g2913 ( 
.A1(n_2910),
.A2(n_2899),
.B1(n_2903),
.B2(n_2904),
.C(n_2907),
.Y(n_2913)
);

AND2x4_ASAP7_75t_L g2914 ( 
.A(n_2912),
.B(n_486),
.Y(n_2914)
);

INVx4_ASAP7_75t_L g2915 ( 
.A(n_2909),
.Y(n_2915)
);

OAI221xp5_ASAP7_75t_R g2916 ( 
.A1(n_2908),
.A2(n_486),
.B1(n_487),
.B2(n_488),
.C(n_489),
.Y(n_2916)
);

AOI21xp5_ASAP7_75t_L g2917 ( 
.A1(n_2911),
.A2(n_488),
.B(n_489),
.Y(n_2917)
);

HB1xp67_ASAP7_75t_L g2918 ( 
.A(n_2915),
.Y(n_2918)
);

INVx2_ASAP7_75t_SL g2919 ( 
.A(n_2914),
.Y(n_2919)
);

BUFx2_ASAP7_75t_L g2920 ( 
.A(n_2916),
.Y(n_2920)
);

AO21x2_ASAP7_75t_L g2921 ( 
.A1(n_2918),
.A2(n_2913),
.B(n_2917),
.Y(n_2921)
);

OAI21xp5_ASAP7_75t_L g2922 ( 
.A1(n_2920),
.A2(n_490),
.B(n_491),
.Y(n_2922)
);

AOI22xp33_ASAP7_75t_L g2923 ( 
.A1(n_2919),
.A2(n_490),
.B1(n_492),
.B2(n_493),
.Y(n_2923)
);

XNOR2xp5_ASAP7_75t_L g2924 ( 
.A(n_2921),
.B(n_492),
.Y(n_2924)
);

OAI21xp33_ASAP7_75t_SL g2925 ( 
.A1(n_2922),
.A2(n_493),
.B(n_494),
.Y(n_2925)
);

OAI22xp5_ASAP7_75t_L g2926 ( 
.A1(n_2924),
.A2(n_2925),
.B1(n_2923),
.B2(n_497),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2925),
.B(n_495),
.Y(n_2927)
);

AOI22xp5_ASAP7_75t_L g2928 ( 
.A1(n_2925),
.A2(n_495),
.B1(n_496),
.B2(n_497),
.Y(n_2928)
);

NOR2x1_ASAP7_75t_SL g2929 ( 
.A(n_2926),
.B(n_496),
.Y(n_2929)
);

AOI22xp5_ASAP7_75t_L g2930 ( 
.A1(n_2929),
.A2(n_2927),
.B1(n_2928),
.B2(n_502),
.Y(n_2930)
);

OA21x2_ASAP7_75t_L g2931 ( 
.A1(n_2930),
.A2(n_499),
.B(n_500),
.Y(n_2931)
);

AOI221xp5_ASAP7_75t_L g2932 ( 
.A1(n_2931),
.A2(n_500),
.B1(n_502),
.B2(n_503),
.C(n_504),
.Y(n_2932)
);

AOI21xp33_ASAP7_75t_SL g2933 ( 
.A1(n_2932),
.A2(n_503),
.B(n_504),
.Y(n_2933)
);

AOI211xp5_ASAP7_75t_L g2934 ( 
.A1(n_2933),
.A2(n_505),
.B(n_506),
.C(n_507),
.Y(n_2934)
);


endmodule