module fake_netlist_1_4557_n_476 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_476);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_476;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g71 ( .A(n_54), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_37), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_51), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_28), .Y(n_74) );
INVx2_ASAP7_75t_L g75 ( .A(n_18), .Y(n_75) );
INVx2_ASAP7_75t_L g76 ( .A(n_23), .Y(n_76) );
INVxp33_ASAP7_75t_L g77 ( .A(n_10), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_36), .Y(n_78) );
INVxp33_ASAP7_75t_SL g79 ( .A(n_33), .Y(n_79) );
NOR2xp67_ASAP7_75t_L g80 ( .A(n_14), .B(n_42), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_49), .Y(n_81) );
CKINVDCx14_ASAP7_75t_R g82 ( .A(n_7), .Y(n_82) );
INVxp33_ASAP7_75t_SL g83 ( .A(n_67), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_46), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_65), .Y(n_85) );
INVxp67_ASAP7_75t_L g86 ( .A(n_10), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_62), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_32), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_61), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_12), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_59), .Y(n_91) );
INVx1_ASAP7_75t_SL g92 ( .A(n_45), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_57), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_31), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_14), .Y(n_95) );
CKINVDCx16_ASAP7_75t_R g96 ( .A(n_69), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_12), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_52), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_19), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_1), .Y(n_100) );
CKINVDCx14_ASAP7_75t_R g101 ( .A(n_6), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_60), .Y(n_102) );
CKINVDCx12_ASAP7_75t_R g103 ( .A(n_16), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_47), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_76), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_75), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_77), .B(n_0), .Y(n_107) );
AND2x4_ASAP7_75t_L g108 ( .A(n_75), .B(n_0), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_76), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_76), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_1), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_94), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_99), .B(n_2), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_94), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_82), .B(n_2), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_82), .Y(n_116) );
AND2x2_ASAP7_75t_L g117 ( .A(n_71), .B(n_3), .Y(n_117) );
NAND2xp33_ASAP7_75t_L g118 ( .A(n_94), .B(n_70), .Y(n_118) );
AND2x4_ASAP7_75t_L g119 ( .A(n_75), .B(n_3), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_102), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_90), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_90), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_102), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_101), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_102), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_72), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_72), .Y(n_127) );
NAND3x1_ASAP7_75t_L g128 ( .A(n_117), .B(n_100), .C(n_97), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_126), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_108), .A2(n_100), .B1(n_95), .B2(n_97), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_126), .Y(n_131) );
BUFx10_ASAP7_75t_L g132 ( .A(n_124), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_117), .B(n_71), .Y(n_133) );
INVx3_ASAP7_75t_L g134 ( .A(n_108), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_126), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_126), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_127), .B(n_96), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_120), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_120), .Y(n_139) );
AND2x6_ASAP7_75t_L g140 ( .A(n_108), .B(n_73), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_116), .A2(n_96), .B1(n_86), .B2(n_95), .Y(n_141) );
AND2x6_ASAP7_75t_L g142 ( .A(n_108), .B(n_78), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_120), .Y(n_143) );
OR2x2_ASAP7_75t_L g144 ( .A(n_111), .B(n_86), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_120), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_126), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_120), .Y(n_147) );
BUFx3_ASAP7_75t_L g148 ( .A(n_120), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_127), .B(n_104), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_127), .B(n_79), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_119), .B(n_90), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_123), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_126), .Y(n_153) );
XOR2xp5_ASAP7_75t_L g154 ( .A(n_141), .B(n_113), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_134), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_133), .B(n_115), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g157 ( .A1(n_140), .A2(n_119), .B1(n_115), .B2(n_107), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_137), .B(n_119), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_144), .B(n_83), .Y(n_159) );
INVx1_ASAP7_75t_SL g160 ( .A(n_132), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_134), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_140), .Y(n_162) );
AND2x2_ASAP7_75t_SL g163 ( .A(n_151), .B(n_119), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_140), .A2(n_103), .B1(n_93), .B2(n_85), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_144), .B(n_92), .Y(n_165) );
NOR2x1p5_ASAP7_75t_L g166 ( .A(n_132), .B(n_85), .Y(n_166) );
NAND2xp33_ASAP7_75t_R g167 ( .A(n_134), .B(n_87), .Y(n_167) );
INVx1_ASAP7_75t_SL g168 ( .A(n_132), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_134), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_151), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_150), .B(n_121), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_151), .B(n_80), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_143), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_140), .A2(n_125), .B1(n_123), .B2(n_112), .Y(n_174) );
BUFx3_ASAP7_75t_L g175 ( .A(n_140), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_140), .A2(n_118), .B1(n_73), .B2(n_78), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_140), .B(n_121), .Y(n_177) );
INVx2_ASAP7_75t_SL g178 ( .A(n_132), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g180 ( .A1(n_130), .A2(n_112), .B(n_105), .C(n_109), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_140), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_142), .B(n_80), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g183 ( .A1(n_128), .A2(n_105), .B1(n_114), .B2(n_110), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
BUFx2_ASAP7_75t_L g185 ( .A(n_142), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_142), .A2(n_74), .B1(n_81), .B2(n_84), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_147), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_155), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_163), .A2(n_142), .B1(n_156), .B2(n_179), .Y(n_189) );
BUFx2_ASAP7_75t_L g190 ( .A(n_162), .Y(n_190) );
INVxp67_ASAP7_75t_L g191 ( .A(n_160), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_156), .B(n_142), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_163), .A2(n_142), .B1(n_128), .B2(n_149), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_165), .B(n_142), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_159), .B(n_178), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_155), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_162), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_162), .Y(n_198) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_168), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_157), .A2(n_142), .B1(n_114), .B2(n_110), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_161), .Y(n_201) );
INVx2_ASAP7_75t_SL g202 ( .A(n_175), .Y(n_202) );
INVx11_ASAP7_75t_L g203 ( .A(n_178), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_161), .Y(n_204) );
BUFx2_ASAP7_75t_L g205 ( .A(n_185), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_181), .A2(n_92), .B1(n_105), .B2(n_109), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_158), .A2(n_114), .B(n_110), .C(n_109), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_170), .B(n_121), .Y(n_208) );
OR2x2_ASAP7_75t_L g209 ( .A(n_154), .B(n_121), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_169), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_169), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_166), .Y(n_212) );
CKINVDCx8_ASAP7_75t_R g213 ( .A(n_185), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_175), .Y(n_214) );
INVx3_ASAP7_75t_L g215 ( .A(n_170), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_179), .Y(n_216) );
OAI21x1_ASAP7_75t_SL g217 ( .A1(n_186), .A2(n_74), .B(n_81), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_181), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_184), .Y(n_219) );
INVx6_ASAP7_75t_L g220 ( .A(n_172), .Y(n_220) );
OAI211xp5_ASAP7_75t_L g221 ( .A1(n_193), .A2(n_164), .B(n_154), .C(n_171), .Y(n_221) );
INVx4_ASAP7_75t_L g222 ( .A(n_198), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_192), .B(n_166), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_196), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_192), .B(n_172), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_198), .Y(n_226) );
OAI21x1_ASAP7_75t_L g227 ( .A1(n_217), .A2(n_180), .B(n_174), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_196), .Y(n_228) );
INVxp67_ASAP7_75t_L g229 ( .A(n_199), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_190), .B(n_172), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_196), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_201), .Y(n_232) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_200), .A2(n_177), .B(n_176), .Y(n_233) );
OAI22xp33_ASAP7_75t_L g234 ( .A1(n_209), .A2(n_167), .B1(n_183), .B2(n_182), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_209), .A2(n_182), .B1(n_187), .B2(n_184), .Y(n_235) );
AOI22xp33_ASAP7_75t_SL g236 ( .A1(n_191), .A2(n_182), .B1(n_84), .B2(n_89), .Y(n_236) );
INVx1_ASAP7_75t_SL g237 ( .A(n_220), .Y(n_237) );
BUFx2_ASAP7_75t_L g238 ( .A(n_205), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_201), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_189), .A2(n_187), .B1(n_89), .B2(n_91), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_201), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_204), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_203), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_193), .B(n_106), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_205), .B(n_106), .Y(n_245) );
OAI21x1_ASAP7_75t_SL g246 ( .A1(n_241), .A2(n_224), .B(n_228), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_234), .A2(n_195), .B1(n_220), .B2(n_212), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_241), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_226), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_223), .A2(n_220), .B1(n_217), .B2(n_194), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_221), .A2(n_200), .B(n_207), .C(n_215), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_222), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_224), .A2(n_213), .B1(n_203), .B2(n_218), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_228), .B(n_216), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_241), .Y(n_255) );
AOI22xp33_ASAP7_75t_SL g256 ( .A1(n_238), .A2(n_220), .B1(n_218), .B2(n_190), .Y(n_256) );
NOR2x1_ASAP7_75t_L g257 ( .A(n_231), .B(n_206), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_231), .B(n_216), .Y(n_258) );
AOI221xp5_ASAP7_75t_L g259 ( .A1(n_229), .A2(n_208), .B1(n_188), .B2(n_210), .C(n_211), .Y(n_259) );
OAI211xp5_ASAP7_75t_L g260 ( .A1(n_236), .A2(n_122), .B(n_91), .C(n_98), .Y(n_260) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_227), .A2(n_145), .B(n_139), .Y(n_261) );
INVx1_ASAP7_75t_SL g262 ( .A(n_238), .Y(n_262) );
OAI211xp5_ASAP7_75t_SL g263 ( .A1(n_235), .A2(n_122), .B(n_98), .C(n_153), .Y(n_263) );
AOI221xp5_ASAP7_75t_L g264 ( .A1(n_240), .A2(n_188), .B1(n_210), .B2(n_211), .C(n_215), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_232), .A2(n_213), .B1(n_220), .B2(n_204), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_223), .B(n_215), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_265), .A2(n_232), .B1(n_239), .B2(n_242), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_246), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_248), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_252), .B(n_239), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_248), .Y(n_271) );
AOI22xp33_ASAP7_75t_SL g272 ( .A1(n_253), .A2(n_223), .B1(n_230), .B2(n_225), .Y(n_272) );
OAI222xp33_ASAP7_75t_L g273 ( .A1(n_262), .A2(n_242), .B1(n_244), .B2(n_223), .C1(n_230), .C2(n_245), .Y(n_273) );
AOI33xp33_ASAP7_75t_L g274 ( .A1(n_247), .A2(n_245), .A3(n_237), .B1(n_225), .B2(n_129), .B3(n_131), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_262), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_248), .B(n_230), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_246), .Y(n_277) );
INVxp67_ASAP7_75t_L g278 ( .A(n_258), .Y(n_278) );
NAND4xp25_ASAP7_75t_SL g279 ( .A(n_256), .B(n_243), .C(n_233), .D(n_6), .Y(n_279) );
OAI21x1_ASAP7_75t_L g280 ( .A1(n_261), .A2(n_227), .B(n_219), .Y(n_280) );
INVx4_ASAP7_75t_L g281 ( .A(n_252), .Y(n_281) );
OAI211xp5_ASAP7_75t_L g282 ( .A1(n_260), .A2(n_222), .B(n_88), .C(n_125), .Y(n_282) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_255), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_255), .B(n_258), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_255), .Y(n_285) );
OAI22xp33_ASAP7_75t_L g286 ( .A1(n_259), .A2(n_230), .B1(n_222), .B2(n_225), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_250), .A2(n_225), .B1(n_222), .B2(n_204), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_254), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_270), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_284), .B(n_252), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_269), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_284), .B(n_252), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_285), .B(n_254), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_285), .B(n_254), .Y(n_294) );
BUFx2_ASAP7_75t_L g295 ( .A(n_268), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_277), .Y(n_296) );
NAND3xp33_ASAP7_75t_L g297 ( .A(n_277), .B(n_251), .C(n_257), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_275), .B(n_254), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_288), .B(n_261), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_269), .B(n_261), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_279), .A2(n_263), .B1(n_266), .B2(n_257), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_271), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_271), .B(n_261), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_283), .B(n_249), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_288), .Y(n_305) );
OAI33xp33_ASAP7_75t_L g306 ( .A1(n_286), .A2(n_129), .A3(n_131), .B1(n_135), .B2(n_136), .B3(n_146), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_270), .B(n_249), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g308 ( .A1(n_278), .A2(n_264), .B1(n_215), .B2(n_123), .C(n_125), .Y(n_308) );
AOI33xp33_ASAP7_75t_L g309 ( .A1(n_272), .A2(n_135), .A3(n_136), .B1(n_146), .B2(n_153), .B3(n_145), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_273), .B(n_4), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_267), .A2(n_249), .B1(n_226), .B2(n_219), .Y(n_311) );
OAI31xp33_ASAP7_75t_L g312 ( .A1(n_267), .A2(n_197), .A3(n_219), .B(n_202), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_270), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_270), .B(n_249), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_276), .B(n_249), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_276), .B(n_249), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g317 ( .A1(n_287), .A2(n_226), .B1(n_219), .B2(n_197), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_281), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_281), .B(n_226), .Y(n_319) );
CKINVDCx16_ASAP7_75t_R g320 ( .A(n_289), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_305), .B(n_281), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_293), .B(n_274), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_313), .B(n_281), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_293), .B(n_280), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_318), .B(n_282), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_305), .B(n_280), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_296), .B(n_123), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_319), .Y(n_328) );
OAI22xp33_ASAP7_75t_L g329 ( .A1(n_318), .A2(n_226), .B1(n_197), .B2(n_198), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_294), .B(n_4), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_289), .Y(n_331) );
AOI21xp33_ASAP7_75t_L g332 ( .A1(n_310), .A2(n_123), .B(n_125), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_294), .B(n_5), .Y(n_333) );
NAND3xp33_ASAP7_75t_L g334 ( .A(n_301), .B(n_123), .C(n_125), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_296), .B(n_125), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_302), .Y(n_336) );
INVx1_ASAP7_75t_SL g337 ( .A(n_319), .Y(n_337) );
NAND4xp25_ASAP7_75t_L g338 ( .A(n_301), .B(n_138), .C(n_139), .D(n_145), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_298), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_298), .B(n_5), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_290), .B(n_7), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_290), .B(n_8), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_292), .B(n_8), .Y(n_343) );
NOR3xp33_ASAP7_75t_L g344 ( .A(n_309), .B(n_138), .C(n_139), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_291), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_307), .B(n_9), .Y(n_346) );
AOI211x1_ASAP7_75t_L g347 ( .A1(n_297), .A2(n_9), .B(n_11), .C(n_13), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_291), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_295), .Y(n_349) );
OAI32xp33_ASAP7_75t_L g350 ( .A1(n_313), .A2(n_11), .A3(n_13), .B1(n_15), .B2(n_16), .Y(n_350) );
NOR3xp33_ASAP7_75t_L g351 ( .A(n_306), .B(n_138), .C(n_214), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_292), .B(n_15), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_307), .B(n_17), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_314), .B(n_17), .Y(n_354) );
INVx1_ASAP7_75t_SL g355 ( .A(n_289), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_314), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_299), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_300), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_304), .B(n_18), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_304), .B(n_19), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_316), .B(n_315), .Y(n_361) );
OA211x2_ASAP7_75t_L g362 ( .A1(n_325), .A2(n_312), .B(n_308), .C(n_311), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_361), .B(n_316), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_339), .B(n_303), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_357), .B(n_300), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_320), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_361), .B(n_315), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_328), .B(n_299), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_340), .B(n_306), .Y(n_369) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_345), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_359), .B(n_297), .Y(n_371) );
OAI31xp33_ASAP7_75t_L g372 ( .A1(n_352), .A2(n_312), .A3(n_308), .B(n_317), .Y(n_372) );
AOI211xp5_ASAP7_75t_SL g373 ( .A1(n_359), .A2(n_317), .B(n_197), .C(n_214), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_360), .B(n_152), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_358), .B(n_152), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_358), .B(n_152), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_337), .B(n_226), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_356), .B(n_326), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_331), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_326), .B(n_152), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_336), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_320), .Y(n_382) );
OAI21xp33_ASAP7_75t_L g383 ( .A1(n_349), .A2(n_152), .B(n_143), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_360), .B(n_152), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_341), .B(n_342), .Y(n_385) );
NAND4xp25_ASAP7_75t_L g386 ( .A(n_347), .B(n_148), .C(n_147), .D(n_214), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_331), .B(n_20), .Y(n_387) );
NOR2xp67_ASAP7_75t_SL g388 ( .A(n_334), .B(n_198), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_324), .B(n_321), .Y(n_389) );
NOR2x1p5_ASAP7_75t_L g390 ( .A(n_352), .B(n_143), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_341), .B(n_143), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_342), .B(n_143), .Y(n_392) );
OAI21xp5_ASAP7_75t_SL g393 ( .A1(n_346), .A2(n_198), .B(n_22), .Y(n_393) );
XNOR2xp5_ASAP7_75t_L g394 ( .A(n_346), .B(n_21), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_353), .B(n_148), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_322), .B(n_24), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_321), .B(n_25), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_353), .B(n_26), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_363), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_363), .Y(n_400) );
NOR3xp33_ASAP7_75t_L g401 ( .A(n_386), .B(n_350), .C(n_338), .Y(n_401) );
INVx3_ASAP7_75t_L g402 ( .A(n_366), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_382), .B(n_355), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_367), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_389), .B(n_354), .Y(n_405) );
NOR2xp67_ASAP7_75t_L g406 ( .A(n_393), .B(n_323), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_389), .B(n_354), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_378), .B(n_323), .Y(n_408) );
NOR2x1_ASAP7_75t_L g409 ( .A(n_390), .B(n_329), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_371), .B(n_335), .Y(n_410) );
OAI21xp33_ASAP7_75t_L g411 ( .A1(n_379), .A2(n_343), .B(n_330), .Y(n_411) );
XNOR2xp5_ASAP7_75t_L g412 ( .A(n_394), .B(n_333), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_378), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_365), .B(n_348), .Y(n_414) );
NAND4xp25_ASAP7_75t_L g415 ( .A(n_362), .B(n_332), .C(n_327), .D(n_344), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_387), .B(n_327), .Y(n_416) );
NAND2x1p5_ASAP7_75t_L g417 ( .A(n_387), .B(n_198), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_381), .B(n_351), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_368), .Y(n_419) );
XOR2x2_ASAP7_75t_L g420 ( .A(n_385), .B(n_27), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_387), .B(n_173), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_364), .B(n_29), .Y(n_422) );
OAI21xp5_ASAP7_75t_SL g423 ( .A1(n_373), .A2(n_30), .B(n_34), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_369), .B(n_35), .Y(n_424) );
NOR3xp33_ASAP7_75t_L g425 ( .A(n_396), .B(n_38), .C(n_39), .Y(n_425) );
NAND5xp2_ASAP7_75t_L g426 ( .A(n_372), .B(n_40), .C(n_41), .D(n_43), .E(n_44), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_370), .B(n_48), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_370), .B(n_50), .Y(n_428) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_369), .A2(n_173), .B1(n_55), .B2(n_56), .C(n_58), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_380), .B(n_53), .Y(n_430) );
OAI21xp5_ASAP7_75t_L g431 ( .A1(n_397), .A2(n_63), .B(n_64), .Y(n_431) );
XNOR2x1_ASAP7_75t_L g432 ( .A(n_397), .B(n_66), .Y(n_432) );
OAI21xp33_ASAP7_75t_L g433 ( .A1(n_396), .A2(n_173), .B(n_68), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_398), .A2(n_374), .B1(n_384), .B2(n_391), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_392), .A2(n_173), .B1(n_395), .B2(n_375), .Y(n_435) );
OAI22xp33_ASAP7_75t_L g436 ( .A1(n_388), .A2(n_393), .B1(n_373), .B2(n_382), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_383), .A2(n_393), .B(n_373), .Y(n_437) );
AOI21xp33_ASAP7_75t_SL g438 ( .A1(n_376), .A2(n_394), .B(n_382), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_363), .Y(n_439) );
AOI21xp33_ASAP7_75t_L g440 ( .A1(n_369), .A2(n_396), .B(n_394), .Y(n_440) );
NOR3xp33_ASAP7_75t_L g441 ( .A(n_386), .B(n_279), .C(n_396), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_389), .B(n_378), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_393), .A2(n_362), .B1(n_369), .B2(n_390), .Y(n_443) );
NOR2x1p5_ASAP7_75t_SL g444 ( .A(n_377), .B(n_352), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_366), .B(n_382), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_363), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_443), .A2(n_445), .B1(n_406), .B2(n_441), .Y(n_447) );
OAI22xp33_ASAP7_75t_L g448 ( .A1(n_402), .A2(n_437), .B1(n_438), .B2(n_417), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_440), .A2(n_411), .B1(n_407), .B2(n_405), .C(n_404), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g450 ( .A1(n_440), .A2(n_400), .B1(n_439), .B2(n_399), .C(n_446), .Y(n_450) );
INVxp67_ASAP7_75t_L g451 ( .A(n_418), .Y(n_451) );
NOR2x1_ASAP7_75t_SL g452 ( .A(n_403), .B(n_416), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_401), .B(n_424), .C(n_423), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g454 ( .A1(n_426), .A2(n_436), .B(n_415), .C(n_431), .Y(n_454) );
OAI211xp5_ASAP7_75t_L g455 ( .A1(n_409), .A2(n_431), .B(n_433), .C(n_434), .Y(n_455) );
AOI221x1_ASAP7_75t_L g456 ( .A1(n_453), .A2(n_426), .B1(n_425), .B2(n_422), .C(n_418), .Y(n_456) );
OAI211xp5_ASAP7_75t_SL g457 ( .A1(n_447), .A2(n_429), .B(n_435), .C(n_419), .Y(n_457) );
OAI211xp5_ASAP7_75t_SL g458 ( .A1(n_454), .A2(n_430), .B(n_410), .C(n_421), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_451), .B(n_414), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_452), .A2(n_420), .B(n_432), .Y(n_460) );
AO22x2_ASAP7_75t_L g461 ( .A1(n_451), .A2(n_413), .B1(n_428), .B2(n_427), .Y(n_461) );
OAI31xp33_ASAP7_75t_L g462 ( .A1(n_448), .A2(n_412), .A3(n_442), .B(n_408), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_450), .B(n_444), .Y(n_463) );
XNOR2xp5_ASAP7_75t_L g464 ( .A(n_460), .B(n_455), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_459), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_461), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_461), .Y(n_467) );
NAND4xp75_ASAP7_75t_L g468 ( .A(n_466), .B(n_462), .C(n_456), .D(n_463), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_465), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_464), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_469), .Y(n_471) );
NOR3xp33_ASAP7_75t_SL g472 ( .A(n_468), .B(n_464), .C(n_467), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_471), .Y(n_473) );
INVx2_ASAP7_75t_SL g474 ( .A(n_473), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_474), .A2(n_470), .B1(n_458), .B2(n_457), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_475), .A2(n_472), .B(n_449), .Y(n_476) );
endmodule