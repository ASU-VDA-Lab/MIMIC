module fake_jpeg_14247_n_217 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_217);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx5_ASAP7_75t_SL g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_5),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_52),
.Y(n_77)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_24),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

CKINVDCx9p33_ASAP7_75t_R g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_33),
.Y(n_91)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_63),
.Y(n_74)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_62),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

AND2x4_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_25),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_0),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_73),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_35),
.B1(n_27),
.B2(n_28),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_87),
.B1(n_63),
.B2(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_38),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_31),
.B1(n_27),
.B2(n_35),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_76),
.A2(n_85),
.B1(n_55),
.B2(n_58),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_28),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_26),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_60),
.B1(n_47),
.B2(n_26),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_18),
.B1(n_36),
.B2(n_33),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_37),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_29),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_92),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_116),
.B1(n_102),
.B2(n_66),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_67),
.A2(n_36),
.B1(n_29),
.B2(n_17),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_99),
.A2(n_110),
.B1(n_72),
.B2(n_64),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_104),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_107),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_77),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

BUFx2_ASAP7_75t_SL g134 ( 
.A(n_105),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_68),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_111),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_67),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_74),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_115),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_71),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_118),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_2),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_114),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

AOI22x1_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_86),
.B1(n_66),
.B2(n_64),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_79),
.B(n_118),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_86),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_70),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_106),
.B(n_107),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_140),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_113),
.B1(n_103),
.B2(n_117),
.Y(n_146)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_93),
.B(n_83),
.CI(n_3),
.CON(n_137),
.SN(n_137)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_83),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_139),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_7),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_120),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_143),
.B(n_148),
.Y(n_165)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_146),
.A2(n_154),
.B1(n_157),
.B2(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_103),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_102),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_153),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_133),
.B1(n_127),
.B2(n_137),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_152),
.B(n_156),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_132),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_134),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_131),
.A2(n_97),
.B1(n_92),
.B2(n_79),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_70),
.B1(n_82),
.B2(n_101),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_158),
.A2(n_128),
.B1(n_141),
.B2(n_142),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_133),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_9),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_10),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_169),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_164),
.A2(n_168),
.B1(n_175),
.B2(n_125),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_123),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_162),
.Y(n_188)
);

AOI22x1_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_127),
.B1(n_137),
.B2(n_128),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_147),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_160),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_153),
.B1(n_145),
.B2(n_154),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_176),
.B(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_181),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_159),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_186),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_152),
.B(n_145),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_169),
.A2(n_158),
.B1(n_149),
.B2(n_157),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_182),
.A2(n_175),
.B1(n_162),
.B2(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_185),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_172),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_184),
.B(n_188),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_165),
.B(n_125),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_135),
.C(n_126),
.Y(n_186)
);

OAI211xp5_ASAP7_75t_L g196 ( 
.A1(n_187),
.A2(n_166),
.B(n_168),
.C(n_170),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_126),
.C(n_136),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_172),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_194),
.A2(n_187),
.B1(n_188),
.B2(n_181),
.Y(n_202)
);

NAND4xp25_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_182),
.C(n_171),
.D(n_15),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_179),
.Y(n_200)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_189),
.Y(n_199)
);

OAI21x1_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_204),
.B(n_205),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_201),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_192),
.B(n_180),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_202),
.A2(n_197),
.B1(n_194),
.B2(n_198),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_191),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_180),
.C(n_168),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_205),
.A2(n_193),
.B1(n_190),
.B2(n_195),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_210),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_207),
.A2(n_204),
.B(n_200),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_212),
.A2(n_213),
.B(n_211),
.Y(n_214)
);

AOI31xp33_ASAP7_75t_L g213 ( 
.A1(n_206),
.A2(n_209),
.A3(n_171),
.B(n_210),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_215),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g217 ( 
.A(n_216),
.Y(n_217)
);


endmodule