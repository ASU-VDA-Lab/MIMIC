module real_aes_6876_n_271 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_271);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_271;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_769;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_0), .A2(n_74), .B1(n_407), .B2(n_576), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_1), .A2(n_40), .B1(n_389), .B2(n_390), .Y(n_759) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_2), .A2(n_204), .B1(n_479), .B2(n_480), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_3), .Y(n_742) );
AOI22xp33_ASAP7_75t_SL g758 ( .A1(n_4), .A2(n_264), .B1(n_553), .B2(n_554), .Y(n_758) );
AOI22xp33_ASAP7_75t_SL g574 ( .A1(n_5), .A2(n_98), .B1(n_327), .B2(n_486), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_6), .A2(n_122), .B1(n_389), .B2(n_666), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_7), .A2(n_134), .B1(n_403), .B2(n_615), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_8), .A2(n_101), .B1(n_375), .B2(n_378), .Y(n_435) );
AOI22xp33_ASAP7_75t_SL g446 ( .A1(n_9), .A2(n_228), .B1(n_385), .B2(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g428 ( .A(n_10), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_11), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_12), .A2(n_224), .B1(n_407), .B2(n_409), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_13), .A2(n_127), .B1(n_725), .B2(n_726), .C(n_727), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_14), .A2(n_34), .B1(n_390), .B2(n_482), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_15), .A2(n_141), .B1(n_369), .B2(n_430), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_16), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_17), .A2(n_152), .B1(n_352), .B2(n_359), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_18), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_19), .B(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_20), .A2(n_135), .B1(n_414), .B2(n_567), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_21), .A2(n_263), .B1(n_399), .B2(n_400), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_22), .A2(n_131), .B1(n_516), .B2(n_517), .Y(n_515) );
AO22x2_ASAP7_75t_L g305 ( .A1(n_23), .A2(n_91), .B1(n_297), .B2(n_302), .Y(n_305) );
INVx1_ASAP7_75t_L g842 ( .A(n_23), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_24), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_25), .A2(n_46), .B1(n_615), .B2(n_767), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_26), .A2(n_242), .B1(n_389), .B2(n_390), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_27), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_28), .Y(n_781) );
AOI22xp33_ASAP7_75t_SL g438 ( .A1(n_29), .A2(n_212), .B1(n_439), .B2(n_441), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g849 ( .A(n_30), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_31), .A2(n_236), .B1(n_444), .B2(n_599), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_32), .A2(n_257), .B1(n_486), .B2(n_664), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_33), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_35), .A2(n_136), .B1(n_556), .B2(n_558), .Y(n_555) );
AOI22xp33_ASAP7_75t_SL g578 ( .A1(n_36), .A2(n_42), .B1(n_314), .B2(n_340), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_37), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_38), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_39), .A2(n_164), .B1(n_335), .B2(n_580), .Y(n_579) );
AO22x2_ASAP7_75t_L g307 ( .A1(n_41), .A2(n_94), .B1(n_297), .B2(n_298), .Y(n_307) );
INVx1_ASAP7_75t_L g843 ( .A(n_41), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_43), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_44), .Y(n_350) );
AOI22xp33_ASAP7_75t_SL g433 ( .A1(n_45), .A2(n_219), .B1(n_399), .B2(n_434), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_47), .Y(n_670) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_48), .A2(n_192), .B1(n_404), .B2(n_407), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_49), .B(n_397), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_50), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_51), .A2(n_209), .B1(n_340), .B2(n_485), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_52), .A2(n_210), .B1(n_558), .B2(n_661), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_53), .A2(n_89), .B1(n_329), .B2(n_404), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_54), .A2(n_95), .B1(n_475), .B2(n_476), .Y(n_777) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_55), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_56), .A2(n_107), .B1(n_292), .B2(n_526), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_57), .A2(n_156), .B1(n_365), .B2(n_594), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_58), .A2(n_77), .B1(n_580), .B2(n_870), .Y(n_869) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_59), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_60), .A2(n_230), .B1(n_415), .B2(n_461), .Y(n_540) );
AOI22xp33_ASAP7_75t_SL g552 ( .A1(n_61), .A2(n_234), .B1(n_553), .B2(n_554), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_62), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_63), .A2(n_176), .B1(n_354), .B2(n_400), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_64), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g851 ( .A(n_65), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_66), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_67), .A2(n_118), .B1(n_464), .B2(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_68), .Y(n_630) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_69), .A2(n_125), .B1(n_484), .B2(n_485), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_70), .A2(n_130), .B1(n_329), .B2(n_444), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_71), .A2(n_137), .B1(n_414), .B2(n_505), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_72), .Y(n_332) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_73), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_75), .A2(n_199), .B1(n_519), .B2(n_521), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_76), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_78), .Y(n_675) );
AOI222xp33_ASAP7_75t_L g410 ( .A1(n_79), .A2(n_161), .B1(n_172), .B2(n_411), .C1(n_413), .C2(n_415), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_80), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_81), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g822 ( .A(n_82), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_83), .A2(n_115), .B1(n_597), .B2(n_866), .Y(n_865) );
AOI22xp33_ASAP7_75t_SL g459 ( .A1(n_84), .A2(n_222), .B1(n_460), .B2(n_461), .Y(n_459) );
AOI222xp33_ASAP7_75t_L g600 ( .A1(n_85), .A2(n_93), .B1(n_124), .B2(n_348), .C1(n_371), .C2(n_601), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_86), .A2(n_188), .B1(n_407), .B2(n_666), .Y(n_756) );
AOI22xp33_ASAP7_75t_SL g465 ( .A1(n_87), .A2(n_142), .B1(n_466), .B2(n_467), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_88), .A2(n_154), .B1(n_367), .B2(n_371), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_90), .A2(n_155), .B1(n_772), .B2(n_775), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_92), .Y(n_508) );
INVx1_ASAP7_75t_L g279 ( .A(n_96), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_97), .A2(n_191), .B1(n_313), .B2(n_320), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_99), .A2(n_267), .B1(n_556), .B2(n_769), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_100), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_102), .A2(n_268), .B1(n_556), .B2(n_580), .Y(n_590) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_103), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_104), .A2(n_611), .B1(n_644), .B2(n_645), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_104), .Y(n_644) );
INVx1_ASAP7_75t_L g277 ( .A(n_105), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_106), .A2(n_175), .B1(n_403), .B2(n_404), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_108), .A2(n_114), .B1(n_389), .B2(n_390), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g338 ( .A(n_109), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_110), .A2(n_189), .B1(n_291), .B2(n_308), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_111), .A2(n_243), .B1(n_375), .B2(n_378), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_112), .A2(n_238), .B1(n_658), .B2(n_659), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_113), .A2(n_261), .B1(n_361), .B2(n_567), .Y(n_748) );
AOI22xp33_ASAP7_75t_SL g689 ( .A1(n_116), .A2(n_120), .B1(n_400), .B2(n_567), .Y(n_689) );
OA22x2_ASAP7_75t_L g677 ( .A1(n_117), .A2(n_678), .B1(n_679), .B2(n_697), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_117), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_119), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_121), .B(n_688), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_123), .A2(n_128), .B1(n_385), .B2(n_386), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_126), .Y(n_783) );
AOI22xp5_ASAP7_75t_SL g422 ( .A1(n_129), .A2(n_423), .B1(n_424), .B2(n_449), .Y(n_422) );
INVx1_ASAP7_75t_L g449 ( .A(n_129), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_132), .A2(n_139), .B1(n_375), .B2(n_378), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_133), .A2(n_162), .B1(n_517), .B2(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_138), .A2(n_173), .B1(n_308), .B2(n_444), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g643 ( .A(n_140), .Y(n_643) );
XNOR2x2_ASAP7_75t_L g286 ( .A(n_143), .B(n_287), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_144), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_145), .B(n_466), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_146), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_147), .Y(n_712) );
INVx2_ASAP7_75t_L g280 ( .A(n_148), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_149), .A2(n_165), .B1(n_479), .B2(n_864), .Y(n_863) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_150), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_151), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_153), .B(n_686), .Y(n_685) );
AOI222xp33_ASAP7_75t_L g730 ( .A1(n_157), .A2(n_218), .B1(n_250), .B2(n_352), .C1(n_411), .C2(n_731), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_158), .Y(n_790) );
AND2x6_ASAP7_75t_L g276 ( .A(n_159), .B(n_277), .Y(n_276) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_159), .Y(n_836) );
AO22x2_ASAP7_75t_L g296 ( .A1(n_160), .A2(n_223), .B1(n_297), .B2(n_298), .Y(n_296) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_163), .A2(n_227), .B1(n_409), .B2(n_471), .Y(n_470) );
AOI22xp33_ASAP7_75t_SL g364 ( .A1(n_166), .A2(n_239), .B1(n_365), .B2(n_369), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_167), .B(n_378), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_168), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_169), .Y(n_854) );
INVx1_ASAP7_75t_L g860 ( .A(n_170), .Y(n_860) );
AOI22xp33_ASAP7_75t_SL g473 ( .A1(n_171), .A2(n_260), .B1(n_474), .B2(n_476), .Y(n_473) );
AOI22xp33_ASAP7_75t_SL g463 ( .A1(n_174), .A2(n_226), .B1(n_372), .B2(n_464), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_177), .A2(n_186), .B1(n_367), .B2(n_460), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_178), .Y(n_325) );
AOI22xp33_ASAP7_75t_SL g696 ( .A1(n_179), .A2(n_255), .B1(n_335), .B2(n_666), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_180), .A2(n_205), .B1(n_340), .B2(n_447), .Y(n_816) );
AOI22xp33_ASAP7_75t_SL g695 ( .A1(n_181), .A2(n_246), .B1(n_516), .B2(n_659), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_182), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_183), .A2(n_270), .B1(n_517), .B2(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_184), .A2(n_216), .B1(n_320), .B2(n_617), .Y(n_616) );
AO22x2_ASAP7_75t_L g301 ( .A1(n_185), .A2(n_244), .B1(n_297), .B2(n_302), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_187), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_190), .B(n_731), .Y(n_855) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_193), .A2(n_225), .B1(n_314), .B2(n_580), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_194), .A2(n_206), .B1(n_313), .B2(n_385), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g622 ( .A(n_195), .Y(n_622) );
AOI22xp33_ASAP7_75t_SL g683 ( .A1(n_196), .A2(n_245), .B1(n_414), .B2(n_460), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_197), .A2(n_249), .B1(n_523), .B2(n_524), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_198), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_200), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_201), .Y(n_808) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_202), .A2(n_221), .B1(n_414), .B2(n_567), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_203), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_207), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_208), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_211), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_213), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_214), .B(n_397), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_215), .A2(n_702), .B1(n_732), .B2(n_733), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_215), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_217), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_220), .B(n_359), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_223), .B(n_841), .Y(n_840) );
OA22x2_ASAP7_75t_L g453 ( .A1(n_229), .A2(n_454), .B1(n_455), .B2(n_487), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_229), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_231), .Y(n_636) );
INVx1_ASAP7_75t_L g654 ( .A(n_232), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_233), .Y(n_709) );
INVx1_ASAP7_75t_L g760 ( .A(n_235), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_237), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_240), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_241), .A2(n_846), .B1(n_871), .B2(n_872), .Y(n_845) );
INVx1_ASAP7_75t_L g871 ( .A(n_241), .Y(n_871) );
INVx1_ASAP7_75t_L g839 ( .A(n_244), .Y(n_839) );
XNOR2x2_ASAP7_75t_L g586 ( .A(n_247), .B(n_587), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_248), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_251), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_252), .Y(n_819) );
INVx1_ASAP7_75t_L g882 ( .A(n_253), .Y(n_882) );
OA22x2_ASAP7_75t_SL g883 ( .A1(n_253), .A2(n_846), .B1(n_872), .B2(n_882), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_254), .A2(n_763), .B1(n_791), .B2(n_792), .Y(n_762) );
INVx1_ASAP7_75t_L g791 ( .A(n_254), .Y(n_791) );
INVx1_ASAP7_75t_L g297 ( .A(n_256), .Y(n_297) );
INVx1_ASAP7_75t_L g299 ( .A(n_256), .Y(n_299) );
AOI211xp5_ASAP7_75t_L g271 ( .A1(n_258), .A2(n_272), .B(n_281), .C(n_844), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_259), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_262), .Y(n_813) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_265), .Y(n_785) );
OA22x2_ASAP7_75t_L g795 ( .A1(n_266), .A2(n_796), .B1(n_797), .B2(n_798), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_266), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_269), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_273), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_277), .Y(n_835) );
OAI21xp5_ASAP7_75t_L g880 ( .A1(n_278), .A2(n_834), .B(n_881), .Y(n_880) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_606), .B1(n_829), .B2(n_830), .C(n_831), .Y(n_281) );
INVx1_ASAP7_75t_L g829 ( .A(n_282), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B1(n_418), .B2(n_605), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_286), .B1(n_380), .B2(n_417), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_288), .B(n_345), .Y(n_287) );
NOR3xp33_ASAP7_75t_L g288 ( .A(n_289), .B(n_324), .C(n_337), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_312), .Y(n_289) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx3_ASAP7_75t_L g479 ( .A(n_292), .Y(n_479) );
BUFx3_ASAP7_75t_L g615 ( .A(n_292), .Y(n_615) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g408 ( .A(n_293), .Y(n_408) );
BUFx2_ASAP7_75t_SL g444 ( .A(n_293), .Y(n_444) );
BUFx2_ASAP7_75t_SL g821 ( .A(n_293), .Y(n_821) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_303), .Y(n_293) );
AND2x6_ASAP7_75t_L g329 ( .A(n_294), .B(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g340 ( .A(n_294), .B(n_319), .Y(n_340) );
AND2x6_ASAP7_75t_L g348 ( .A(n_294), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_300), .Y(n_294) );
AND2x2_ASAP7_75t_L g336 ( .A(n_295), .B(n_301), .Y(n_336) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_296), .B(n_301), .Y(n_311) );
AND2x2_ASAP7_75t_L g317 ( .A(n_296), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g358 ( .A(n_296), .B(n_305), .Y(n_358) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g302 ( .A(n_299), .Y(n_302) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g318 ( .A(n_301), .Y(n_318) );
INVx1_ASAP7_75t_L g357 ( .A(n_301), .Y(n_357) );
AND2x4_ASAP7_75t_L g309 ( .A(n_303), .B(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g335 ( .A(n_303), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_303), .B(n_317), .Y(n_344) );
AND2x2_ASAP7_75t_L g405 ( .A(n_303), .B(n_317), .Y(n_405) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
AND2x2_ASAP7_75t_L g319 ( .A(n_304), .B(n_307), .Y(n_319) );
OR2x2_ASAP7_75t_L g331 ( .A(n_304), .B(n_307), .Y(n_331) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g349 ( .A(n_305), .B(n_307), .Y(n_349) );
AND2x2_ASAP7_75t_L g356 ( .A(n_306), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g559 ( .A(n_306), .Y(n_559) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g323 ( .A(n_307), .Y(n_323) );
BUFx2_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
BUFx3_ASAP7_75t_L g409 ( .A(n_309), .Y(n_409) );
BUFx3_ASAP7_75t_L g526 ( .A(n_309), .Y(n_526) );
BUFx3_ASAP7_75t_L g576 ( .A(n_309), .Y(n_576) );
BUFx2_ASAP7_75t_SL g599 ( .A(n_309), .Y(n_599) );
BUFx2_ASAP7_75t_L g666 ( .A(n_309), .Y(n_666) );
BUFx3_ASAP7_75t_L g866 ( .A(n_309), .Y(n_866) );
AND2x2_ASAP7_75t_L g558 ( .A(n_310), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x6_ASAP7_75t_L g322 ( .A(n_311), .B(n_323), .Y(n_322) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g520 ( .A(n_314), .Y(n_520) );
INVx4_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx3_ASAP7_75t_L g387 ( .A(n_315), .Y(n_387) );
INVx1_ASAP7_75t_L g447 ( .A(n_315), .Y(n_447) );
INVx2_ASAP7_75t_L g475 ( .A(n_315), .Y(n_475) );
INVx3_ASAP7_75t_L g554 ( .A(n_315), .Y(n_554) );
INVx5_ASAP7_75t_L g661 ( .A(n_315), .Y(n_661) );
INVx8_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_317), .B(n_319), .Y(n_711) );
INVx1_ASAP7_75t_L g373 ( .A(n_318), .Y(n_373) );
AND2x6_ASAP7_75t_L g379 ( .A(n_319), .B(n_336), .Y(n_379) );
NAND2x1p5_ASAP7_75t_L g395 ( .A(n_319), .B(n_336), .Y(n_395) );
BUFx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g390 ( .A(n_321), .Y(n_390) );
BUFx2_ASAP7_75t_L g476 ( .A(n_321), .Y(n_476) );
BUFx2_ASAP7_75t_L g521 ( .A(n_321), .Y(n_521) );
INVx6_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g580 ( .A(n_322), .Y(n_580) );
INVx1_ASAP7_75t_L g368 ( .A(n_323), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B1(n_332), .B2(n_333), .Y(n_324) );
INVx2_ASAP7_75t_L g767 ( .A(n_326), .Y(n_767) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_327), .Y(n_722) );
INVx5_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g403 ( .A(n_328), .Y(n_403) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_328), .Y(n_472) );
INVx4_ASAP7_75t_L g549 ( .A(n_328), .Y(n_549) );
INVx11_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx11_ASAP7_75t_L g440 ( .A(n_329), .Y(n_440) );
AND2x4_ASAP7_75t_L g377 ( .A(n_330), .B(n_336), .Y(n_377) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g498 ( .A(n_331), .B(n_499), .Y(n_498) );
INVx4_ASAP7_75t_L g523 ( .A(n_333), .Y(n_523) );
INVx4_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx3_ASAP7_75t_L g389 ( .A(n_335), .Y(n_389) );
BUFx3_ASAP7_75t_L g482 ( .A(n_335), .Y(n_482) );
INVx2_ASAP7_75t_L g557 ( .A(n_335), .Y(n_557) );
INVx1_ASAP7_75t_L g499 ( .A(n_336), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_339), .B1(n_341), .B2(n_342), .Y(n_337) );
INVx2_ASAP7_75t_L g385 ( .A(n_339), .Y(n_385) );
INVx3_ASAP7_75t_L g516 ( .A(n_339), .Y(n_516) );
INVx2_ASAP7_75t_L g553 ( .A(n_339), .Y(n_553) );
INVx2_ASAP7_75t_L g621 ( .A(n_339), .Y(n_621) );
INVx6_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx3_ASAP7_75t_L g484 ( .A(n_340), .Y(n_484) );
BUFx3_ASAP7_75t_L g664 ( .A(n_340), .Y(n_664) );
BUFx3_ASAP7_75t_L g774 ( .A(n_340), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_342), .A2(n_825), .B1(n_826), .B2(n_827), .Y(n_824) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g623 ( .A(n_343), .Y(n_623) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_363), .Y(n_345) );
OAI21xp5_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_350), .B(n_351), .Y(n_346) );
OAI21xp5_ASAP7_75t_SL g457 ( .A1(n_347), .A2(n_458), .B(n_459), .Y(n_457) );
OAI21xp5_ASAP7_75t_SL g564 ( .A1(n_347), .A2(n_565), .B(n_566), .Y(n_564) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx4_ASAP7_75t_L g412 ( .A(n_348), .Y(n_412) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_348), .Y(n_539) );
BUFx3_ASAP7_75t_L g674 ( .A(n_348), .Y(n_674) );
AND2x4_ASAP7_75t_L g372 ( .A(n_349), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g511 ( .A(n_349), .Y(n_511) );
INVx3_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx4_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g784 ( .A(n_354), .Y(n_784) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_355), .Y(n_399) );
BUFx4f_ASAP7_75t_SL g460 ( .A(n_355), .Y(n_460) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_355), .Y(n_505) );
AND2x4_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
INVx1_ASAP7_75t_L g362 ( .A(n_357), .Y(n_362) );
AND2x4_ASAP7_75t_L g361 ( .A(n_358), .B(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g367 ( .A(n_358), .B(n_368), .Y(n_367) );
NAND2x1p5_ASAP7_75t_L g631 ( .A(n_358), .B(n_559), .Y(n_631) );
BUFx4f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx12f_ASAP7_75t_L g414 ( .A(n_361), .Y(n_414) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_361), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_374), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx3_ASAP7_75t_L g400 ( .A(n_367), .Y(n_400) );
BUFx2_ASAP7_75t_L g434 ( .A(n_367), .Y(n_434) );
BUFx2_ASAP7_75t_L g464 ( .A(n_367), .Y(n_464) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx2_ASAP7_75t_SL g415 ( .A(n_372), .Y(n_415) );
BUFx2_ASAP7_75t_SL g567 ( .A(n_372), .Y(n_567) );
INVx1_ASAP7_75t_L g512 ( .A(n_373), .Y(n_512) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g397 ( .A(n_376), .Y(n_397) );
INVx2_ASAP7_75t_L g466 ( .A(n_376), .Y(n_466) );
INVx5_ASAP7_75t_L g688 ( .A(n_376), .Y(n_688) );
INVx4_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g468 ( .A(n_379), .Y(n_468) );
BUFx4f_ASAP7_75t_L g544 ( .A(n_379), .Y(n_544) );
BUFx2_ASAP7_75t_L g726 ( .A(n_379), .Y(n_726) );
INVx1_ASAP7_75t_L g417 ( .A(n_380), .Y(n_417) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
XOR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_416), .Y(n_381) );
NAND4xp75_ASAP7_75t_L g382 ( .A(n_383), .B(n_391), .C(n_401), .D(n_410), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_388), .Y(n_383) );
INVx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OA211x2_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B(n_396), .C(n_398), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_393), .A2(n_497), .B1(n_780), .B2(n_781), .Y(n_779) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g501 ( .A(n_394), .Y(n_501) );
INVx1_ASAP7_75t_L g745 ( .A(n_394), .Y(n_745) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx3_ASAP7_75t_L g669 ( .A(n_395), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_399), .Y(n_812) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_406), .Y(n_401) );
INVx2_ASAP7_75t_L g825 ( .A(n_403), .Y(n_825) );
BUFx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx3_ASAP7_75t_L g442 ( .A(n_405), .Y(n_442) );
BUFx3_ASAP7_75t_L g486 ( .A(n_405), .Y(n_486) );
BUFx3_ASAP7_75t_L g517 ( .A(n_405), .Y(n_517) );
INVx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx3_ASAP7_75t_L g658 ( .A(n_408), .Y(n_658) );
INVxp67_ASAP7_75t_L g627 ( .A(n_409), .Y(n_627) );
INVx2_ASAP7_75t_L g427 ( .A(n_411), .Y(n_427) );
INVx4_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI21xp5_ASAP7_75t_SL g746 ( .A1(n_412), .A2(n_747), .B(n_748), .Y(n_746) );
BUFx4f_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g431 ( .A(n_414), .Y(n_431) );
INVx1_ASAP7_75t_L g605 ( .A(n_418), .Y(n_605) );
XNOR2xp5_ASAP7_75t_SL g418 ( .A(n_419), .B(n_450), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_425), .B(n_436), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_432), .Y(n_425) );
OAI21xp5_ASAP7_75t_SL g426 ( .A1(n_427), .A2(n_428), .B(n_429), .Y(n_426) );
OAI21xp33_ASAP7_75t_SL g502 ( .A1(n_427), .A2(n_503), .B(n_504), .Y(n_502) );
OAI221xp5_ASAP7_75t_L g635 ( .A1(n_427), .A2(n_636), .B1(n_637), .B2(n_638), .C(n_639), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g782 ( .A1(n_427), .A2(n_783), .B1(n_784), .B2(n_785), .C(n_786), .Y(n_782) );
OAI221xp5_ASAP7_75t_L g852 ( .A1(n_427), .A2(n_784), .B1(n_853), .B2(n_854), .C(n_855), .Y(n_852) );
INVx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_435), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_445), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_443), .Y(n_437) );
INVx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx4_ASAP7_75t_L g597 ( .A(n_440), .Y(n_597) );
INVx4_ASAP7_75t_L g659 ( .A(n_440), .Y(n_659) );
BUFx4f_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_447), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_529), .B1(n_603), .B2(n_604), .Y(n_450) );
INVx1_ASAP7_75t_L g603 ( .A(n_451), .Y(n_603) );
OAI22xp5_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_453), .B1(n_488), .B2(n_528), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_SL g487 ( .A(n_455), .Y(n_487) );
NAND3x1_ASAP7_75t_L g455 ( .A(n_456), .B(n_469), .C(n_477), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_462), .Y(n_456) );
INVx2_ASAP7_75t_L g507 ( .A(n_461), .Y(n_507) );
BUFx2_ASAP7_75t_L g640 ( .A(n_461), .Y(n_640) );
BUFx3_ASAP7_75t_L g731 ( .A(n_461), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_465), .Y(n_462) );
INVx1_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_SL g686 ( .A(n_468), .Y(n_686) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_473), .Y(n_469) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVxp67_ASAP7_75t_L g713 ( .A(n_476), .Y(n_713) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_483), .Y(n_477) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_481), .A2(n_625), .B1(n_626), .B2(n_627), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_481), .A2(n_720), .B1(n_721), .B2(n_723), .Y(n_719) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_L g864 ( .A(n_482), .Y(n_864) );
BUFx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g528 ( .A(n_488), .Y(n_528) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
XNOR2x1_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_514), .Y(n_491) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_502), .C(n_506), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_500), .B2(n_501), .Y(n_493) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_497), .A2(n_501), .B1(n_642), .B2(n_643), .Y(n_641) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g667 ( .A1(n_498), .A2(n_668), .B1(n_669), .B2(n_670), .C(n_671), .Y(n_667) );
BUFx3_ASAP7_75t_L g743 ( .A(n_498), .Y(n_743) );
INVx2_ASAP7_75t_L g802 ( .A(n_498), .Y(n_802) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_505), .Y(n_594) );
OAI22xp5_ASAP7_75t_SL g506 ( .A1(n_507), .A2(n_508), .B1(n_509), .B2(n_513), .Y(n_506) );
INVx1_ASAP7_75t_L g601 ( .A(n_507), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_509), .A2(n_788), .B1(n_789), .B2(n_790), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_509), .A2(n_857), .B1(n_858), .B2(n_860), .Y(n_856) );
BUFx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
CKINVDCx16_ASAP7_75t_R g634 ( .A(n_510), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_510), .A2(n_631), .B1(n_728), .B2(n_729), .Y(n_727) );
OR2x6_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
AND4x1_ASAP7_75t_L g514 ( .A(n_515), .B(n_518), .C(n_522), .D(n_527), .Y(n_514) );
INVx1_ASAP7_75t_L g776 ( .A(n_517), .Y(n_776) );
INVx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_525), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_704) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g604 ( .A(n_529), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B1(n_583), .B2(n_584), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OAI22x1_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B1(n_561), .B2(n_582), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_532), .A2(n_533), .B1(n_586), .B2(n_602), .Y(n_585) );
INVx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
XOR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_560), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_535), .B(n_546), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_541), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_538), .B(n_540), .Y(n_536) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .C(n_545), .Y(n_541) );
NOR2x1_ASAP7_75t_L g546 ( .A(n_547), .B(n_551), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
INVxp67_ASAP7_75t_L g717 ( .A(n_553), .Y(n_717) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx3_ASAP7_75t_L g582 ( .A(n_561), .Y(n_582) );
XOR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_581), .Y(n_561) );
NAND2x1_ASAP7_75t_SL g562 ( .A(n_563), .B(n_572), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_568), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .C(n_571), .Y(n_568) );
NOR2x1_ASAP7_75t_L g572 ( .A(n_573), .B(n_577), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
BUFx2_ASAP7_75t_L g769 ( .A(n_576), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g602 ( .A(n_586), .Y(n_602) );
NAND4xp75_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .C(n_595), .D(n_600), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
AND2x2_ASAP7_75t_SL g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx2_ASAP7_75t_SL g637 ( .A(n_594), .Y(n_637) );
INVx2_ASAP7_75t_SL g751 ( .A(n_594), .Y(n_751) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
INVx1_ASAP7_75t_SL g823 ( .A(n_599), .Y(n_823) );
INVx1_ASAP7_75t_L g830 ( .A(n_606), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B1(n_646), .B2(n_647), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g645 ( .A(n_611), .Y(n_645) );
AND2x2_ASAP7_75t_SL g611 ( .A(n_612), .B(n_628), .Y(n_611) );
NOR3xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_618), .C(n_624), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B1(n_622), .B2(n_623), .Y(n_618) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_623), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_715) );
NOR3xp33_ASAP7_75t_SL g628 ( .A(n_629), .B(n_635), .C(n_641), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B1(n_632), .B2(n_633), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_631), .A2(n_750), .B1(n_751), .B2(n_752), .Y(n_749) );
BUFx3_ASAP7_75t_L g789 ( .A(n_631), .Y(n_789) );
INVx4_ASAP7_75t_L g859 ( .A(n_631), .Y(n_859) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
XNOR2xp5_ASAP7_75t_SL g647 ( .A(n_648), .B(n_734), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI22xp5_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_652), .B1(n_700), .B2(n_701), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_677), .B1(n_698), .B2(n_699), .Y(n_652) );
INVx2_ASAP7_75t_SL g698 ( .A(n_653), .Y(n_698) );
XNOR2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
NOR4xp75_ASAP7_75t_L g655 ( .A(n_656), .B(n_662), .C(n_667), .D(n_672), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_657), .B(n_660), .Y(n_656) );
INVxp67_ASAP7_75t_L g706 ( .A(n_658), .Y(n_706) );
BUFx6f_ASAP7_75t_L g870 ( .A(n_661), .Y(n_870) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_663), .B(n_665), .Y(n_662) );
INVx2_ASAP7_75t_L g805 ( .A(n_669), .Y(n_805) );
OAI21xp5_ASAP7_75t_SL g672 ( .A1(n_673), .A2(n_675), .B(n_676), .Y(n_672) );
OAI21xp5_ASAP7_75t_SL g681 ( .A1(n_673), .A2(n_682), .B(n_683), .Y(n_681) );
OAI21xp33_ASAP7_75t_L g807 ( .A1(n_673), .A2(n_808), .B(n_809), .Y(n_807) );
INVx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g699 ( .A(n_677), .Y(n_699) );
INVx1_ASAP7_75t_L g697 ( .A(n_679), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_690), .Y(n_679) );
NOR2xp67_ASAP7_75t_L g680 ( .A(n_681), .B(n_684), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .C(n_689), .Y(n_684) );
BUFx6f_ASAP7_75t_L g725 ( .A(n_688), .Y(n_725) );
NOR2x1_ASAP7_75t_L g690 ( .A(n_691), .B(n_694), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g733 ( .A(n_702), .Y(n_733) );
AND4x1_ASAP7_75t_L g702 ( .A(n_703), .B(n_714), .C(n_724), .D(n_730), .Y(n_702) );
NOR2xp33_ASAP7_75t_SL g703 ( .A(n_704), .B(n_708), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_710), .B1(n_712), .B2(n_713), .Y(n_708) );
BUFx2_ASAP7_75t_R g710 ( .A(n_711), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_719), .Y(n_714) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B1(n_793), .B2(n_794), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OAI22xp5_ASAP7_75t_SL g736 ( .A1(n_737), .A2(n_738), .B1(n_761), .B2(n_762), .Y(n_736) );
OAI22xp5_ASAP7_75t_SL g794 ( .A1(n_737), .A2(n_738), .B1(n_795), .B2(n_828), .Y(n_794) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
XOR2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_760), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_753), .Y(n_739) );
NOR3xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_746), .C(n_749), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_757), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g792 ( .A(n_763), .Y(n_792) );
AND2x2_ASAP7_75t_SL g763 ( .A(n_764), .B(n_778), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_765), .B(n_770), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_768), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_777), .Y(n_770) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx3_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NOR3xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_782), .C(n_787), .Y(n_778) );
OAI22xp33_ASAP7_75t_L g810 ( .A1(n_789), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_810) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx2_ASAP7_75t_L g828 ( .A(n_795), .Y(n_828) );
INVx2_ASAP7_75t_SL g797 ( .A(n_798), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_799), .B(n_814), .Y(n_798) );
NOR3xp33_ASAP7_75t_L g799 ( .A(n_800), .B(n_807), .C(n_810), .Y(n_799) );
OAI22xp5_ASAP7_75t_SL g800 ( .A1(n_801), .A2(n_803), .B1(n_804), .B2(n_806), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g850 ( .A(n_802), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_804), .A2(n_849), .B1(n_850), .B2(n_851), .Y(n_848) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NOR3xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_818), .C(n_824), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_820), .B1(n_822), .B2(n_823), .Y(n_818) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_SL g831 ( .A(n_832), .Y(n_831) );
NOR2x1_ASAP7_75t_L g832 ( .A(n_833), .B(n_837), .Y(n_832) );
OR2x2_ASAP7_75t_SL g886 ( .A(n_833), .B(n_838), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_834), .B(n_836), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g875 ( .A(n_834), .Y(n_875) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_835), .B(n_878), .Y(n_881) );
CKINVDCx16_ASAP7_75t_R g878 ( .A(n_836), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_838), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
OAI322xp33_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_873), .A3(n_876), .B1(n_879), .B2(n_882), .C1(n_883), .C2(n_884), .Y(n_844) );
INVx2_ASAP7_75t_L g872 ( .A(n_846), .Y(n_872) );
AND2x2_ASAP7_75t_SL g846 ( .A(n_847), .B(n_861), .Y(n_846) );
NOR3xp33_ASAP7_75t_L g847 ( .A(n_848), .B(n_852), .C(n_856), .Y(n_847) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_862), .B(n_867), .Y(n_861) );
NAND2xp5_ASAP7_75t_SL g862 ( .A(n_863), .B(n_865), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_869), .Y(n_867) );
HB1xp67_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
HB1xp67_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g879 ( .A(n_880), .Y(n_879) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_885), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_886), .Y(n_885) );
endmodule