module fake_jpeg_21638_n_153 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_22),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_26),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_6),
.B(n_32),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_24),
.B1(n_38),
.B2(n_34),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_61),
.B1(n_46),
.B2(n_70),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_77),
.Y(n_81)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_83),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_84),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_65),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_48),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_97),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_43),
.B(n_66),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_99),
.C(n_100),
.Y(n_115)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_60),
.B1(n_48),
.B2(n_64),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_91),
.B1(n_96),
.B2(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_43),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_98),
.B(n_101),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_66),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_85),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_47),
.B1(n_45),
.B2(n_4),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_99),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_112),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_114),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_45),
.A3(n_47),
.B1(n_68),
.B2(n_44),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_54),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_121),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_123),
.B1(n_13),
.B2(n_15),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_116),
.C(n_103),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_3),
.B(n_5),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_112),
.A2(n_63),
.B1(n_62),
.B2(n_51),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_53),
.B1(n_50),
.B2(n_5),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_125),
.B(n_129),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_58),
.B1(n_55),
.B2(n_59),
.Y(n_129)
);

AO21x1_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_2),
.B(n_3),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_135),
.C(n_128),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_124),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_134),
.B(n_138),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_127),
.B(n_10),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_122),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_137),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_143),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_144),
.A2(n_130),
.B(n_141),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_136),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_146),
.B(n_135),
.Y(n_147)
);

INVxp33_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_140),
.C(n_18),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g150 ( 
.A(n_149),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_16),
.C(n_21),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_23),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_25),
.Y(n_153)
);


endmodule