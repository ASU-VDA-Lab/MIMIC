module fake_jpeg_16918_n_363 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_363);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_363;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_55),
.Y(n_72)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_41),
.Y(n_86)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_9),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_20),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx9p33_ASAP7_75t_R g84 ( 
.A(n_59),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_60),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_19),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_63),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_64),
.B(n_65),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_39),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_20),
.C(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_39),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_75),
.B(n_76),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NOR2xp67_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_34),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_51),
.B1(n_34),
.B2(n_37),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g143 ( 
.A(n_87),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_38),
.B1(n_29),
.B2(n_46),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_88),
.A2(n_91),
.B1(n_92),
.B2(n_54),
.Y(n_144)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_42),
.B1(n_52),
.B2(n_46),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_90),
.A2(n_67),
.B1(n_55),
.B2(n_47),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_38),
.B1(n_50),
.B2(n_52),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_64),
.A2(n_50),
.B1(n_42),
.B2(n_55),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_95),
.Y(n_141)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_SL g101 ( 
.A1(n_63),
.A2(n_59),
.B(n_48),
.Y(n_101)
);

AOI32xp33_ASAP7_75t_L g147 ( 
.A1(n_101),
.A2(n_53),
.A3(n_59),
.B1(n_57),
.B2(n_48),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_28),
.B1(n_30),
.B2(n_35),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_106),
.B1(n_116),
.B2(n_118),
.Y(n_138)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

BUFx2_ASAP7_75t_SL g133 ( 
.A(n_104),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_105),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_35),
.B1(n_30),
.B2(n_28),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_70),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_114),
.Y(n_121)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_81),
.A2(n_28),
.B1(n_30),
.B2(n_35),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_73),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_63),
.B(n_86),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_137),
.B(n_147),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_75),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_95),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_21),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_81),
.B1(n_79),
.B2(n_61),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_131),
.B1(n_139),
.B2(n_97),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_81),
.B1(n_79),
.B2(n_61),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_72),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_99),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_135),
.A2(n_142),
.B1(n_144),
.B2(n_118),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_96),
.B(n_69),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g139 ( 
.A1(n_96),
.A2(n_72),
.A3(n_76),
.B1(n_77),
.B2(n_63),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_145),
.B(n_148),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_112),
.A2(n_47),
.B1(n_40),
.B2(n_36),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_54),
.B(n_67),
.C(n_82),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_96),
.A2(n_33),
.B(n_71),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_160),
.B1(n_123),
.B2(n_136),
.Y(n_178)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_100),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_138),
.A2(n_94),
.B1(n_71),
.B2(n_97),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_158),
.A2(n_161),
.B1(n_124),
.B2(n_33),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_159),
.A2(n_171),
.B(n_176),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_145),
.A2(n_118),
.B1(n_22),
.B2(n_26),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_144),
.A2(n_82),
.B1(n_107),
.B2(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_89),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_164),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_114),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_170),
.B(n_174),
.Y(n_186)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_167),
.B(n_169),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

FAx1_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_73),
.CI(n_68),
.CON(n_169),
.SN(n_169)
);

AO22x1_ASAP7_75t_L g170 ( 
.A1(n_131),
.A2(n_49),
.B1(n_93),
.B2(n_99),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_68),
.Y(n_171)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_111),
.Y(n_174)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_119),
.C(n_135),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_179),
.C(n_187),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_178),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_139),
.Y(n_179)
);

OAI22x1_ASAP7_75t_SL g181 ( 
.A1(n_163),
.A2(n_169),
.B1(n_159),
.B2(n_156),
.Y(n_181)
);

OAI22x1_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_58),
.B1(n_60),
.B2(n_146),
.Y(n_214)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_136),
.C(n_147),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_121),
.C(n_141),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_194),
.C(n_196),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_191),
.B(n_60),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_26),
.B(n_21),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_193),
.A2(n_176),
.B(n_37),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_124),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_68),
.C(n_117),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_163),
.A2(n_154),
.B1(n_158),
.B2(n_161),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_200),
.B1(n_201),
.B2(n_173),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_60),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_203),
.C(n_58),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_170),
.A2(n_126),
.B1(n_120),
.B2(n_49),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_170),
.A2(n_49),
.B1(n_134),
.B2(n_122),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_153),
.B(n_134),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_167),
.B(n_165),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_150),
.B(n_146),
.C(n_143),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_205),
.B(n_217),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_207),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_157),
.Y(n_208)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_230),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_181),
.A2(n_153),
.B1(n_175),
.B2(n_172),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_210),
.A2(n_202),
.B1(n_201),
.B2(n_200),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_175),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_212),
.B(n_215),
.Y(n_250)
);

NOR2x1_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_122),
.Y(n_213)
);

AO22x1_ASAP7_75t_L g253 ( 
.A1(n_213),
.A2(n_93),
.B1(n_104),
.B2(n_58),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_214),
.B(n_227),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_216),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_192),
.B(n_22),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_218),
.A2(n_228),
.B1(n_231),
.B2(n_196),
.Y(n_235)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_168),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_220),
.B(n_221),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_168),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_178),
.B(n_36),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_229),
.Y(n_237)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_225),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_198),
.A2(n_23),
.B(n_24),
.C(n_8),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_166),
.B1(n_143),
.B2(n_149),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_177),
.A2(n_166),
.B1(n_143),
.B2(n_105),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_194),
.C(n_186),
.Y(n_236)
);

NOR3xp33_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_24),
.C(n_23),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_12),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_105),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_202),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_235),
.A2(n_260),
.B1(n_227),
.B2(n_1),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_211),
.C(n_206),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_245),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_223),
.A2(n_197),
.B1(n_186),
.B2(n_188),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_245),
.B1(n_261),
.B2(n_226),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

NOR4xp25_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_179),
.C(n_191),
.D(n_104),
.Y(n_244)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_87),
.C(n_9),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_230),
.B1(n_226),
.B2(n_234),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_246),
.B(n_205),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_257),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_210),
.B(n_218),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_249),
.A2(n_207),
.B(n_224),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_206),
.B(n_41),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_232),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_208),
.B(n_115),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_222),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_209),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_240),
.A2(n_213),
.B(n_217),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_281),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_264),
.A2(n_277),
.B1(n_282),
.B2(n_237),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_225),
.Y(n_265)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_278),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_248),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_279),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_273),
.C(n_275),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_261),
.Y(n_270)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_271),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_258),
.A2(n_255),
.B(n_249),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_258),
.B1(n_239),
.B2(n_238),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_211),
.C(n_219),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_236),
.B(n_216),
.C(n_229),
.Y(n_275)
);

NOR3xp33_ASAP7_75t_SL g279 ( 
.A(n_255),
.B(n_241),
.C(n_244),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_280),
.B(n_259),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_41),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_253),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_247),
.A2(n_10),
.B1(n_18),
.B2(n_17),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_253),
.C(n_257),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_241),
.B(n_7),
.Y(n_284)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_270),
.Y(n_314)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_286),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_256),
.B1(n_237),
.B2(n_251),
.Y(n_289)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_289),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_293),
.Y(n_310)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_294),
.Y(n_319)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_295),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_243),
.C(n_239),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_266),
.C(n_270),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_252),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_271),
.C(n_11),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_300),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_259),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_262),
.A2(n_248),
.B1(n_1),
.B2(n_2),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_276),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_272),
.B(n_273),
.Y(n_304)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_304),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_278),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_305),
.B(n_294),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_316),
.C(n_317),
.Y(n_327)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_311),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_293),
.A2(n_279),
.B(n_283),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_313),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_314),
.A2(n_299),
.B1(n_287),
.B2(n_3),
.Y(n_324)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_0),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_288),
.C(n_296),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_0),
.C(n_2),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_3),
.C(n_4),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_314),
.A2(n_291),
.B(n_297),
.Y(n_320)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_287),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_321),
.B(n_324),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_322),
.A2(n_308),
.B(n_317),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_291),
.B1(n_301),
.B2(n_303),
.Y(n_323)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_323),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_325),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_306),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_328),
.A2(n_310),
.B1(n_313),
.B2(n_319),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_11),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_309),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_334),
.B(n_335),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_318),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_336),
.A2(n_341),
.B1(n_324),
.B2(n_330),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_15),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_331),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_341)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_343),
.Y(n_353)
);

OA21x2_ASAP7_75t_SL g344 ( 
.A1(n_336),
.A2(n_327),
.B(n_326),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_345),
.Y(n_354)
);

O2A1O1Ixp33_ASAP7_75t_SL g345 ( 
.A1(n_337),
.A2(n_332),
.B(n_327),
.C(n_321),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_340),
.B(n_12),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_347),
.Y(n_355)
);

AO21x1_ASAP7_75t_L g347 ( 
.A1(n_333),
.A2(n_12),
.B(n_13),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_342),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_348),
.B(n_349),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_350),
.B(n_341),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_352),
.A2(n_349),
.B(n_346),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_356),
.B(n_357),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_353),
.B(n_338),
.C(n_18),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_338),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_359),
.A2(n_355),
.B(n_351),
.Y(n_360)
);

BUFx24_ASAP7_75t_SL g361 ( 
.A(n_360),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_361),
.B(n_354),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_362),
.B(n_18),
.Y(n_363)
);


endmodule