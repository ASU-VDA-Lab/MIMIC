module fake_jpeg_15514_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

BUFx3_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_4),
.B(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_13),
.B(n_17),
.Y(n_23)
);

AOI32xp33_ASAP7_75t_L g14 ( 
.A1(n_8),
.A2(n_12),
.A3(n_10),
.B1(n_11),
.B2(n_6),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_15),
.Y(n_27)
);

INVx4_ASAP7_75t_SL g15 ( 
.A(n_6),
.Y(n_15)
);

INVx3_ASAP7_75t_SL g16 ( 
.A(n_11),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_20),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_10),
.A2(n_0),
.B1(n_2),
.B2(n_5),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_7),
.B1(n_9),
.B2(n_17),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_6),
.A2(n_0),
.B1(n_2),
.B2(n_5),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_12),
.B1(n_7),
.B2(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_13),
.A2(n_2),
.B(n_7),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_16),
.B(n_15),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_26),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_9),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_31),
.B(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_27),
.C(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_35),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_30),
.Y(n_38)
);

AO21x2_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_29),
.B(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_36),
.Y(n_40)
);


endmodule