module fake_netlist_6_3300_n_1811 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1811);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1811;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1737;
wire n_236;
wire n_653;
wire n_1464;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_32),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_174),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_56),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_83),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_145),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_18),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_2),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_118),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_98),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_57),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_141),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_29),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_121),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_105),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_64),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_82),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_127),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_100),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_19),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_104),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_177),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_171),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_10),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_30),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_96),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_9),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_18),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_66),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_1),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_86),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_61),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_45),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_43),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_52),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_58),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_134),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_49),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_135),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_78),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_169),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_42),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_6),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_110),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_124),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_28),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_187),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_24),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_111),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_93),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_58),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_51),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_19),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_185),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_87),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_8),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_159),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_114),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_13),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_147),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_112),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_107),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_142),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_39),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_170),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_168),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_92),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_20),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_17),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_102),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_10),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_71),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_12),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_12),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_54),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_6),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_188),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_139),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_173),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_45),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_23),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_144),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_3),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_36),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_3),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_60),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_109),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_94),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_23),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_54),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_42),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_68),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_9),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_95),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_17),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_137),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_5),
.Y(n_291)
);

BUFx2_ASAP7_75t_SL g292 ( 
.A(n_38),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_50),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_43),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_157),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_129),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_156),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_67),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_75),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_80),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_128),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_34),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_26),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_1),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_182),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_103),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_158),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_70),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_90),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_181),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_34),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_8),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_130),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_29),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_13),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_0),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_123),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_4),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_32),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_89),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_136),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_55),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_11),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_108),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_154),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_57),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_180),
.Y(n_327)
);

BUFx10_ASAP7_75t_L g328 ( 
.A(n_39),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_138),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_37),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_47),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_15),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_49),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_56),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_176),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_53),
.Y(n_336)
);

BUFx2_ASAP7_75t_SL g337 ( 
.A(n_120),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_186),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_25),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_148),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_79),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_99),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_183),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_26),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_48),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_74),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_133),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_36),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_153),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_175),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_116),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_44),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_88),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_91),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_152),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_38),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_178),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_60),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_61),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_143),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_69),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_132),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_16),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_97),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_47),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_126),
.Y(n_366)
);

BUFx10_ASAP7_75t_L g367 ( 
.A(n_119),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_16),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_59),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_44),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_40),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_149),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_76),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_203),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_203),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_203),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_203),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_190),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_203),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_203),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_220),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_203),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_203),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_214),
.Y(n_384)
);

BUFx6f_ASAP7_75t_SL g385 ( 
.A(n_367),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_282),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_358),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_220),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_193),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_358),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_358),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_197),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_202),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_205),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_358),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_288),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_216),
.B(n_0),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_313),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_207),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_209),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_358),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_195),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_195),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_327),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_357),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_257),
.B(n_2),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_225),
.Y(n_407)
);

INVxp33_ASAP7_75t_SL g408 ( 
.A(n_279),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_257),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_279),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_189),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_192),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_192),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_357),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_211),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_254),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_198),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_198),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_212),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_217),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_225),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_267),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_267),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_319),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_223),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_233),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_227),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_234),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_237),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_238),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_242),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_243),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_247),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_208),
.B(n_4),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_248),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_208),
.B(n_5),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_301),
.B(n_7),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_250),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_251),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_319),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_255),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_196),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_260),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_196),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_215),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_264),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_266),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_215),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_224),
.Y(n_449)
);

CKINVDCx14_ASAP7_75t_R g450 ( 
.A(n_245),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_271),
.Y(n_451)
);

INVxp33_ASAP7_75t_SL g452 ( 
.A(n_191),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_272),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_224),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_241),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_301),
.B(n_14),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_241),
.Y(n_457)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_245),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_249),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_245),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_276),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_286),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_249),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_200),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_199),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_284),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_254),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_290),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_378),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_467),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_405),
.B(n_228),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_387),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_389),
.B(n_308),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_392),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_393),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_394),
.B(n_308),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_399),
.B(n_194),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_384),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_386),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_374),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_400),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_387),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_419),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_411),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_425),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_390),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_390),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_374),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_426),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_414),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_391),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_391),
.B(n_194),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_395),
.B(n_320),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_381),
.B(n_206),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_428),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_450),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_395),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_416),
.B(n_467),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_401),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_429),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_430),
.B(n_320),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_431),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_375),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_401),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_432),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_433),
.B(n_355),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_375),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_376),
.Y(n_508)
);

CKINVDCx8_ASAP7_75t_R g509 ( 
.A(n_435),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_376),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_407),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_377),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_377),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_439),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_407),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_396),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_441),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_442),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_443),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_442),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_447),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_444),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_451),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_452),
.B(n_232),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_453),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_412),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_462),
.B(n_355),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_444),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_379),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_415),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_445),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_388),
.B(n_305),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_458),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_445),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_398),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_409),
.B(n_307),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_420),
.Y(n_537)
);

OA21x2_ASAP7_75t_L g538 ( 
.A1(n_379),
.A2(n_382),
.B(n_380),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_464),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_380),
.Y(n_540)
);

BUFx6f_ASAP7_75t_SL g541 ( 
.A(n_413),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_438),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_406),
.B(n_302),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_427),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_448),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_446),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_461),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_543),
.B(n_524),
.Y(n_548)
);

OA22x2_ASAP7_75t_L g549 ( 
.A1(n_470),
.A2(n_410),
.B1(n_427),
.B2(n_418),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_526),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_470),
.B(n_417),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_526),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_529),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_480),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_477),
.B(n_408),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_526),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_544),
.Y(n_557)
);

NAND3xp33_ASAP7_75t_L g558 ( 
.A(n_543),
.B(n_436),
.C(n_434),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_498),
.B(n_460),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_544),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_498),
.B(n_465),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_501),
.B(n_382),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_529),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_540),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_538),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_538),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_540),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_469),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_538),
.A2(n_456),
.B1(n_437),
.B2(n_465),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_506),
.B(n_383),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_480),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_527),
.B(n_468),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_480),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_532),
.B(n_397),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_488),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_540),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_488),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_529),
.Y(n_578)
);

AO22x2_ASAP7_75t_L g579 ( 
.A1(n_471),
.A2(n_292),
.B1(n_365),
.B2(n_289),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_536),
.B(n_448),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_530),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_540),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_473),
.B(n_383),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_529),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_494),
.B(n_199),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_488),
.Y(n_586)
);

CKINVDCx6p67_ASAP7_75t_R g587 ( 
.A(n_478),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_503),
.Y(n_588)
);

BUFx10_ASAP7_75t_L g589 ( 
.A(n_474),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_476),
.B(n_201),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_539),
.B(n_262),
.Y(n_591)
);

INVx4_ASAP7_75t_SL g592 ( 
.A(n_529),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_509),
.B(n_201),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_538),
.B(n_295),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_529),
.B(n_296),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_503),
.Y(n_596)
);

OR2x6_ASAP7_75t_L g597 ( 
.A(n_490),
.B(n_484),
.Y(n_597)
);

AND2x6_ASAP7_75t_L g598 ( 
.A(n_503),
.B(n_204),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_475),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_509),
.B(n_204),
.Y(n_600)
);

AND2x2_ASAP7_75t_SL g601 ( 
.A(n_490),
.B(n_213),
.Y(n_601)
);

NAND2xp33_ASAP7_75t_R g602 ( 
.A(n_481),
.B(n_210),
.Y(n_602)
);

OR2x6_ASAP7_75t_L g603 ( 
.A(n_496),
.B(n_292),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_479),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_472),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_472),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_492),
.Y(n_607)
);

BUFx10_ASAP7_75t_L g608 ( 
.A(n_483),
.Y(n_608)
);

INVxp67_ASAP7_75t_SL g609 ( 
.A(n_507),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_472),
.Y(n_610)
);

INVx4_ASAP7_75t_SL g611 ( 
.A(n_541),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_SL g612 ( 
.A(n_541),
.B(n_236),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_485),
.B(n_489),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_507),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_492),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_495),
.A2(n_502),
.B1(n_505),
.B2(n_500),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_514),
.B(n_213),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_518),
.A2(n_311),
.B1(n_345),
.B2(n_339),
.Y(n_618)
);

NAND2xp33_ASAP7_75t_L g619 ( 
.A(n_507),
.B(n_222),
.Y(n_619)
);

BUFx6f_ASAP7_75t_SL g620 ( 
.A(n_518),
.Y(n_620)
);

INVxp67_ASAP7_75t_SL g621 ( 
.A(n_508),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_508),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_508),
.Y(n_623)
);

OR2x6_ASAP7_75t_L g624 ( 
.A(n_533),
.B(n_337),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_517),
.B(n_449),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_519),
.B(n_222),
.Y(n_626)
);

INVx8_ASAP7_75t_L g627 ( 
.A(n_521),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_523),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_525),
.B(n_240),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_510),
.B(n_297),
.Y(n_630)
);

AND3x2_ASAP7_75t_L g631 ( 
.A(n_492),
.B(n_256),
.C(n_240),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_472),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_520),
.B(n_466),
.Y(n_633)
);

NAND3xp33_ASAP7_75t_L g634 ( 
.A(n_520),
.B(n_219),
.C(n_218),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_510),
.B(n_512),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_522),
.Y(n_636)
);

BUFx8_ASAP7_75t_SL g637 ( 
.A(n_516),
.Y(n_637)
);

AND2x6_ASAP7_75t_L g638 ( 
.A(n_510),
.B(n_256),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_512),
.B(n_298),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_522),
.B(n_285),
.Y(n_640)
);

AOI21x1_ASAP7_75t_L g641 ( 
.A1(n_513),
.A2(n_273),
.B(n_259),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_513),
.B(n_299),
.Y(n_642)
);

AND3x2_ASAP7_75t_L g643 ( 
.A(n_492),
.B(n_273),
.C(n_259),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_513),
.B(n_300),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_528),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_482),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_482),
.B(n_306),
.Y(n_647)
);

INVx4_ASAP7_75t_L g648 ( 
.A(n_472),
.Y(n_648)
);

AND2x6_ASAP7_75t_L g649 ( 
.A(n_493),
.B(n_281),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_472),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_528),
.Y(n_651)
);

AND2x6_ASAP7_75t_L g652 ( 
.A(n_493),
.B(n_281),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_531),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_486),
.B(n_487),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_486),
.B(n_309),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_487),
.B(n_385),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_491),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_493),
.B(n_324),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_497),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_534),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_534),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_493),
.B(n_324),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_497),
.B(n_310),
.Y(n_663)
);

NOR2x1p5_ASAP7_75t_L g664 ( 
.A(n_537),
.B(n_227),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_499),
.B(n_317),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_541),
.A2(n_291),
.B1(n_315),
.B2(n_314),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_545),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_545),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_499),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_504),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_504),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_491),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_491),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_511),
.B(n_329),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_491),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_491),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_541),
.A2(n_385),
.B1(n_404),
.B2(n_321),
.Y(n_677)
);

INVxp33_ASAP7_75t_L g678 ( 
.A(n_511),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_491),
.B(n_325),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_515),
.B(n_385),
.Y(n_680)
);

INVxp67_ASAP7_75t_SL g681 ( 
.A(n_515),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_542),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_546),
.B(n_449),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_547),
.B(n_338),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_535),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_470),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_543),
.B(n_329),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_478),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_544),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_480),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_480),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_529),
.Y(n_692)
);

BUFx4f_ASAP7_75t_L g693 ( 
.A(n_538),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_529),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_538),
.A2(n_336),
.B1(n_339),
.B2(n_345),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_470),
.Y(n_696)
);

INVx4_ASAP7_75t_L g697 ( 
.A(n_529),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_498),
.B(n_342),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_583),
.B(n_574),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_555),
.B(n_221),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_554),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_557),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_607),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_693),
.B(n_343),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_607),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_615),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_562),
.B(n_335),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_554),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_571),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_615),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_693),
.B(n_346),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_683),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_570),
.B(n_335),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_561),
.B(n_340),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_555),
.B(n_226),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_563),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_561),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_548),
.A2(n_347),
.B1(n_362),
.B2(n_366),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_561),
.B(n_340),
.Y(n_719)
);

BUFx5_ASAP7_75t_L g720 ( 
.A(n_565),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_550),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_571),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_580),
.B(n_302),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_573),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_552),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_625),
.B(n_302),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_548),
.B(n_229),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_563),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_558),
.A2(n_354),
.B1(n_373),
.B2(n_372),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_683),
.B(n_231),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_594),
.A2(n_569),
.B(n_566),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_565),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_681),
.B(n_341),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_566),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_695),
.B(n_349),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_572),
.A2(n_687),
.B1(n_559),
.B2(n_556),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_551),
.B(n_316),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_695),
.A2(n_331),
.B1(n_284),
.B2(n_289),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_572),
.B(n_686),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_636),
.B(n_341),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_651),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_687),
.B(n_235),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_668),
.B(n_350),
.Y(n_743)
);

BUFx12f_ASAP7_75t_L g744 ( 
.A(n_589),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_560),
.Y(n_745)
);

INVx8_ASAP7_75t_L g746 ( 
.A(n_627),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_573),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_569),
.A2(n_331),
.B1(n_293),
.B2(n_294),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_551),
.B(n_351),
.Y(n_749)
);

BUFx8_ASAP7_75t_L g750 ( 
.A(n_620),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_653),
.B(n_350),
.Y(n_751)
);

NAND2xp33_ASAP7_75t_L g752 ( 
.A(n_649),
.B(n_353),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_551),
.B(n_360),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_564),
.B(n_361),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_591),
.B(n_246),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_SL g756 ( 
.A1(n_601),
.A2(n_258),
.B1(n_326),
.B2(n_367),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_689),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_678),
.B(n_239),
.Y(n_758)
);

NOR2x1_ASAP7_75t_L g759 ( 
.A(n_684),
.B(n_337),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_660),
.B(n_364),
.Y(n_760)
);

INVxp67_ASAP7_75t_SL g761 ( 
.A(n_563),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_661),
.B(n_454),
.Y(n_762)
);

INVxp67_ASAP7_75t_SL g763 ( 
.A(n_563),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_667),
.B(n_454),
.Y(n_764)
);

NOR2xp67_ASAP7_75t_L g765 ( 
.A(n_599),
.B(n_63),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_640),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_664),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_678),
.B(n_244),
.Y(n_768)
);

NOR2x1p5_ASAP7_75t_L g769 ( 
.A(n_568),
.B(n_246),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_686),
.B(n_228),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_696),
.B(n_316),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_L g772 ( 
.A1(n_549),
.A2(n_645),
.B1(n_585),
.B2(n_600),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_696),
.B(n_455),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_609),
.B(n_621),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_633),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_575),
.Y(n_776)
);

INVxp33_ASAP7_75t_L g777 ( 
.A(n_637),
.Y(n_777)
);

A2O1A1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_567),
.A2(n_277),
.B(n_294),
.C(n_304),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_669),
.B(n_455),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_671),
.B(n_457),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_630),
.B(n_457),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_575),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_577),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_604),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_639),
.B(n_459),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_646),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_642),
.B(n_459),
.Y(n_787)
);

INVx8_ASAP7_75t_L g788 ( 
.A(n_627),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_644),
.B(n_463),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_646),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_698),
.B(n_463),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_617),
.B(n_252),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_576),
.A2(n_336),
.B(n_365),
.C(n_334),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_582),
.B(n_466),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_659),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_617),
.B(n_263),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_590),
.B(n_265),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_590),
.B(n_268),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_SL g799 ( 
.A(n_628),
.B(n_367),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_601),
.B(n_367),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_626),
.B(n_269),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_647),
.B(n_270),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_670),
.B(n_626),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_618),
.A2(n_579),
.B1(n_619),
.B2(n_649),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_629),
.B(n_228),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_SL g806 ( 
.A(n_589),
.B(n_230),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_585),
.A2(n_330),
.B(n_293),
.C(n_304),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_655),
.B(n_274),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_603),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_663),
.B(n_275),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_629),
.B(n_278),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_603),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_584),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_673),
.B(n_230),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_654),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_665),
.B(n_280),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_577),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_604),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_602),
.A2(n_230),
.B1(n_253),
.B2(n_261),
.Y(n_819)
);

NOR2xp67_ASAP7_75t_L g820 ( 
.A(n_616),
.B(n_65),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_553),
.B(n_283),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_674),
.B(n_402),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_593),
.B(n_253),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_584),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_553),
.B(n_694),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_584),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_688),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_694),
.B(n_287),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_674),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_614),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_600),
.B(n_253),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_595),
.B(n_679),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_677),
.B(n_261),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_673),
.B(n_261),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_586),
.B(n_303),
.Y(n_835)
);

INVx4_ASAP7_75t_L g836 ( 
.A(n_692),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_588),
.B(n_596),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_614),
.B(n_312),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_674),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_603),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_634),
.B(n_318),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_622),
.B(n_322),
.Y(n_842)
);

AOI221xp5_ASAP7_75t_L g843 ( 
.A1(n_618),
.A2(n_311),
.B1(n_330),
.B2(n_334),
.C(n_359),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_658),
.B(n_662),
.Y(n_844)
);

AND2x6_ASAP7_75t_SL g845 ( 
.A(n_597),
.B(n_402),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_624),
.B(n_323),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_623),
.Y(n_847)
);

AND2x6_ASAP7_75t_SL g848 ( 
.A(n_597),
.B(n_403),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_690),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_690),
.B(n_332),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_691),
.B(n_333),
.Y(n_851)
);

BUFx8_ASAP7_75t_L g852 ( 
.A(n_620),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_691),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_579),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_624),
.B(n_344),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_624),
.B(n_348),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_692),
.B(n_371),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_635),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_602),
.A2(n_369),
.B1(n_352),
.B2(n_356),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_579),
.A2(n_619),
.B1(n_649),
.B2(n_652),
.Y(n_860)
);

NAND2xp33_ASAP7_75t_L g861 ( 
.A(n_649),
.B(n_652),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_692),
.B(n_363),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_649),
.A2(n_316),
.B1(n_328),
.B2(n_368),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_731),
.A2(n_676),
.B(n_675),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_832),
.A2(n_658),
.B(n_662),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_712),
.B(n_613),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_699),
.B(n_656),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_SL g868 ( 
.A(n_744),
.B(n_581),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_700),
.A2(n_656),
.B(n_680),
.C(n_612),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_717),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_734),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_717),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_815),
.B(n_652),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_702),
.Y(n_874)
);

AOI21x1_ASAP7_75t_L g875 ( 
.A1(n_704),
.A2(n_641),
.B(n_666),
.Y(n_875)
);

BUFx12f_ASAP7_75t_L g876 ( 
.A(n_750),
.Y(n_876)
);

NOR3xp33_ASAP7_75t_L g877 ( 
.A(n_700),
.B(n_613),
.C(n_612),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_715),
.A2(n_652),
.B1(n_682),
.B2(n_680),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_715),
.B(n_652),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_791),
.B(n_610),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_702),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_786),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_730),
.B(n_610),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_730),
.B(n_650),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_774),
.A2(n_697),
.B(n_578),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_790),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_748),
.B(n_650),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_792),
.A2(n_682),
.B(n_627),
.C(n_685),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_795),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_748),
.B(n_692),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_844),
.A2(n_598),
.B1(n_638),
.B2(n_589),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_732),
.B(n_598),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_766),
.B(n_608),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_739),
.B(n_608),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_772),
.A2(n_440),
.B(n_424),
.C(n_403),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_726),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_854),
.B(n_608),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_732),
.A2(n_697),
.B(n_578),
.Y(n_898)
);

OAI321xp33_ASAP7_75t_L g899 ( 
.A1(n_792),
.A2(n_423),
.A3(n_440),
.B1(n_421),
.B2(n_422),
.C(n_424),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_844),
.A2(n_736),
.B1(n_727),
.B2(n_803),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_704),
.A2(n_598),
.B(n_638),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_734),
.A2(n_581),
.B1(n_370),
.B2(n_688),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_745),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_858),
.B(n_598),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_723),
.B(n_587),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_758),
.B(n_611),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_861),
.A2(n_672),
.B(n_657),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_825),
.A2(n_672),
.B(n_657),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_711),
.A2(n_598),
.B(n_638),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_757),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_720),
.B(n_611),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_720),
.B(n_611),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_711),
.A2(n_648),
.B(n_605),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_781),
.B(n_638),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_758),
.B(n_328),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_761),
.A2(n_648),
.B(n_605),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_763),
.A2(n_632),
.B(n_606),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_741),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_738),
.A2(n_423),
.B(n_328),
.C(n_643),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_720),
.B(n_592),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_716),
.A2(n_826),
.B(n_728),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_720),
.B(n_592),
.Y(n_922)
);

NAND3xp33_ASAP7_75t_L g923 ( 
.A(n_796),
.B(n_631),
.C(n_632),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_827),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_785),
.B(n_638),
.Y(n_925)
);

AOI21x1_ASAP7_75t_L g926 ( 
.A1(n_837),
.A2(n_592),
.B(n_606),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_720),
.B(n_131),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_738),
.A2(n_637),
.B1(n_15),
.B2(n_20),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_771),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_829),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_716),
.A2(n_184),
.B(n_167),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_772),
.A2(n_14),
.B(n_21),
.C(n_22),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_787),
.B(n_21),
.Y(n_933)
);

NAND3xp33_ASAP7_75t_L g934 ( 
.A(n_796),
.B(n_22),
.C(n_24),
.Y(n_934)
);

OAI22x1_ASAP7_75t_L g935 ( 
.A1(n_819),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_935)
);

AO22x1_ASAP7_75t_L g936 ( 
.A1(n_801),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_720),
.B(n_77),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_728),
.A2(n_81),
.B(n_163),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_839),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_768),
.B(n_31),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_768),
.B(n_33),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_826),
.A2(n_84),
.B(n_162),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_800),
.A2(n_35),
.B(n_37),
.C(n_40),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_703),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_789),
.B(n_773),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_836),
.A2(n_85),
.B(n_161),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_836),
.A2(n_73),
.B(n_160),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_775),
.B(n_35),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_734),
.A2(n_72),
.B1(n_155),
.B2(n_151),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_701),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_801),
.A2(n_165),
.B1(n_150),
.B2(n_140),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_708),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_746),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_734),
.A2(n_117),
.B(n_115),
.Y(n_954)
);

NOR2xp67_ASAP7_75t_SL g955 ( 
.A(n_813),
.B(n_41),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_811),
.A2(n_113),
.B1(n_106),
.B2(n_101),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_804),
.A2(n_41),
.B1(n_46),
.B2(n_48),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_813),
.A2(n_46),
.B(n_50),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_800),
.B(n_51),
.Y(n_959)
);

NAND2x1p5_ASAP7_75t_L g960 ( 
.A(n_813),
.B(n_52),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_746),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_707),
.B(n_53),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_811),
.A2(n_55),
.B(n_59),
.C(n_62),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_713),
.B(n_62),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_813),
.A2(n_824),
.B(n_821),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_SL g966 ( 
.A1(n_735),
.A2(n_807),
.B(n_805),
.C(n_793),
.Y(n_966)
);

AND2x2_ASAP7_75t_SL g967 ( 
.A(n_860),
.B(n_804),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_820),
.B(n_860),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_824),
.A2(n_828),
.B(n_714),
.Y(n_969)
);

NAND3xp33_ASAP7_75t_L g970 ( 
.A(n_756),
.B(n_742),
.C(n_799),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_824),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_705),
.A2(n_706),
.B1(n_710),
.B2(n_863),
.Y(n_972)
);

NOR2x1p5_ASAP7_75t_SL g973 ( 
.A(n_709),
.B(n_722),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_824),
.A2(n_719),
.B(n_857),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_802),
.B(n_808),
.Y(n_975)
);

AOI22x1_ASAP7_75t_L g976 ( 
.A1(n_721),
.A2(n_725),
.B1(n_724),
.B2(n_782),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_747),
.A2(n_817),
.B(n_830),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_733),
.A2(n_838),
.B(n_851),
.C(n_751),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_822),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_863),
.A2(n_816),
.B1(n_810),
.B2(n_742),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_759),
.B(n_765),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_797),
.A2(n_798),
.B1(n_840),
.B2(n_760),
.Y(n_982)
);

O2A1O1Ixp5_ASAP7_75t_L g983 ( 
.A1(n_754),
.A2(n_851),
.B(n_838),
.C(n_862),
.Y(n_983)
);

O2A1O1Ixp5_ASAP7_75t_L g984 ( 
.A1(n_754),
.A2(n_850),
.B(n_740),
.C(n_743),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_752),
.A2(n_776),
.B(n_783),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_822),
.B(n_737),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_847),
.A2(n_849),
.B(n_853),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_835),
.A2(n_842),
.B(n_794),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_809),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_841),
.A2(n_805),
.B1(n_753),
.B2(n_749),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_749),
.A2(n_753),
.B(n_780),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_755),
.B(n_859),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_823),
.B(n_831),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_762),
.B(n_764),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_841),
.B(n_809),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_746),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_784),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_779),
.A2(n_770),
.B(n_834),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_812),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_718),
.B(n_729),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_778),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_846),
.A2(n_856),
.B(n_855),
.C(n_843),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_814),
.A2(n_834),
.B(n_767),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_814),
.A2(n_833),
.B(n_855),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_846),
.A2(n_856),
.B(n_812),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_806),
.B(n_788),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_788),
.A2(n_818),
.B(n_777),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_788),
.B(n_750),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_769),
.B(n_845),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_848),
.A2(n_693),
.B(n_774),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_852),
.A2(n_693),
.B(n_774),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_852),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_712),
.B(n_723),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_748),
.A2(n_731),
.B1(n_712),
.B2(n_736),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_702),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_774),
.A2(n_693),
.B(n_832),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_699),
.B(n_815),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_SL g1018 ( 
.A1(n_700),
.A2(n_715),
.B1(n_799),
.B2(n_543),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_699),
.B(n_815),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_774),
.A2(n_693),
.B(n_832),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_717),
.Y(n_1021)
);

NAND2xp33_ASAP7_75t_L g1022 ( 
.A(n_720),
.B(n_734),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_717),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_774),
.A2(n_693),
.B(n_832),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_717),
.Y(n_1025)
);

AO22x1_ASAP7_75t_L g1026 ( 
.A1(n_700),
.A2(n_715),
.B1(n_730),
.B2(n_792),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_717),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_772),
.A2(n_548),
.B(n_687),
.C(n_699),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_699),
.B(n_815),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_774),
.A2(n_693),
.B(n_832),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_774),
.A2(n_693),
.B(n_832),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_734),
.Y(n_1032)
);

AO21x1_ASAP7_75t_L g1033 ( 
.A1(n_800),
.A2(n_711),
.B(n_704),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_700),
.A2(n_715),
.B(n_796),
.C(n_792),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_699),
.B(n_815),
.Y(n_1035)
);

INVx11_ASAP7_75t_L g1036 ( 
.A(n_750),
.Y(n_1036)
);

AO22x1_ASAP7_75t_L g1037 ( 
.A1(n_700),
.A2(n_715),
.B1(n_730),
.B2(n_792),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_774),
.A2(n_693),
.B(n_832),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_731),
.A2(n_693),
.B(n_594),
.Y(n_1039)
);

INVxp67_ASAP7_75t_L g1040 ( 
.A(n_702),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_700),
.A2(n_715),
.B(n_796),
.C(n_792),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_699),
.B(n_815),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_717),
.Y(n_1043)
);

NAND3xp33_ASAP7_75t_SL g1044 ( 
.A(n_756),
.B(n_715),
.C(n_700),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_712),
.B(n_700),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_717),
.Y(n_1046)
);

AOI21x1_ASAP7_75t_L g1047 ( 
.A1(n_704),
.A2(n_711),
.B(n_594),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_699),
.B(n_815),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1045),
.B(n_1017),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_977),
.A2(n_926),
.B(n_985),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_1047),
.A2(n_1020),
.B(n_1016),
.Y(n_1051)
);

AOI21x1_ASAP7_75t_SL g1052 ( 
.A1(n_879),
.A2(n_1000),
.B(n_873),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_871),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1045),
.B(n_1019),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_1015),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_SL g1056 ( 
.A1(n_1034),
.A2(n_1041),
.B(n_968),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_1024),
.A2(n_1031),
.B(n_1030),
.Y(n_1057)
);

NOR2xp67_ASAP7_75t_L g1058 ( 
.A(n_896),
.B(n_929),
.Y(n_1058)
);

AO31x2_ASAP7_75t_L g1059 ( 
.A1(n_1033),
.A2(n_1014),
.A3(n_980),
.B(n_972),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_1038),
.A2(n_1039),
.B(n_968),
.Y(n_1060)
);

O2A1O1Ixp5_ASAP7_75t_L g1061 ( 
.A1(n_1026),
.A2(n_1037),
.B(n_884),
.C(n_883),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_965),
.A2(n_969),
.B(n_974),
.Y(n_1062)
);

INVx1_ASAP7_75t_SL g1063 ( 
.A(n_1015),
.Y(n_1063)
);

AOI221xp5_ASAP7_75t_SL g1064 ( 
.A1(n_1002),
.A2(n_957),
.B1(n_959),
.B2(n_932),
.C(n_1028),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1029),
.B(n_1035),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1042),
.B(n_1048),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_945),
.B(n_867),
.Y(n_1067)
);

AOI21x1_ASAP7_75t_L g1068 ( 
.A1(n_913),
.A2(n_875),
.B(n_991),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_900),
.A2(n_1018),
.B1(n_967),
.B2(n_990),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_874),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_SL g1071 ( 
.A1(n_871),
.A2(n_865),
.B(n_901),
.Y(n_1071)
);

AOI21x1_ASAP7_75t_L g1072 ( 
.A1(n_892),
.A2(n_885),
.B(n_914),
.Y(n_1072)
);

AOI21xp33_ASAP7_75t_L g1073 ( 
.A1(n_970),
.A2(n_915),
.B(n_866),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1013),
.B(n_905),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1022),
.A2(n_925),
.B(n_994),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_975),
.A2(n_880),
.B(n_907),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_866),
.B(n_940),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_1044),
.A2(n_959),
.B(n_941),
.C(n_877),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_908),
.A2(n_976),
.B(n_898),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_987),
.A2(n_864),
.B(n_909),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_890),
.A2(n_887),
.B(n_983),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_967),
.B(n_918),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_916),
.A2(n_917),
.B(n_921),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_963),
.A2(n_869),
.A3(n_1001),
.B(n_982),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_986),
.B(n_930),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_920),
.A2(n_922),
.B(n_904),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_984),
.A2(n_978),
.B(n_988),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_911),
.A2(n_912),
.B(n_998),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_939),
.B(n_933),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_881),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_995),
.B(n_894),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_966),
.A2(n_981),
.B(n_927),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_966),
.A2(n_981),
.B(n_927),
.Y(n_1093)
);

AO31x2_ASAP7_75t_L g1094 ( 
.A1(n_963),
.A2(n_888),
.A3(n_964),
.B(n_962),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_996),
.Y(n_1095)
);

NAND2x1p5_ASAP7_75t_L g1096 ( 
.A(n_871),
.B(n_996),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_937),
.A2(n_1004),
.B(n_1010),
.Y(n_1097)
);

O2A1O1Ixp5_ASAP7_75t_L g1098 ( 
.A1(n_937),
.A2(n_1011),
.B(n_995),
.C(n_1003),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_928),
.A2(n_943),
.B(n_895),
.C(n_934),
.Y(n_1099)
);

O2A1O1Ixp5_ASAP7_75t_L g1100 ( 
.A1(n_993),
.A2(n_948),
.B(n_936),
.C(n_1005),
.Y(n_1100)
);

NAND2x2_ASAP7_75t_L g1101 ( 
.A(n_997),
.B(n_903),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_950),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_SL g1103 ( 
.A(n_868),
.B(n_953),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_952),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_993),
.A2(n_894),
.B(n_878),
.C(n_992),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_870),
.A2(n_1021),
.B(n_872),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_886),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1027),
.A2(n_1046),
.B(n_1043),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_906),
.A2(n_899),
.B(n_1025),
.Y(n_1109)
);

OAI21xp33_ASAP7_75t_SL g1110 ( 
.A1(n_928),
.A2(n_944),
.B(n_889),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_SL g1111 ( 
.A1(n_891),
.A2(n_931),
.B(n_947),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1023),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1032),
.A2(n_938),
.B(n_946),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1032),
.Y(n_1114)
);

AOI21x1_ASAP7_75t_SL g1115 ( 
.A1(n_1009),
.A2(n_999),
.B(n_989),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_996),
.B(n_979),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_942),
.A2(n_954),
.B(n_949),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_924),
.B(n_1040),
.Y(n_1118)
);

NOR2x1_ASAP7_75t_R g1119 ( 
.A(n_876),
.B(n_961),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_923),
.A2(n_871),
.B(n_1006),
.Y(n_1120)
);

OR2x6_ASAP7_75t_L g1121 ( 
.A(n_996),
.B(n_1007),
.Y(n_1121)
);

OAI22x1_ASAP7_75t_L g1122 ( 
.A1(n_989),
.A2(n_999),
.B1(n_897),
.B2(n_893),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_897),
.A2(n_956),
.B(n_951),
.C(n_893),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_979),
.B(n_971),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_971),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_958),
.A2(n_960),
.B(n_1006),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_971),
.A2(n_979),
.B(n_919),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_979),
.B(n_919),
.Y(n_1128)
);

NAND2x1_ASAP7_75t_L g1129 ( 
.A(n_971),
.B(n_955),
.Y(n_1129)
);

AOI21x1_ASAP7_75t_L g1130 ( 
.A1(n_973),
.A2(n_935),
.B(n_902),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_960),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_910),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1008),
.B(n_1012),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1036),
.A2(n_977),
.B(n_926),
.Y(n_1134)
);

AOI221x1_ASAP7_75t_L g1135 ( 
.A1(n_1034),
.A2(n_1041),
.B1(n_1044),
.B2(n_877),
.C(n_970),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1045),
.B(n_1017),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_977),
.A2(n_926),
.B(n_985),
.Y(n_1137)
);

INVx4_ASAP7_75t_L g1138 ( 
.A(n_996),
.Y(n_1138)
);

NOR3xp33_ASAP7_75t_L g1139 ( 
.A(n_1044),
.B(n_1037),
.C(n_1026),
.Y(n_1139)
);

OAI21xp33_ASAP7_75t_L g1140 ( 
.A1(n_1045),
.A2(n_700),
.B(n_715),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1045),
.B(n_1017),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_871),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1013),
.B(n_712),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1045),
.B(n_1017),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1034),
.A2(n_1041),
.B(n_731),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1045),
.B(n_1017),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_977),
.A2(n_926),
.B(n_985),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1016),
.A2(n_1024),
.B(n_1020),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1016),
.A2(n_1024),
.B(n_1020),
.Y(n_1149)
);

NOR2xp67_ASAP7_75t_L g1150 ( 
.A(n_896),
.B(n_599),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1045),
.B(n_1017),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_977),
.A2(n_926),
.B(n_985),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1034),
.A2(n_1041),
.B(n_731),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_1033),
.A2(n_1041),
.A3(n_1034),
.B(n_1014),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1045),
.B(n_1017),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1034),
.A2(n_1041),
.B(n_731),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_996),
.B(n_979),
.Y(n_1157)
);

OAI211xp5_ASAP7_75t_L g1158 ( 
.A1(n_928),
.A2(n_756),
.B(n_1018),
.C(n_700),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_977),
.A2(n_926),
.B(n_985),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1016),
.A2(n_1024),
.B(n_1020),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1045),
.B(n_1017),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1016),
.A2(n_1024),
.B(n_1020),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1013),
.B(n_712),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1034),
.A2(n_1041),
.B(n_731),
.Y(n_1164)
);

OAI22x1_ASAP7_75t_L g1165 ( 
.A1(n_970),
.A2(n_1045),
.B1(n_548),
.B2(n_866),
.Y(n_1165)
);

AND3x4_ASAP7_75t_L g1166 ( 
.A(n_877),
.B(n_818),
.C(n_784),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_996),
.B(n_979),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1013),
.B(n_712),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_882),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_882),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_996),
.B(n_979),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_871),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1034),
.A2(n_1041),
.B(n_1044),
.C(n_1045),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1016),
.A2(n_1024),
.B(n_1020),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1045),
.B(n_1017),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_977),
.A2(n_926),
.B(n_985),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_977),
.A2(n_926),
.B(n_985),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1045),
.B(n_1017),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1015),
.Y(n_1179)
);

OAI22x1_ASAP7_75t_L g1180 ( 
.A1(n_970),
.A2(n_1045),
.B1(n_548),
.B2(n_866),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1045),
.B(n_712),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1016),
.A2(n_1024),
.B(n_1020),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_871),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1034),
.A2(n_1041),
.B(n_1044),
.C(n_1045),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_977),
.A2(n_926),
.B(n_985),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_977),
.A2(n_926),
.B(n_985),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1034),
.B(n_1041),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1034),
.A2(n_1041),
.B1(n_900),
.B2(n_1018),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1045),
.B(n_1017),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_SL g1190 ( 
.A1(n_1018),
.A2(n_756),
.B(n_715),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1045),
.B(n_1017),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1034),
.B(n_1041),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1036),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1034),
.A2(n_1041),
.B(n_1044),
.C(n_1045),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_977),
.A2(n_926),
.B(n_985),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_977),
.A2(n_926),
.B(n_985),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1036),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_977),
.A2(n_926),
.B(n_985),
.Y(n_1198)
);

AO21x1_ASAP7_75t_L g1199 ( 
.A1(n_1014),
.A2(n_980),
.B(n_968),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1016),
.A2(n_1024),
.B(n_1020),
.Y(n_1200)
);

NAND2x1p5_ASAP7_75t_L g1201 ( 
.A(n_1095),
.B(n_1138),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1067),
.B(n_1065),
.Y(n_1202)
);

OR2x6_ASAP7_75t_L g1203 ( 
.A(n_1121),
.B(n_1131),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1169),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1193),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1066),
.B(n_1049),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1142),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1050),
.A2(n_1147),
.B(n_1137),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1197),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1170),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1102),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_1179),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1104),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1090),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1142),
.Y(n_1215)
);

NAND2x1p5_ASAP7_75t_L g1216 ( 
.A(n_1095),
.B(n_1138),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1143),
.B(n_1163),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1142),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1054),
.B(n_1136),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_R g1220 ( 
.A(n_1103),
.B(n_1130),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1112),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1168),
.B(n_1074),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_SL g1223 ( 
.A(n_1140),
.B(n_1190),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1139),
.A2(n_1069),
.B1(n_1188),
.B2(n_1073),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1132),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_1118),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1183),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1141),
.A2(n_1146),
.B1(n_1189),
.B2(n_1144),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1091),
.B(n_1151),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_1101),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1155),
.B(n_1161),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1085),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1070),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1187),
.A2(n_1192),
.B(n_1056),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1175),
.B(n_1178),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1058),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_SL g1237 ( 
.A(n_1173),
.B(n_1184),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1191),
.A2(n_1158),
.B1(n_1194),
.B2(n_1164),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1116),
.B(n_1157),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1183),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1077),
.B(n_1181),
.Y(n_1241)
);

BUFx2_ASAP7_75t_SL g1242 ( 
.A(n_1167),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1082),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1158),
.A2(n_1145),
.B1(n_1156),
.B2(n_1153),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1089),
.Y(n_1245)
);

NAND2x1p5_ASAP7_75t_L g1246 ( 
.A(n_1167),
.B(n_1171),
.Y(n_1246)
);

INVx3_ASAP7_75t_SL g1247 ( 
.A(n_1133),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1133),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1105),
.B(n_1064),
.Y(n_1249)
);

NAND3xp33_ASAP7_75t_L g1250 ( 
.A(n_1139),
.B(n_1135),
.C(n_1078),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1192),
.A2(n_1099),
.B1(n_1123),
.B2(n_1166),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1165),
.B(n_1180),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_1128),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1114),
.Y(n_1254)
);

BUFx10_ASAP7_75t_L g1255 ( 
.A(n_1131),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1150),
.B(n_1122),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1125),
.Y(n_1257)
);

BUFx4f_ASAP7_75t_SL g1258 ( 
.A(n_1131),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1166),
.A2(n_1110),
.B1(n_1199),
.B2(n_1123),
.Y(n_1259)
);

INVx6_ASAP7_75t_SL g1260 ( 
.A(n_1121),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_R g1261 ( 
.A(n_1053),
.B(n_1172),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1154),
.B(n_1099),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1172),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1057),
.A2(n_1200),
.B(n_1182),
.Y(n_1264)
);

AO21x2_ASAP7_75t_L g1265 ( 
.A1(n_1057),
.A2(n_1200),
.B(n_1182),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1183),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1120),
.B(n_1124),
.Y(n_1267)
);

AOI221xp5_ASAP7_75t_L g1268 ( 
.A1(n_1100),
.A2(n_1092),
.B1(n_1093),
.B2(n_1061),
.C(n_1081),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1100),
.B(n_1120),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1121),
.B(n_1127),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1071),
.A2(n_1129),
.B1(n_1127),
.B2(n_1109),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1084),
.B(n_1154),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1126),
.A2(n_1097),
.B1(n_1109),
.B2(n_1106),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1060),
.A2(n_1075),
.B1(n_1096),
.B2(n_1183),
.Y(n_1274)
);

NAND2x1p5_ASAP7_75t_L g1275 ( 
.A(n_1134),
.B(n_1086),
.Y(n_1275)
);

INVx5_ASAP7_75t_L g1276 ( 
.A(n_1052),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1154),
.B(n_1059),
.Y(n_1277)
);

AND2x2_ASAP7_75t_SL g1278 ( 
.A(n_1154),
.B(n_1119),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1059),
.B(n_1084),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_SL g1280 ( 
.A(n_1115),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1098),
.A2(n_1061),
.B(n_1060),
.C(n_1097),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1108),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1059),
.B(n_1075),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1094),
.Y(n_1284)
);

INVx5_ASAP7_75t_L g1285 ( 
.A(n_1052),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1094),
.Y(n_1286)
);

INVxp67_ASAP7_75t_L g1287 ( 
.A(n_1115),
.Y(n_1287)
);

O2A1O1Ixp5_ASAP7_75t_L g1288 ( 
.A1(n_1098),
.A2(n_1148),
.B(n_1174),
.C(n_1162),
.Y(n_1288)
);

NAND2x1p5_ASAP7_75t_L g1289 ( 
.A(n_1117),
.B(n_1088),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1051),
.B(n_1068),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1148),
.A2(n_1174),
.B(n_1162),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1152),
.A2(n_1198),
.B(n_1176),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_SL g1293 ( 
.A(n_1149),
.B(n_1160),
.C(n_1111),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1080),
.A2(n_1160),
.B(n_1149),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1113),
.B(n_1062),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1072),
.Y(n_1296)
);

INVx4_ASAP7_75t_L g1297 ( 
.A(n_1159),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1177),
.Y(n_1298)
);

AOI221xp5_ASAP7_75t_L g1299 ( 
.A1(n_1079),
.A2(n_1083),
.B1(n_1185),
.B2(n_1186),
.C(n_1195),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1196),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1116),
.B(n_1157),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1140),
.A2(n_1044),
.B1(n_1018),
.B2(n_1139),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1076),
.A2(n_1020),
.B(n_1016),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1063),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1116),
.B(n_1157),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1107),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1116),
.B(n_1157),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1142),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1067),
.B(n_1065),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1076),
.A2(n_1020),
.B(n_1016),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1193),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1076),
.A2(n_1020),
.B(n_1016),
.Y(n_1312)
);

NOR2x1p5_ASAP7_75t_L g1313 ( 
.A(n_1077),
.B(n_587),
.Y(n_1313)
);

BUFx10_ASAP7_75t_L g1314 ( 
.A(n_1133),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1067),
.B(n_1065),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1140),
.B(n_1045),
.Y(n_1316)
);

NAND2x1p5_ASAP7_75t_L g1317 ( 
.A(n_1095),
.B(n_1138),
.Y(n_1317)
);

OR2x6_ASAP7_75t_L g1318 ( 
.A(n_1121),
.B(n_746),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1143),
.B(n_1013),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1143),
.B(n_1013),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1055),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1055),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1076),
.A2(n_1020),
.B(n_1016),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1076),
.A2(n_1020),
.B(n_1016),
.Y(n_1324)
);

OR2x6_ASAP7_75t_L g1325 ( 
.A(n_1121),
.B(n_746),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1076),
.A2(n_1020),
.B(n_1016),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1140),
.B(n_1045),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1055),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1055),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1090),
.Y(n_1330)
);

OR2x6_ASAP7_75t_L g1331 ( 
.A(n_1121),
.B(n_746),
.Y(n_1331)
);

NAND2xp33_ASAP7_75t_L g1332 ( 
.A(n_1140),
.B(n_1034),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1076),
.A2(n_1020),
.B(n_1016),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1076),
.A2(n_1020),
.B(n_1016),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1143),
.B(n_1013),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1107),
.Y(n_1336)
);

CKINVDCx11_ASAP7_75t_R g1337 ( 
.A(n_1101),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1205),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1224),
.A2(n_1332),
.B(n_1327),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1203),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1260),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1306),
.Y(n_1342)
);

CKINVDCx14_ASAP7_75t_R g1343 ( 
.A(n_1209),
.Y(n_1343)
);

NAND2x1p5_ASAP7_75t_L g1344 ( 
.A(n_1253),
.B(n_1270),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1208),
.A2(n_1292),
.B(n_1303),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1223),
.B(n_1243),
.Y(n_1346)
);

BUFx2_ASAP7_75t_R g1347 ( 
.A(n_1311),
.Y(n_1347)
);

OA21x2_ASAP7_75t_L g1348 ( 
.A1(n_1288),
.A2(n_1294),
.B(n_1291),
.Y(n_1348)
);

AO21x1_ASAP7_75t_L g1349 ( 
.A1(n_1251),
.A2(n_1244),
.B(n_1237),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1223),
.B(n_1253),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_1226),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1203),
.Y(n_1352)
);

BUFx8_ASAP7_75t_L g1353 ( 
.A(n_1212),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1204),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1310),
.A2(n_1323),
.B(n_1312),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1210),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1233),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1321),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1324),
.A2(n_1333),
.B(n_1326),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1211),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1334),
.A2(n_1264),
.B(n_1275),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1213),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1302),
.B(n_1251),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1254),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1265),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1255),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1260),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1322),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1221),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1257),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1245),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1329),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1237),
.A2(n_1316),
.B1(n_1244),
.B2(n_1250),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1232),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1250),
.A2(n_1220),
.B1(n_1238),
.B2(n_1278),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1222),
.B(n_1217),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1263),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1293),
.A2(n_1294),
.B(n_1281),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1238),
.A2(n_1228),
.B1(n_1234),
.B2(n_1206),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1252),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1296),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1255),
.Y(n_1382)
);

CKINVDCx11_ASAP7_75t_R g1383 ( 
.A(n_1247),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1202),
.B(n_1309),
.Y(n_1384)
);

AO21x1_ASAP7_75t_L g1385 ( 
.A1(n_1269),
.A2(n_1271),
.B(n_1259),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1252),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1258),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1241),
.A2(n_1249),
.B1(n_1228),
.B2(n_1319),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1282),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1276),
.B(n_1285),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1286),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1206),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1202),
.B(n_1315),
.Y(n_1393)
);

AOI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1313),
.A2(n_1248),
.B1(n_1315),
.B2(n_1335),
.Y(n_1394)
);

AOI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1271),
.A2(n_1295),
.B(n_1300),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1249),
.A2(n_1320),
.B1(n_1256),
.B2(n_1262),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1262),
.A2(n_1267),
.B1(n_1235),
.B2(n_1231),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1304),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1266),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1219),
.A2(n_1231),
.B1(n_1235),
.B2(n_1225),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1328),
.Y(n_1401)
);

INVx6_ASAP7_75t_L g1402 ( 
.A(n_1314),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1308),
.Y(n_1403)
);

AOI21xp33_ASAP7_75t_SL g1404 ( 
.A1(n_1230),
.A2(n_1236),
.B(n_1219),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1308),
.Y(n_1405)
);

AO21x1_ASAP7_75t_L g1406 ( 
.A1(n_1283),
.A2(n_1274),
.B(n_1273),
.Y(n_1406)
);

CKINVDCx11_ASAP7_75t_R g1407 ( 
.A(n_1337),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1268),
.A2(n_1272),
.B1(n_1284),
.B2(n_1280),
.Y(n_1408)
);

AO21x2_ASAP7_75t_L g1409 ( 
.A1(n_1290),
.A2(n_1274),
.B(n_1295),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1214),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1330),
.A2(n_1331),
.B1(n_1325),
.B2(n_1318),
.Y(n_1411)
);

AO21x2_ASAP7_75t_L g1412 ( 
.A1(n_1277),
.A2(n_1279),
.B(n_1287),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1207),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1318),
.A2(n_1331),
.B1(n_1325),
.B2(n_1242),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1275),
.A2(n_1289),
.B(n_1299),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1289),
.A2(n_1298),
.B(n_1325),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1331),
.A2(n_1277),
.B1(n_1279),
.B2(n_1305),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1261),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1239),
.B(n_1301),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1276),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1307),
.A2(n_1276),
.B1(n_1285),
.B2(n_1246),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1215),
.B(n_1218),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1246),
.B(n_1240),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1201),
.A2(n_1317),
.B(n_1216),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_SL g1425 ( 
.A1(n_1285),
.A2(n_1215),
.B1(n_1218),
.B2(n_1227),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1297),
.A2(n_1158),
.B1(n_806),
.B2(n_799),
.Y(n_1426)
);

INVx6_ASAP7_75t_L g1427 ( 
.A(n_1314),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1223),
.A2(n_1044),
.B1(n_1018),
.B2(n_1140),
.Y(n_1428)
);

OAI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1223),
.A2(n_799),
.B1(n_806),
.B2(n_1190),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1226),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1223),
.A2(n_1044),
.B1(n_1018),
.B2(n_1140),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1223),
.A2(n_1044),
.B1(n_1018),
.B2(n_1140),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1336),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1336),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1223),
.A2(n_1044),
.B1(n_1018),
.B2(n_1140),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1270),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1288),
.A2(n_1087),
.B(n_1294),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1223),
.B(n_1243),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1223),
.B(n_1243),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1229),
.B(n_1202),
.Y(n_1440)
);

BUFx12f_ASAP7_75t_SL g1441 ( 
.A(n_1203),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1429),
.A2(n_1339),
.B1(n_1440),
.B2(n_1394),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1344),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1363),
.B(n_1384),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1391),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1342),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1363),
.B(n_1384),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1398),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1393),
.B(n_1380),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1412),
.B(n_1386),
.Y(n_1450)
);

OR2x6_ASAP7_75t_L g1451 ( 
.A(n_1416),
.B(n_1385),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1340),
.A2(n_1352),
.B(n_1344),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1393),
.B(n_1350),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_1381),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1412),
.Y(n_1455)
);

NOR2xp67_ASAP7_75t_L g1456 ( 
.A(n_1404),
.B(n_1376),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1346),
.B(n_1438),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1438),
.B(n_1439),
.Y(n_1458)
);

INVx4_ASAP7_75t_L g1459 ( 
.A(n_1402),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1389),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1345),
.A2(n_1415),
.B(n_1361),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1418),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1402),
.Y(n_1463)
);

BUFx4f_ASAP7_75t_SL g1464 ( 
.A(n_1418),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1401),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1370),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1353),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1354),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1356),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1436),
.B(n_1349),
.Y(n_1470)
);

OR2x6_ASAP7_75t_L g1471 ( 
.A(n_1385),
.B(n_1395),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1360),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1410),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1362),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1364),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1400),
.B(n_1392),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1409),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1371),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1374),
.Y(n_1479)
);

CKINVDCx11_ASAP7_75t_R g1480 ( 
.A(n_1407),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1433),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1409),
.Y(n_1482)
);

OAI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1428),
.A2(n_1431),
.B(n_1432),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1434),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1365),
.Y(n_1485)
);

INVx6_ASAP7_75t_L g1486 ( 
.A(n_1353),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1349),
.B(n_1373),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1353),
.Y(n_1488)
);

OA21x2_ASAP7_75t_L g1489 ( 
.A1(n_1355),
.A2(n_1359),
.B(n_1406),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1378),
.B(n_1437),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1397),
.B(n_1396),
.Y(n_1491)
);

CKINVDCx20_ASAP7_75t_R g1492 ( 
.A(n_1351),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1409),
.Y(n_1493)
);

NOR2x1_ASAP7_75t_SL g1494 ( 
.A(n_1378),
.B(n_1420),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1406),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1357),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_1351),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1348),
.Y(n_1498)
);

INVx4_ASAP7_75t_L g1499 ( 
.A(n_1427),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1375),
.B(n_1379),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1410),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1355),
.A2(n_1359),
.B(n_1390),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1357),
.Y(n_1503)
);

INVx4_ASAP7_75t_R g1504 ( 
.A(n_1358),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1369),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1377),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1399),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1403),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1424),
.A2(n_1411),
.B(n_1421),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1450),
.B(n_1408),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1470),
.B(n_1417),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1450),
.B(n_1388),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1455),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1470),
.B(n_1435),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1495),
.B(n_1426),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1454),
.B(n_1487),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1445),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1483),
.A2(n_1500),
.B1(n_1442),
.B2(n_1487),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1490),
.B(n_1368),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1498),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1471),
.B(n_1405),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1460),
.B(n_1414),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1491),
.A2(n_1430),
.B1(n_1441),
.B2(n_1383),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1471),
.B(n_1423),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1471),
.B(n_1423),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1485),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1471),
.B(n_1413),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1460),
.B(n_1425),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1477),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1477),
.B(n_1422),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1482),
.B(n_1422),
.Y(n_1531)
);

INVxp67_ASAP7_75t_L g1532 ( 
.A(n_1448),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1444),
.B(n_1382),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1482),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1494),
.B(n_1422),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1493),
.B(n_1419),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1493),
.B(n_1419),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1519),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1536),
.B(n_1457),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1516),
.B(n_1453),
.Y(n_1540)
);

NOR3xp33_ASAP7_75t_L g1541 ( 
.A(n_1522),
.B(n_1476),
.C(n_1456),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_SL g1542 ( 
.A1(n_1514),
.A2(n_1451),
.B1(n_1486),
.B2(n_1458),
.Y(n_1542)
);

OA21x2_ASAP7_75t_L g1543 ( 
.A1(n_1520),
.A2(n_1461),
.B(n_1502),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1518),
.A2(n_1451),
.B1(n_1486),
.B2(n_1473),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1536),
.B(n_1457),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1537),
.B(n_1458),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1518),
.A2(n_1451),
.B1(n_1486),
.B2(n_1497),
.Y(n_1547)
);

AND2x2_ASAP7_75t_SL g1548 ( 
.A(n_1511),
.B(n_1489),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1516),
.B(n_1449),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1519),
.B(n_1449),
.Y(n_1550)
);

OAI221xp5_ASAP7_75t_L g1551 ( 
.A1(n_1523),
.A2(n_1367),
.B1(n_1341),
.B2(n_1462),
.C(n_1465),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1523),
.B(n_1459),
.Y(n_1552)
);

NOR2xp67_ASAP7_75t_L g1553 ( 
.A(n_1520),
.B(n_1463),
.Y(n_1553)
);

NAND3xp33_ASAP7_75t_L g1554 ( 
.A(n_1515),
.B(n_1501),
.C(n_1507),
.Y(n_1554)
);

OAI221xp5_ASAP7_75t_SL g1555 ( 
.A1(n_1514),
.A2(n_1452),
.B1(n_1341),
.B2(n_1367),
.C(n_1447),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1532),
.B(n_1478),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1530),
.B(n_1446),
.Y(n_1557)
);

NAND3xp33_ASAP7_75t_SL g1558 ( 
.A(n_1522),
.B(n_1492),
.C(n_1497),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1519),
.B(n_1479),
.Y(n_1559)
);

NAND3xp33_ASAP7_75t_L g1560 ( 
.A(n_1515),
.B(n_1481),
.C(n_1484),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1531),
.B(n_1509),
.Y(n_1561)
);

AOI221x1_ASAP7_75t_SL g1562 ( 
.A1(n_1517),
.A2(n_1475),
.B1(n_1474),
.B2(n_1472),
.C(n_1469),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1526),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1524),
.B(n_1509),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1524),
.B(n_1525),
.Y(n_1565)
);

NAND3xp33_ASAP7_75t_L g1566 ( 
.A(n_1515),
.B(n_1505),
.C(n_1506),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1533),
.B(n_1466),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1510),
.A2(n_1452),
.B(n_1443),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1533),
.B(n_1468),
.Y(n_1569)
);

OAI221xp5_ASAP7_75t_SL g1570 ( 
.A1(n_1510),
.A2(n_1462),
.B1(n_1467),
.B2(n_1488),
.C(n_1443),
.Y(n_1570)
);

NOR3xp33_ASAP7_75t_L g1571 ( 
.A(n_1510),
.B(n_1480),
.C(n_1499),
.Y(n_1571)
);

OAI221xp5_ASAP7_75t_SL g1572 ( 
.A1(n_1511),
.A2(n_1488),
.B1(n_1467),
.B2(n_1496),
.C(n_1503),
.Y(n_1572)
);

NAND2xp33_ASAP7_75t_SL g1573 ( 
.A(n_1528),
.B(n_1492),
.Y(n_1573)
);

OAI21xp33_ASAP7_75t_L g1574 ( 
.A1(n_1512),
.A2(n_1503),
.B(n_1496),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1563),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1563),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1538),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1543),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1559),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1559),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1549),
.B(n_1529),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1540),
.B(n_1529),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1556),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1548),
.B(n_1527),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1557),
.Y(n_1585)
);

NOR2xp67_ASAP7_75t_L g1586 ( 
.A(n_1566),
.B(n_1520),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1548),
.B(n_1527),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1550),
.B(n_1534),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1548),
.B(n_1521),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1564),
.B(n_1565),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1565),
.B(n_1521),
.Y(n_1591)
);

NAND3xp33_ASAP7_75t_L g1592 ( 
.A(n_1541),
.B(n_1508),
.C(n_1521),
.Y(n_1592)
);

AND2x4_ASAP7_75t_SL g1593 ( 
.A(n_1571),
.B(n_1535),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1553),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1561),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1564),
.Y(n_1596)
);

OR2x2_ASAP7_75t_SL g1597 ( 
.A(n_1558),
.B(n_1486),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1567),
.B(n_1569),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1562),
.B(n_1513),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1575),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1578),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1580),
.B(n_1562),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1594),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1596),
.B(n_1539),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1586),
.A2(n_1566),
.B(n_1547),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1575),
.Y(n_1606)
);

OAI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1592),
.A2(n_1547),
.B1(n_1544),
.B2(n_1551),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1586),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1576),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1596),
.B(n_1539),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1578),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1594),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1576),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1577),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1577),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1588),
.Y(n_1616)
);

AOI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1592),
.A2(n_1544),
.B1(n_1573),
.B2(n_1552),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1596),
.B(n_1545),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1595),
.B(n_1584),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1579),
.B(n_1583),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1588),
.Y(n_1621)
);

NAND2x1p5_ASAP7_75t_L g1622 ( 
.A(n_1589),
.B(n_1553),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1588),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1584),
.B(n_1546),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1581),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1585),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1584),
.B(n_1546),
.Y(n_1627)
);

OAI21xp33_ASAP7_75t_L g1628 ( 
.A1(n_1617),
.A2(n_1574),
.B(n_1555),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1600),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1600),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1603),
.Y(n_1631)
);

AOI21xp33_ASAP7_75t_L g1632 ( 
.A1(n_1607),
.A2(n_1599),
.B(n_1554),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1624),
.B(n_1587),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1602),
.B(n_1583),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1602),
.B(n_1480),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1606),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1603),
.B(n_1593),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1606),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1624),
.B(n_1598),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1609),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1609),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1624),
.B(n_1587),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1613),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1627),
.B(n_1598),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1627),
.B(n_1587),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1608),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1613),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1614),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1616),
.B(n_1582),
.Y(n_1649)
);

NOR2xp67_ASAP7_75t_L g1650 ( 
.A(n_1605),
.B(n_1589),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1625),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1627),
.B(n_1589),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1622),
.B(n_1590),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1622),
.B(n_1590),
.Y(n_1654)
);

INVx2_ASAP7_75t_SL g1655 ( 
.A(n_1622),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1614),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_SL g1657 ( 
.A(n_1605),
.B(n_1572),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1615),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1616),
.B(n_1582),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1619),
.Y(n_1660)
);

OAI21xp33_ASAP7_75t_L g1661 ( 
.A1(n_1617),
.A2(n_1574),
.B(n_1599),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1622),
.B(n_1590),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1604),
.B(n_1610),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1615),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1621),
.B(n_1591),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1612),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1626),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1621),
.B(n_1591),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1604),
.B(n_1590),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1619),
.Y(n_1670)
);

NAND2xp33_ASAP7_75t_SL g1671 ( 
.A(n_1657),
.B(n_1504),
.Y(n_1671)
);

INVx1_ASAP7_75t_SL g1672 ( 
.A(n_1666),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1639),
.B(n_1623),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1661),
.B(n_1623),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1644),
.B(n_1625),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1663),
.B(n_1612),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1632),
.A2(n_1593),
.B1(n_1542),
.B2(n_1568),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1629),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1648),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1663),
.B(n_1604),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1633),
.B(n_1610),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1629),
.Y(n_1682)
);

INVx4_ASAP7_75t_L g1683 ( 
.A(n_1631),
.Y(n_1683)
);

CKINVDCx16_ASAP7_75t_R g1684 ( 
.A(n_1635),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1631),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1648),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1633),
.B(n_1610),
.Y(n_1687)
);

NAND3x1_ASAP7_75t_SL g1688 ( 
.A(n_1653),
.B(n_1347),
.C(n_1568),
.Y(n_1688)
);

INVx3_ASAP7_75t_SL g1689 ( 
.A(n_1637),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1628),
.B(n_1618),
.Y(n_1690)
);

INVxp67_ASAP7_75t_L g1691 ( 
.A(n_1634),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1630),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1658),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1658),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1642),
.B(n_1618),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1664),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1646),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1642),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1651),
.B(n_1620),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1637),
.B(n_1593),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1650),
.B(n_1618),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1664),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1637),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1649),
.B(n_1620),
.Y(n_1704)
);

OAI21x1_ASAP7_75t_L g1705 ( 
.A1(n_1653),
.A2(n_1611),
.B(n_1601),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1645),
.B(n_1652),
.Y(n_1706)
);

INVx2_ASAP7_75t_SL g1707 ( 
.A(n_1689),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1689),
.B(n_1645),
.Y(n_1708)
);

NAND4xp75_ASAP7_75t_L g1709 ( 
.A(n_1674),
.B(n_1655),
.C(n_1662),
.D(n_1654),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1683),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1678),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1672),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1684),
.B(n_1655),
.Y(n_1713)
);

OAI21xp33_ASAP7_75t_L g1714 ( 
.A1(n_1690),
.A2(n_1670),
.B(n_1660),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1678),
.Y(n_1715)
);

NAND2xp33_ASAP7_75t_SL g1716 ( 
.A(n_1697),
.B(n_1654),
.Y(n_1716)
);

OAI21xp33_ASAP7_75t_L g1717 ( 
.A1(n_1701),
.A2(n_1670),
.B(n_1660),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1706),
.B(n_1665),
.Y(n_1718)
);

INVx2_ASAP7_75t_SL g1719 ( 
.A(n_1700),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1691),
.B(n_1652),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1703),
.B(n_1407),
.Y(n_1721)
);

OAI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1698),
.A2(n_1554),
.B1(n_1560),
.B2(n_1668),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1683),
.B(n_1669),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1676),
.B(n_1669),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1682),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1676),
.B(n_1685),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1682),
.Y(n_1727)
);

INVx1_ASAP7_75t_SL g1728 ( 
.A(n_1671),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1680),
.B(n_1662),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1692),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1683),
.Y(n_1731)
);

AOI21xp33_ASAP7_75t_SL g1732 ( 
.A1(n_1677),
.A2(n_1338),
.B(n_1570),
.Y(n_1732)
);

AOI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1728),
.A2(n_1671),
.B1(n_1700),
.B2(n_1698),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1723),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1731),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1719),
.B(n_1700),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1712),
.A2(n_1680),
.B1(n_1687),
.B2(n_1681),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1711),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1707),
.B(n_1681),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1721),
.B(n_1687),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1707),
.B(n_1695),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1715),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1725),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1719),
.B(n_1695),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1727),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1721),
.B(n_1699),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_SL g1747 ( 
.A(n_1716),
.B(n_1723),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1708),
.B(n_1675),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1730),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1716),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1710),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_R g1752 ( 
.A(n_1710),
.B(n_1343),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_SL g1753 ( 
.A(n_1750),
.B(n_1709),
.Y(n_1753)
);

A2O1A1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1747),
.A2(n_1732),
.B(n_1713),
.C(n_1726),
.Y(n_1754)
);

NAND3xp33_ASAP7_75t_L g1755 ( 
.A(n_1747),
.B(n_1713),
.C(n_1735),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1736),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1736),
.Y(n_1757)
);

AO21x1_ASAP7_75t_L g1758 ( 
.A1(n_1736),
.A2(n_1734),
.B(n_1751),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1733),
.B(n_1722),
.Y(n_1759)
);

OAI211xp5_ASAP7_75t_L g1760 ( 
.A1(n_1737),
.A2(n_1714),
.B(n_1717),
.C(n_1708),
.Y(n_1760)
);

OAI31xp33_ASAP7_75t_L g1761 ( 
.A1(n_1740),
.A2(n_1723),
.A3(n_1720),
.B(n_1724),
.Y(n_1761)
);

AOI21xp5_ASAP7_75t_SL g1762 ( 
.A1(n_1746),
.A2(n_1338),
.B(n_1387),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1737),
.A2(n_1597),
.B1(n_1718),
.B2(n_1729),
.Y(n_1763)
);

AOI221xp5_ASAP7_75t_L g1764 ( 
.A1(n_1739),
.A2(n_1729),
.B1(n_1692),
.B2(n_1686),
.C(n_1694),
.Y(n_1764)
);

AOI32xp33_ASAP7_75t_L g1765 ( 
.A1(n_1748),
.A2(n_1679),
.A3(n_1693),
.B1(n_1696),
.B2(n_1702),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1757),
.Y(n_1766)
);

NOR3xp33_ASAP7_75t_L g1767 ( 
.A(n_1755),
.B(n_1741),
.C(n_1734),
.Y(n_1767)
);

NAND4xp25_ASAP7_75t_L g1768 ( 
.A(n_1753),
.B(n_1744),
.C(n_1742),
.D(n_1743),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1762),
.B(n_1748),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1758),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1756),
.B(n_1752),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1761),
.B(n_1738),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1760),
.B(n_1745),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1759),
.B(n_1749),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1764),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1754),
.B(n_1752),
.Y(n_1776)
);

XNOR2x1_ASAP7_75t_SL g1777 ( 
.A(n_1765),
.B(n_1387),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_L g1778 ( 
.A(n_1770),
.B(n_1763),
.C(n_1699),
.Y(n_1778)
);

NAND3xp33_ASAP7_75t_L g1779 ( 
.A(n_1775),
.B(n_1675),
.C(n_1704),
.Y(n_1779)
);

OAI211xp5_ASAP7_75t_SL g1780 ( 
.A1(n_1773),
.A2(n_1343),
.B(n_1673),
.C(n_1383),
.Y(n_1780)
);

NAND2x1p5_ASAP7_75t_L g1781 ( 
.A(n_1771),
.B(n_1358),
.Y(n_1781)
);

NAND3xp33_ASAP7_75t_SL g1782 ( 
.A(n_1767),
.B(n_1704),
.C(n_1673),
.Y(n_1782)
);

NOR3xp33_ASAP7_75t_L g1783 ( 
.A(n_1768),
.B(n_1688),
.C(n_1705),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1779),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1782),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1778),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_SL g1787 ( 
.A1(n_1781),
.A2(n_1769),
.B1(n_1766),
.B2(n_1776),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1783),
.B(n_1774),
.Y(n_1788)
);

NOR2xp67_ASAP7_75t_L g1789 ( 
.A(n_1780),
.B(n_1768),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1781),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1787),
.B(n_1772),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1785),
.Y(n_1792)
);

AND4x2_ASAP7_75t_L g1793 ( 
.A(n_1789),
.B(n_1777),
.C(n_1788),
.D(n_1786),
.Y(n_1793)
);

AOI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1784),
.A2(n_1656),
.B1(n_1630),
.B2(n_1643),
.C(n_1636),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1790),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_SL g1796 ( 
.A(n_1788),
.B(n_1464),
.C(n_1688),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1795),
.B(n_1636),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1792),
.Y(n_1798)
);

INVxp33_ASAP7_75t_L g1799 ( 
.A(n_1791),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1797),
.Y(n_1800)
);

NAND4xp25_ASAP7_75t_L g1801 ( 
.A(n_1800),
.B(n_1798),
.C(n_1796),
.D(n_1793),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_SL g1802 ( 
.A1(n_1801),
.A2(n_1799),
.B1(n_1372),
.B2(n_1794),
.Y(n_1802)
);

AOI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1801),
.A2(n_1705),
.B1(n_1638),
.B2(n_1640),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1803),
.Y(n_1804)
);

OAI21x1_ASAP7_75t_L g1805 ( 
.A1(n_1802),
.A2(n_1667),
.B(n_1640),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1804),
.B(n_1649),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1804),
.A2(n_1805),
.B(n_1372),
.Y(n_1807)
);

OAI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1806),
.A2(n_1641),
.B(n_1638),
.Y(n_1808)
);

NAND3xp33_ASAP7_75t_L g1809 ( 
.A(n_1808),
.B(n_1807),
.C(n_1643),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1809),
.A2(n_1641),
.B1(n_1647),
.B2(n_1667),
.Y(n_1810)
);

AOI211xp5_ASAP7_75t_L g1811 ( 
.A1(n_1810),
.A2(n_1647),
.B(n_1659),
.C(n_1366),
.Y(n_1811)
);


endmodule