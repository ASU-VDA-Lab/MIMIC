module fake_jpeg_13116_n_316 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_17),
.B(n_6),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_62),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_8),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_46),
.B(n_69),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_29),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_50),
.B(n_59),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_33),
.B(n_13),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_56),
.Y(n_73)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_54),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_13),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_14),
.B(n_34),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_26),
.B(n_18),
.Y(n_101)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

CKINVDCx9p33_ASAP7_75t_R g68 ( 
.A(n_31),
.Y(n_68)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_27),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_11),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_70),
.B(n_9),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_80),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_68),
.A2(n_14),
.B1(n_34),
.B2(n_28),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_76),
.A2(n_87),
.B1(n_93),
.B2(n_106),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_35),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_83),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_40),
.A2(n_28),
.B1(n_23),
.B2(n_16),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_35),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_92),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_27),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_41),
.A2(n_22),
.B1(n_32),
.B2(n_31),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_97),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_40),
.B(n_27),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_109),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_113),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_102),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_44),
.B(n_26),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_59),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_51),
.A2(n_32),
.B1(n_18),
.B2(n_15),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_55),
.B(n_37),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_60),
.A2(n_23),
.B1(n_19),
.B2(n_37),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_111),
.A2(n_117),
.B1(n_118),
.B2(n_4),
.Y(n_163)
);

AND2x4_ASAP7_75t_SL g113 ( 
.A(n_47),
.B(n_37),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_115),
.Y(n_154)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_45),
.A2(n_19),
.B1(n_23),
.B2(n_37),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_54),
.A2(n_23),
.B1(n_19),
.B2(n_21),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_152),
.Y(n_166)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_108),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_127),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_78),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_112),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_142),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_99),
.A2(n_55),
.B1(n_19),
.B2(n_50),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

NAND2x1p5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_98),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_134),
.A2(n_147),
.B(n_71),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_135),
.Y(n_181)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_113),
.Y(n_139)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_143),
.B(n_155),
.Y(n_183)
);

AO22x1_ASAP7_75t_L g144 ( 
.A1(n_86),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_144),
.B(n_159),
.Y(n_168)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_146),
.A2(n_151),
.B1(n_162),
.B2(n_143),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_82),
.A2(n_76),
.B1(n_87),
.B2(n_103),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_93),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_151)
);

AO22x1_ASAP7_75t_SL g152 ( 
.A1(n_107),
.A2(n_3),
.B1(n_4),
.B2(n_9),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_161),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_74),
.B(n_10),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_95),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_75),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_158),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_77),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_3),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_72),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_3),
.B1(n_4),
.B2(n_94),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_136),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_104),
.B1(n_88),
.B2(n_89),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_194),
.B1(n_130),
.B2(n_161),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_154),
.B(n_89),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_173),
.B(n_184),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_120),
.B(n_104),
.C(n_71),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_153),
.C(n_123),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_79),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_81),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_185),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_193),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_137),
.A2(n_136),
.B1(n_148),
.B2(n_159),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_187),
.A2(n_188),
.B1(n_198),
.B2(n_130),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_136),
.A2(n_134),
.B1(n_163),
.B2(n_125),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_191),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_131),
.B(n_126),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_196),
.Y(n_220)
);

O2A1O1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_134),
.A2(n_147),
.B(n_144),
.C(n_152),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_186),
.B(n_185),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_132),
.B(n_125),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_144),
.A2(n_149),
.B1(n_121),
.B2(n_160),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_166),
.B(n_132),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_199),
.B(n_201),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_178),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_208),
.Y(n_239)
);

A2O1A1O1Ixp25_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_152),
.B(n_135),
.C(n_142),
.D(n_156),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_211),
.B1(n_177),
.B2(n_169),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_179),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_206),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_224),
.B1(n_225),
.B2(n_175),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_207),
.C(n_203),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_123),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_138),
.C(n_145),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_171),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_172),
.A2(n_140),
.B1(n_122),
.B2(n_129),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_187),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_216),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_217),
.B(n_176),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_167),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_222),
.B(n_226),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_165),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_185),
.A2(n_180),
.B(n_172),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_170),
.B(n_167),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_193),
.B1(n_183),
.B2(n_173),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_191),
.A2(n_182),
.B1(n_164),
.B2(n_174),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_181),
.A2(n_174),
.B(n_176),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_229),
.A2(n_242),
.B(n_220),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_234),
.B(n_218),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_235),
.A2(n_237),
.B1(n_227),
.B2(n_225),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_215),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_241),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_212),
.A2(n_169),
.B1(n_177),
.B2(n_189),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_175),
.B1(n_177),
.B2(n_189),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_250),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_197),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_218),
.A2(n_197),
.B1(n_224),
.B2(n_223),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_213),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_246),
.Y(n_266)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_215),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_248),
.C(n_207),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_216),
.C(n_214),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_251),
.A2(n_254),
.B1(n_255),
.B2(n_258),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_269),
.C(n_254),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_249),
.A2(n_218),
.B1(n_222),
.B2(n_223),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_217),
.B(n_226),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_256),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_206),
.B1(n_201),
.B2(n_199),
.Y(n_258)
);

AO22x1_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_202),
.B1(n_210),
.B2(n_208),
.Y(n_259)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_259),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_260),
.B(n_262),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_239),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_263),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_228),
.B(n_213),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_240),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_237),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_268),
.B1(n_244),
.B2(n_253),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_229),
.A2(n_231),
.B(n_234),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_238),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_230),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_247),
.B1(n_248),
.B2(n_232),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_269),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_262),
.B(n_228),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_277),
.Y(n_286)
);

NAND3xp33_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_245),
.C(n_232),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_273),
.B(n_266),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_255),
.B(n_251),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_264),
.A2(n_230),
.B1(n_233),
.B2(n_250),
.Y(n_275)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_233),
.Y(n_277)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_267),
.C(n_260),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_253),
.A2(n_263),
.B1(n_261),
.B2(n_259),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_274),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_288),
.C(n_289),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_285),
.A2(n_287),
.B1(n_283),
.B2(n_282),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_258),
.C(n_256),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_259),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_292),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_275),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_293),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_281),
.Y(n_296)
);

OAI21x1_ASAP7_75t_SL g304 ( 
.A1(n_296),
.A2(n_302),
.B(n_291),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_300),
.B(n_301),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_272),
.C(n_276),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_278),
.B1(n_272),
.B2(n_268),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_307),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_284),
.B(n_288),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_301),
.C(n_286),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_299),
.A2(n_265),
.B(n_285),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_309),
.B(n_286),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_295),
.C(n_298),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_303),
.B(n_296),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_312),
.C(n_302),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_265),
.B(n_257),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_271),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_257),
.Y(n_316)
);


endmodule