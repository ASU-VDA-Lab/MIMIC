module fake_jpeg_30325_n_371 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_371);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_371;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_SL g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_17),
.B(n_8),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_49),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_53),
.Y(n_97)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx6p67_ASAP7_75t_R g114 ( 
.A(n_52),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_56),
.B(n_59),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_27),
.B(n_8),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_69),
.Y(n_105)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_67),
.Y(n_99)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_0),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_27),
.B(n_31),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_75),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_24),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_21),
.B(n_36),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_82),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_81),
.Y(n_104)
);

BUFx2_ASAP7_75t_R g82 ( 
.A(n_31),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

HAxp5_ASAP7_75t_SL g89 ( 
.A(n_83),
.B(n_86),
.CON(n_89),
.SN(n_89)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_25),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_30),
.B1(n_44),
.B2(n_43),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_88),
.A2(n_91),
.B1(n_94),
.B2(n_118),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_30),
.B1(n_44),
.B2(n_43),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_23),
.B1(n_25),
.B2(n_39),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_93),
.A2(n_98),
.B1(n_102),
.B2(n_109),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_44),
.B1(n_30),
.B2(n_43),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_52),
.A2(n_23),
.B1(n_25),
.B2(n_32),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_60),
.A2(n_23),
.B1(n_32),
.B2(n_20),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_63),
.A2(n_32),
.B1(n_20),
.B2(n_29),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_63),
.A2(n_32),
.B1(n_20),
.B2(n_47),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_33),
.B1(n_36),
.B2(n_21),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_111),
.B(n_107),
.Y(n_180)
);

NAND2x1_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_20),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_115),
.B(n_129),
.Y(n_178)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_33),
.Y(n_117)
);

NOR2x1_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_9),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_65),
.A2(n_45),
.B1(n_41),
.B2(n_38),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_86),
.A2(n_32),
.B1(n_22),
.B2(n_29),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_61),
.B(n_45),
.C(n_41),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_69),
.C(n_9),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_54),
.A2(n_57),
.B1(n_58),
.B2(n_62),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_128),
.B1(n_83),
.B2(n_2),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_85),
.A2(n_38),
.B1(n_35),
.B2(n_26),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_77),
.A2(n_78),
.B1(n_84),
.B2(n_73),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_129),
.A2(n_89),
.B1(n_125),
.B2(n_114),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_66),
.A2(n_26),
.B1(n_35),
.B2(n_11),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_71),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_76),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_139),
.B(n_172),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_83),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_163),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_143),
.B(n_158),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_81),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_148),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_145),
.Y(n_211)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_96),
.B(n_15),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_81),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_150),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_87),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_87),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_162),
.Y(n_184)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_153),
.A2(n_171),
.B1(n_174),
.B2(n_92),
.Y(n_207)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx11_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_15),
.C(n_2),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_168),
.C(n_99),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_117),
.B(n_107),
.Y(n_158)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_95),
.B(n_15),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_106),
.B(n_1),
.Y(n_163)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_87),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_173),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_167),
.Y(n_195)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_115),
.B(n_1),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_126),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_100),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_101),
.B(n_4),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_128),
.A2(n_4),
.B1(n_5),
.B2(n_118),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_178),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_177),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_107),
.B(n_106),
.Y(n_177)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_113),
.Y(n_219)
);

OR2x2_ASAP7_75t_SL g203 ( 
.A(n_180),
.B(n_125),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_199),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_155),
.A2(n_111),
.B1(n_106),
.B2(n_138),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_193),
.A2(n_209),
.B1(n_179),
.B2(n_156),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_203),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_140),
.B(n_87),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_99),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_202),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_139),
.B(n_129),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_178),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_216),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_129),
.C(n_134),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_210),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_207),
.A2(n_208),
.B1(n_212),
.B2(n_214),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_164),
.A2(n_135),
.B1(n_133),
.B2(n_138),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_155),
.A2(n_132),
.B1(n_92),
.B2(n_127),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_104),
.C(n_103),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_153),
.A2(n_127),
.B1(n_89),
.B2(n_121),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_146),
.A2(n_133),
.B1(n_135),
.B2(n_116),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_116),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_112),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_169),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_182),
.B(n_143),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_226),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_172),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_243),
.C(n_210),
.Y(n_258)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

AO22x1_ASAP7_75t_L g224 ( 
.A1(n_197),
.A2(n_175),
.B1(n_203),
.B2(n_217),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_224),
.A2(n_249),
.B(n_189),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_176),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_230),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_175),
.C(n_141),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_229),
.B(n_216),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_176),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_186),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_231),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_184),
.B(n_182),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_235),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_175),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_234),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_146),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_170),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_218),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_207),
.A2(n_141),
.B1(n_142),
.B2(n_181),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_241),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_212),
.A2(n_181),
.B1(n_159),
.B2(n_171),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_197),
.A2(n_165),
.B(n_152),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_242),
.A2(n_209),
.B(n_215),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_192),
.B(n_154),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_197),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_244),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_195),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_247),
.A2(n_214),
.B1(n_199),
.B2(n_195),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_202),
.A2(n_160),
.B(n_113),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_250),
.Y(n_271)
);

AO21x1_ASAP7_75t_L g286 ( 
.A1(n_252),
.A2(n_239),
.B(n_249),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_253),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_206),
.B(n_192),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_257),
.A2(n_211),
.B(n_167),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_266),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_242),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_233),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_263),
.A2(n_211),
.B1(n_187),
.B2(n_220),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_272),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_227),
.B(n_198),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_246),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_275),
.C(n_277),
.Y(n_283)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_274),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_234),
.B(n_201),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_225),
.B(n_213),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_222),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_239),
.B(n_160),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_205),
.C(n_190),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_240),
.B(n_170),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_205),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_259),
.A2(n_224),
.B1(n_245),
.B2(n_247),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_279),
.A2(n_281),
.B1(n_284),
.B2(n_263),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_259),
.A2(n_229),
.B1(n_248),
.B2(n_237),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_240),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_282),
.B(n_289),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_264),
.A2(n_237),
.B1(n_238),
.B2(n_241),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_285),
.A2(n_257),
.B(n_258),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_297),
.B(n_252),
.Y(n_303)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_276),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_299),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_266),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_293),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_160),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_273),
.B(n_147),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_255),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_236),
.Y(n_295)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_295),
.Y(n_306)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_280),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_300),
.B(n_310),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_254),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_318),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_303),
.A2(n_298),
.B(n_285),
.Y(n_324)
);

NOR4xp25_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_262),
.C(n_261),
.D(n_274),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_278),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_308),
.A2(n_314),
.B1(n_298),
.B2(n_281),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_299),
.Y(n_310)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_313),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_284),
.A2(n_277),
.B1(n_253),
.B2(n_269),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_288),
.B(n_271),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_315),
.Y(n_323)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_316),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_278),
.B(n_283),
.C(n_293),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_318),
.C(n_312),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_290),
.B(n_275),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_320),
.B(n_324),
.Y(n_335)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_309),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_283),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_330),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_329),
.C(n_314),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_290),
.C(n_291),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_286),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_303),
.A2(n_319),
.B(n_311),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_332),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_338),
.B(n_341),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_311),
.C(n_308),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_339),
.B(n_342),
.C(n_331),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_333),
.A2(n_302),
.B1(n_313),
.B2(n_306),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_340),
.B(n_327),
.Y(n_348)
);

XNOR2x1_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_304),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_306),
.C(n_315),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_343),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_338),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_321),
.C(n_332),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_346),
.B(n_337),
.C(n_335),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_336),
.A2(n_334),
.B1(n_323),
.B2(n_325),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_347),
.A2(n_251),
.B1(n_270),
.B2(n_145),
.Y(n_356)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_348),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_343),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_350),
.B(n_200),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_342),
.A2(n_324),
.B(n_322),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_357),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_354),
.B(n_345),
.C(n_347),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_351),
.A2(n_341),
.B(n_335),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_356),
.A2(n_358),
.B1(n_161),
.B2(n_185),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_349),
.B(n_185),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_359),
.B(n_361),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_354),
.B(n_194),
.C(n_191),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_362),
.B(n_346),
.C(n_359),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_360),
.A2(n_352),
.B1(n_355),
.B2(n_194),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_364),
.B(n_365),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_365),
.B(n_363),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_366),
.B(n_363),
.Y(n_369)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_367),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_368),
.B(n_369),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_370),
.Y(n_371)
);


endmodule