module fake_jpeg_31288_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_5),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_4),
.B(n_3),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_17),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_22),
.Y(n_24)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_20),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_20),
.A2(n_12),
.B1(n_14),
.B2(n_10),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_23),
.A2(n_27),
.B1(n_15),
.B2(n_21),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_19),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_2),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_30),
.B(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_34),
.C(n_35),
.Y(n_38)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2x1_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_28),
.C(n_24),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_35),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_25),
.C(n_23),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_16),
.C(n_41),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_36),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_45),
.Y(n_47)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_16),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_49),
.A2(n_48),
.B(n_47),
.Y(n_50)
);


endmodule