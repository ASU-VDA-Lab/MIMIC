module fake_jpeg_7559_n_174 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_42),
.Y(n_64)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_19),
.B1(n_30),
.B2(n_32),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_47),
.A2(n_29),
.B1(n_62),
.B2(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_48),
.B(n_50),
.Y(n_79)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_53),
.Y(n_72)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_60),
.B(n_18),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_22),
.C(n_17),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_76),
.C(n_81),
.Y(n_96)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_78),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_26),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_77),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_25),
.B(n_23),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_21),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_23),
.Y(n_81)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_90),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_31),
.B(n_20),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_84),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_31),
.B(n_20),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_45),
.A2(n_30),
.B1(n_29),
.B2(n_18),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_88),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_45),
.A2(n_30),
.B1(n_29),
.B2(n_26),
.Y(n_87)
);

NAND2x1_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_61),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_15),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_92),
.A2(n_107),
.B1(n_109),
.B2(n_82),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_21),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_74),
.Y(n_112)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_115),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_120),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_66),
.B1(n_69),
.B2(n_68),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_118),
.B1(n_73),
.B2(n_72),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

NOR4xp25_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_67),
.C(n_77),
.D(n_78),
.Y(n_116)
);

NOR4xp25_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_91),
.C(n_107),
.D(n_92),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_106),
.B1(n_100),
.B2(n_101),
.Y(n_118)
);

XOR2x2_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_70),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_68),
.C(n_69),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_126),
.C(n_122),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_73),
.B(n_90),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_91),
.B(n_92),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_123),
.B(n_125),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_97),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_23),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_130),
.C(n_121),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_91),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_137),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_85),
.B1(n_56),
.B2(n_65),
.Y(n_148)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_109),
.B(n_98),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_135),
.Y(n_144)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_24),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_111),
.B1(n_110),
.B2(n_115),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_71),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_112),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_145),
.C(n_149),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_142),
.A2(n_148),
.B1(n_127),
.B2(n_139),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_126),
.Y(n_145)
);

BUFx12_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_146),
.B(n_147),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_113),
.C(n_71),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_25),
.B1(n_1),
.B2(n_3),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_130),
.C(n_132),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_154),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_133),
.C(n_134),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_134),
.C(n_24),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_156),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_56),
.C(n_23),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_143),
.B(n_144),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_157),
.A2(n_15),
.B1(n_23),
.B2(n_9),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_160),
.B(n_163),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_146),
.B1(n_85),
.B2(n_10),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_11),
.B1(n_10),
.B2(n_8),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_153),
.B(n_159),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_167),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_158),
.Y(n_170)
);

OAI221xp5_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_160),
.B1(n_158),
.B2(n_25),
.C(n_5),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_SL g171 ( 
.A1(n_168),
.A2(n_165),
.B(n_1),
.C(n_4),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_25),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_172),
.C(n_169),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_0),
.Y(n_174)
);


endmodule