module fake_jpeg_15994_n_190 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_18),
.B(n_1),
.Y(n_34)
);

CKINVDCx11_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_2),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_2),
.Y(n_38)
);

CKINVDCx12_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_2),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_46)
);

AO22x2_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_25),
.B1(n_21),
.B2(n_26),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_50),
.B1(n_19),
.B2(n_16),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_22),
.Y(n_69)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVxp33_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_21),
.B1(n_25),
.B2(n_29),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_61),
.Y(n_83)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_39),
.B(n_36),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_63),
.B(n_54),
.Y(n_81)
);

OR2x2_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_37),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_6),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_34),
.B1(n_28),
.B2(n_16),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_65),
.B1(n_69),
.B2(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_20),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_68),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_20),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_74),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_20),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_53),
.C(n_24),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_50),
.B1(n_4),
.B2(n_6),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_72),
.B(n_76),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_52),
.B(n_19),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_20),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_17),
.B1(n_23),
.B2(n_14),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_17),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_99),
.B(n_97),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_87),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_91),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_53),
.B1(n_44),
.B2(n_14),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_92),
.B1(n_71),
.B2(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_63),
.B(n_66),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_24),
.B1(n_40),
.B2(n_10),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_55),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_69),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_105),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_114),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_89),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_110),
.C(n_99),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_64),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_65),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_93),
.Y(n_137)
);

CKINVDCx10_ASAP7_75t_R g118 ( 
.A(n_80),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_118),
.Y(n_121)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_78),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_126),
.B(n_129),
.C(n_133),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_103),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_131),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_81),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_107),
.C(n_117),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_82),
.B1(n_88),
.B2(n_86),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_87),
.B1(n_99),
.B2(n_92),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_130),
.B(n_84),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_119),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_115),
.B1(n_105),
.B2(n_100),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_119),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_136),
.B(n_94),
.Y(n_151)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_150),
.C(n_125),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

OAI321xp33_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_109),
.A3(n_113),
.B1(n_77),
.B2(n_101),
.C(n_75),
.Y(n_141)
);

OA21x2_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_142),
.B(n_143),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_96),
.C(n_76),
.Y(n_142)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_122),
.B(n_112),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_128),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_144),
.B(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_122),
.B1(n_134),
.B2(n_133),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_152),
.A2(n_138),
.B1(n_130),
.B2(n_150),
.Y(n_165)
);

NOR2xp67_ASAP7_75t_SL g154 ( 
.A(n_142),
.B(n_147),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_SL g169 ( 
.A(n_154),
.B(n_156),
.C(n_7),
.Y(n_169)
);

AOI211xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_135),
.B(n_126),
.C(n_129),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_157),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_121),
.B1(n_108),
.B2(n_120),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_146),
.B1(n_120),
.B2(n_108),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_85),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_145),
.B(n_148),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_152),
.B(n_164),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_165),
.B(n_170),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_169),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_162),
.C(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_9),
.Y(n_168)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_10),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_156),
.B1(n_153),
.B2(n_155),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_174),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_176),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_160),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_181),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_174),
.A2(n_159),
.B1(n_175),
.B2(n_176),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_182),
.A2(n_159),
.B(n_167),
.Y(n_183)
);

MAJx2_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_182),
.C(n_178),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_187),
.B(n_185),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_184),
.A2(n_11),
.B(n_12),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_7),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_7),
.Y(n_190)
);


endmodule