module fake_jpeg_6093_n_307 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_23),
.B(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_41),
.Y(n_48)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_17),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_27),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_20),
.B1(n_31),
.B2(n_23),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_45),
.A2(n_47),
.B1(n_22),
.B2(n_24),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_42),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_20),
.B1(n_31),
.B2(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_27),
.B1(n_31),
.B2(n_33),
.Y(n_56)
);

AO22x1_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_27),
.B1(n_39),
.B2(n_35),
.Y(n_77)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_63),
.Y(n_71)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_59),
.Y(n_75)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_27),
.Y(n_72)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_20),
.B1(n_31),
.B2(n_18),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_16),
.B1(n_30),
.B2(n_22),
.Y(n_89)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_72),
.B(n_90),
.Y(n_111)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_78),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_56),
.B1(n_59),
.B2(n_62),
.Y(n_94)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_20),
.B1(n_29),
.B2(n_28),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_21),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_28),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_56),
.B1(n_61),
.B2(n_40),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_55),
.B(n_29),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_28),
.Y(n_103)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_29),
.B(n_30),
.C(n_16),
.Y(n_90)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_92),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_106),
.B1(n_118),
.B2(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_95),
.B(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_103),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_107),
.B1(n_114),
.B2(n_54),
.Y(n_121)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_44),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_65),
.B1(n_56),
.B2(n_64),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_112),
.Y(n_125)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

BUFx4f_ASAP7_75t_SL g142 ( 
.A(n_109),
.Y(n_142)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_82),
.B(n_61),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_77),
.A2(n_67),
.B1(n_37),
.B2(n_57),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_48),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_27),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_71),
.Y(n_116)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_72),
.A2(n_50),
.B(n_37),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_73),
.B(n_49),
.C(n_75),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_72),
.A2(n_37),
.B1(n_41),
.B2(n_40),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_137),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_133),
.B1(n_107),
.B2(n_95),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_132),
.B1(n_140),
.B2(n_141),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_75),
.C(n_93),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_143),
.C(n_98),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_75),
.B1(n_53),
.B2(n_92),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_105),
.B(n_104),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_49),
.B(n_68),
.C(n_30),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_135),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_101),
.A2(n_40),
.B1(n_41),
.B2(n_93),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_96),
.A2(n_79),
.B1(n_70),
.B2(n_91),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_136),
.B1(n_139),
.B2(n_25),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_68),
.B(n_16),
.C(n_79),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_70),
.B1(n_91),
.B2(n_84),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_105),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_138),
.B(n_118),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_84),
.B1(n_88),
.B2(n_78),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_41),
.B1(n_40),
.B2(n_88),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_41),
.B1(n_88),
.B2(n_74),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_39),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_144),
.B(n_94),
.Y(n_155)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_157),
.B1(n_127),
.B2(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_148),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_129),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_150),
.B(n_151),
.Y(n_184)
);

NAND2x1_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_115),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_125),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_156),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_97),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_33),
.Y(n_194)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_116),
.C(n_112),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_159),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_150),
.C(n_169),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_103),
.B1(n_108),
.B2(n_110),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_99),
.Y(n_162)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_129),
.A2(n_99),
.B(n_98),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_169),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_26),
.B1(n_21),
.B2(n_18),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_26),
.B1(n_21),
.B2(n_18),
.Y(n_166)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_126),
.A2(n_39),
.B(n_35),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_170),
.A2(n_171),
.B1(n_123),
.B2(n_142),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_123),
.A2(n_25),
.B1(n_24),
.B2(n_26),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_173),
.A2(n_181),
.B1(n_185),
.B2(n_189),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_177),
.C(n_190),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_127),
.C(n_133),
.Y(n_177)
);

A2O1A1O1Ixp25_ASAP7_75t_L g178 ( 
.A1(n_151),
.A2(n_120),
.B(n_135),
.C(n_131),
.D(n_122),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_178),
.B(n_194),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_137),
.B1(n_136),
.B2(n_122),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_182),
.A2(n_186),
.B1(n_192),
.B2(n_168),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_128),
.B1(n_123),
.B2(n_142),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_142),
.B1(n_39),
.B2(n_35),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_142),
.B1(n_35),
.B2(n_119),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_32),
.C(n_33),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_32),
.B1(n_33),
.B2(n_2),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_146),
.A2(n_32),
.B1(n_33),
.B2(n_2),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_152),
.B1(n_155),
.B2(n_167),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_197),
.A2(n_208),
.B1(n_181),
.B2(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_199),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_152),
.B(n_148),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_206),
.B(n_214),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_195),
.A2(n_147),
.B1(n_156),
.B2(n_149),
.Y(n_203)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_158),
.C(n_162),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_212),
.C(n_213),
.Y(n_229)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_216),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_164),
.B(n_153),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_158),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_209),
.Y(n_222)
);

AO22x2_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_149),
.B1(n_165),
.B2(n_166),
.Y(n_208)
);

NAND2x1_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_32),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_174),
.B(n_145),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_15),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_217),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_15),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_0),
.C(n_1),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_187),
.B(n_195),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_14),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_194),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_12),
.Y(n_220)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_176),
.Y(n_224)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_172),
.Y(n_225)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_216),
.A2(n_172),
.B1(n_188),
.B2(n_178),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_226),
.A2(n_237),
.B1(n_200),
.B2(n_208),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_228),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_194),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_236),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_11),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_208),
.A2(n_0),
.B(n_1),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_208),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_219),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_0),
.C(n_2),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_213),
.C(n_212),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_246),
.C(n_250),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_242),
.A2(n_236),
.B(n_233),
.Y(n_265)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_204),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_224),
.A2(n_215),
.B1(n_209),
.B2(n_202),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_253),
.B1(n_223),
.B2(n_226),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_222),
.C(n_240),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_211),
.C(n_2),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_255),
.C(n_239),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_225),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_230),
.B(n_11),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_254),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_10),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_245),
.A2(n_231),
.B1(n_221),
.B2(n_238),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_260),
.A2(n_262),
.B1(n_241),
.B2(n_255),
.Y(n_272)
);

AOI21x1_ASAP7_75t_SL g261 ( 
.A1(n_243),
.A2(n_237),
.B(n_230),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_265),
.B(n_252),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_248),
.B1(n_232),
.B2(n_250),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_264),
.C(n_266),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_233),
.C(n_4),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_10),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_268),
.B(n_3),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_275),
.B(n_276),
.Y(n_286)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_278),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_244),
.C(n_246),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_267),
.B(n_244),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_277),
.B(n_258),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_259),
.A2(n_3),
.B(n_4),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_280),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_265),
.B(n_269),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_275),
.A2(n_264),
.B1(n_269),
.B2(n_266),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_5),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_282),
.Y(n_292)
);

NOR2xp67_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_263),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_5),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_271),
.B(n_3),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_288),
.A2(n_5),
.B(n_6),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_273),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_289),
.B(n_6),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_5),
.Y(n_290)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);

AOI21xp33_ASAP7_75t_L g297 ( 
.A1(n_293),
.A2(n_296),
.B(n_6),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_8),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_7),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_299),
.Y(n_301)
);

A2O1A1O1Ixp25_ASAP7_75t_L g303 ( 
.A1(n_301),
.A2(n_302),
.B(n_298),
.C(n_291),
.D(n_286),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_283),
.Y(n_304)
);

OAI21x1_ASAP7_75t_SL g305 ( 
.A1(n_304),
.A2(n_300),
.B(n_7),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_305),
.A2(n_7),
.B(n_8),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_8),
.Y(n_307)
);


endmodule