module fake_jpeg_14655_n_94 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_94);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_94;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx3_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_1),
.B(n_3),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_31),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_1),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_22),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_22),
.B1(n_13),
.B2(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2x1_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_24),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_43),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_47),
.B1(n_48),
.B2(n_20),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_24),
.B(n_21),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_19),
.B(n_14),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_30),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_2),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_26),
.A2(n_13),
.B1(n_16),
.B2(n_15),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_26),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_23),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_23),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_18),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_50),
.B(n_56),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_45),
.B(n_40),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_16),
.B1(n_33),
.B2(n_4),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_62),
.B1(n_3),
.B2(n_4),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_59),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_28),
.C(n_20),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_63),
.B(n_42),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_72),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_71),
.B1(n_20),
.B2(n_28),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_41),
.B(n_35),
.C(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_52),
.B1(n_57),
.B2(n_61),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_74),
.B1(n_78),
.B2(n_79),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_50),
.C(n_53),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_76),
.C(n_77),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_35),
.C(n_52),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_28),
.C(n_37),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_46),
.B1(n_51),
.B2(n_56),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_67),
.C(n_68),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_71),
.C(n_9),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_85),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_71),
.C(n_8),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_88),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_4),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_10),
.C(n_11),
.Y(n_91)
);

BUFx24_ASAP7_75t_SL g92 ( 
.A(n_91),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_86),
.C(n_90),
.Y(n_93)
);

AOI322xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_6),
.A3(n_86),
.B1(n_89),
.B2(n_92),
.C1(n_90),
.C2(n_88),
.Y(n_94)
);


endmodule