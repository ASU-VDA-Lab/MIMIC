module fake_jpeg_19589_n_23 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_23);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_23;

wire n_13;
wire n_21;
wire n_10;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

BUFx3_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

OA22x2_ASAP7_75t_L g11 ( 
.A1(n_3),
.A2(n_9),
.B1(n_0),
.B2(n_7),
.Y(n_11)
);

NAND2xp33_ASAP7_75t_SL g12 ( 
.A(n_2),
.B(n_6),
.Y(n_12)
);

OAI22xp33_ASAP7_75t_L g13 ( 
.A1(n_8),
.A2(n_5),
.B1(n_3),
.B2(n_1),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_1),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_14),
.A2(n_2),
.B(n_4),
.Y(n_17)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

OAI21xp33_ASAP7_75t_SL g18 ( 
.A1(n_15),
.A2(n_16),
.B(n_11),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_12),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_18),
.C(n_11),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_18),
.B(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_20),
.Y(n_21)
);

AOI322xp5_ASAP7_75t_L g22 ( 
.A1(n_21),
.A2(n_13),
.A3(n_11),
.B1(n_16),
.B2(n_15),
.C1(n_4),
.C2(n_5),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_11),
.Y(n_23)
);


endmodule