module real_aes_878_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_552;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AO22x2_ASAP7_75t_L g99 ( .A1(n_0), .A2(n_56), .B1(n_89), .B2(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g161 ( .A(n_1), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_2), .B(n_188), .Y(n_211) );
AOI22xp33_ASAP7_75t_SL g109 ( .A1(n_3), .A2(n_68), .B1(n_110), .B2(n_113), .Y(n_109) );
INVx1_ASAP7_75t_L g233 ( .A(n_4), .Y(n_233) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_5), .A2(n_18), .B1(n_89), .B2(n_97), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_6), .Y(n_249) );
AOI22xp33_ASAP7_75t_SL g539 ( .A1(n_6), .A2(n_80), .B1(n_81), .B2(n_249), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g142 ( .A1(n_7), .A2(n_143), .B1(n_144), .B2(n_147), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_7), .Y(n_143) );
INVx2_ASAP7_75t_L g187 ( .A(n_8), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g136 ( .A1(n_9), .A2(n_11), .B1(n_137), .B2(n_138), .Y(n_136) );
INVx1_ASAP7_75t_L g221 ( .A(n_10), .Y(n_221) );
INVx1_ASAP7_75t_L g218 ( .A(n_12), .Y(n_218) );
INVx1_ASAP7_75t_SL g293 ( .A(n_13), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_14), .B(n_198), .Y(n_197) );
AOI33xp33_ASAP7_75t_L g270 ( .A1(n_15), .A2(n_38), .A3(n_178), .B1(n_193), .B2(n_271), .B3(n_272), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_16), .A2(n_67), .B1(n_145), .B2(n_146), .Y(n_144) );
INVx1_ASAP7_75t_L g146 ( .A(n_16), .Y(n_146) );
INVx1_ASAP7_75t_L g242 ( .A(n_17), .Y(n_242) );
OAI221xp5_ASAP7_75t_L g153 ( .A1(n_18), .A2(n_56), .B1(n_58), .B2(n_154), .C(n_156), .Y(n_153) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_19), .A2(n_70), .B(n_187), .Y(n_186) );
OR2x2_ASAP7_75t_L g189 ( .A(n_19), .B(n_70), .Y(n_189) );
AOI22xp33_ASAP7_75t_SL g124 ( .A1(n_20), .A2(n_66), .B1(n_125), .B2(n_126), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_21), .B(n_231), .Y(n_290) );
INVx3_ASAP7_75t_L g89 ( .A(n_22), .Y(n_89) );
AO222x2_ASAP7_75t_L g84 ( .A1(n_23), .A2(n_41), .B1(n_50), .B2(n_85), .C1(n_101), .C2(n_104), .Y(n_84) );
AOI22xp33_ASAP7_75t_L g115 ( .A1(n_24), .A2(n_44), .B1(n_116), .B2(n_119), .Y(n_115) );
INVx1_ASAP7_75t_SL g90 ( .A(n_25), .Y(n_90) );
INVx1_ASAP7_75t_L g163 ( .A(n_26), .Y(n_163) );
AND2x2_ASAP7_75t_L g182 ( .A(n_26), .B(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g207 ( .A(n_26), .B(n_161), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_27), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_28), .B(n_231), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_29), .A2(n_69), .B1(n_134), .B2(n_135), .Y(n_133) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_30), .A2(n_175), .B1(n_185), .B2(n_188), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_31), .B(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_32), .B(n_198), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_33), .A2(n_80), .B1(n_81), .B2(n_548), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_33), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_34), .B(n_209), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_35), .B(n_198), .Y(n_234) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_36), .A2(n_58), .B1(n_89), .B2(n_93), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_37), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_39), .B(n_198), .Y(n_261) );
INVx1_ASAP7_75t_L g179 ( .A(n_40), .Y(n_179) );
INVx1_ASAP7_75t_L g200 ( .A(n_40), .Y(n_200) );
AND2x2_ASAP7_75t_L g262 ( .A(n_42), .B(n_263), .Y(n_262) );
AOI221xp5_ASAP7_75t_L g230 ( .A1(n_43), .A2(n_60), .B1(n_191), .B2(n_231), .C(n_232), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_45), .B(n_231), .Y(n_285) );
INVx1_ASAP7_75t_L g91 ( .A(n_46), .Y(n_91) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_47), .A2(n_53), .B1(n_129), .B2(n_131), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_48), .B(n_185), .Y(n_251) );
AOI21xp5_ASAP7_75t_SL g281 ( .A1(n_49), .A2(n_191), .B(n_282), .Y(n_281) );
AOI22xp33_ASAP7_75t_SL g79 ( .A1(n_51), .A2(n_80), .B1(n_81), .B2(n_139), .Y(n_79) );
INVx1_ASAP7_75t_L g139 ( .A(n_51), .Y(n_139) );
INVx1_ASAP7_75t_L g214 ( .A(n_52), .Y(n_214) );
INVx1_ASAP7_75t_L g260 ( .A(n_54), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_55), .A2(n_191), .B(n_259), .Y(n_258) );
INVxp33_ASAP7_75t_L g158 ( .A(n_56), .Y(n_158) );
INVx1_ASAP7_75t_L g183 ( .A(n_57), .Y(n_183) );
INVx1_ASAP7_75t_L g202 ( .A(n_57), .Y(n_202) );
INVxp67_ASAP7_75t_L g157 ( .A(n_58), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_59), .B(n_231), .Y(n_273) );
AND2x2_ASAP7_75t_L g295 ( .A(n_61), .B(n_238), .Y(n_295) );
INVx1_ASAP7_75t_L g215 ( .A(n_62), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_63), .A2(n_191), .B(n_292), .Y(n_291) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_64), .A2(n_191), .B(n_196), .C(n_208), .Y(n_190) );
AND2x2_ASAP7_75t_SL g279 ( .A(n_65), .B(n_238), .Y(n_279) );
INVx1_ASAP7_75t_L g145 ( .A(n_67), .Y(n_145) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_67), .A2(n_191), .B1(n_268), .B2(n_269), .Y(n_267) );
INVx1_ASAP7_75t_L g283 ( .A(n_71), .Y(n_283) );
AND2x2_ASAP7_75t_L g274 ( .A(n_72), .B(n_238), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_73), .A2(n_240), .B(n_241), .C(n_243), .Y(n_239) );
INVx1_ASAP7_75t_L g555 ( .A(n_73), .Y(n_555) );
INVx1_ASAP7_75t_L g148 ( .A(n_74), .Y(n_148) );
BUFx2_ASAP7_75t_SL g155 ( .A(n_75), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_76), .B(n_198), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_150), .B1(n_164), .B2(n_535), .C(n_538), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_140), .Y(n_78) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_81), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
AND2x2_ASAP7_75t_L g82 ( .A(n_83), .B(n_122), .Y(n_82) );
NOR2xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_108), .Y(n_83) );
AND2x4_ASAP7_75t_L g85 ( .A(n_86), .B(n_94), .Y(n_85) );
AND2x2_ASAP7_75t_L g113 ( .A(n_86), .B(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g119 ( .A(n_86), .B(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_92), .Y(n_86) );
HB1xp67_ASAP7_75t_L g102 ( .A(n_87), .Y(n_102) );
AND2x2_ASAP7_75t_L g106 ( .A(n_87), .B(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g112 ( .A(n_87), .Y(n_112) );
OAI22x1_ASAP7_75t_L g87 ( .A1(n_88), .A2(n_89), .B1(n_90), .B2(n_91), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g93 ( .A(n_89), .Y(n_93) );
INVx2_ASAP7_75t_L g97 ( .A(n_89), .Y(n_97) );
INVx1_ASAP7_75t_L g100 ( .A(n_89), .Y(n_100) );
INVx2_ASAP7_75t_L g107 ( .A(n_92), .Y(n_107) );
AND2x2_ASAP7_75t_L g111 ( .A(n_92), .B(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g127 ( .A(n_92), .Y(n_127) );
AND2x2_ASAP7_75t_L g129 ( .A(n_94), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g134 ( .A(n_94), .B(n_106), .Y(n_134) );
AND2x6_ASAP7_75t_L g137 ( .A(n_94), .B(n_111), .Y(n_137) );
AND2x4_ASAP7_75t_L g94 ( .A(n_95), .B(n_98), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
AND2x2_ASAP7_75t_L g103 ( .A(n_96), .B(n_99), .Y(n_103) );
AND2x4_ASAP7_75t_L g105 ( .A(n_96), .B(n_98), .Y(n_105) );
INVx1_ASAP7_75t_L g118 ( .A(n_96), .Y(n_118) );
INVxp67_ASAP7_75t_L g114 ( .A(n_98), .Y(n_114) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x2_ASAP7_75t_L g117 ( .A(n_99), .B(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_SL g101 ( .A(n_102), .B(n_103), .Y(n_101) );
AND2x4_ASAP7_75t_L g126 ( .A(n_103), .B(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g135 ( .A(n_103), .B(n_130), .Y(n_135) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
AND2x2_ASAP7_75t_L g110 ( .A(n_105), .B(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g131 ( .A(n_105), .B(n_130), .Y(n_131) );
AND2x4_ASAP7_75t_L g116 ( .A(n_106), .B(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g130 ( .A(n_107), .B(n_112), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_115), .Y(n_108) );
AND2x2_ASAP7_75t_SL g125 ( .A(n_111), .B(n_117), .Y(n_125) );
AND2x6_ASAP7_75t_L g138 ( .A(n_117), .B(n_130), .Y(n_138) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_118), .Y(n_121) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_132), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_128), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_136), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g140 ( .A1(n_141), .A2(n_142), .B1(n_148), .B2(n_149), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g147 ( .A(n_144), .Y(n_147) );
INVx1_ASAP7_75t_L g149 ( .A(n_148), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_151), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_152), .Y(n_151) );
AND3x1_ASAP7_75t_SL g152 ( .A(n_153), .B(n_159), .C(n_162), .Y(n_152) );
INVxp67_ASAP7_75t_L g545 ( .A(n_153), .Y(n_545) );
CKINVDCx8_ASAP7_75t_R g154 ( .A(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
CKINVDCx16_ASAP7_75t_R g543 ( .A(n_159), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_159), .A2(n_176), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g177 ( .A(n_160), .B(n_178), .Y(n_177) );
OR2x2_ASAP7_75t_SL g551 ( .A(n_160), .B(n_162), .Y(n_551) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g195 ( .A(n_161), .B(n_179), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_162), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2x1p5_ASAP7_75t_L g192 ( .A(n_163), .B(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_469), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_392), .Y(n_167) );
NAND3xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_339), .C(n_372), .Y(n_168) );
AOI211xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_296), .B(n_305), .C(n_329), .Y(n_169) );
OAI21xp33_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_225), .B(n_275), .Y(n_170) );
OR2x2_ASAP7_75t_L g349 ( .A(n_171), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g504 ( .A(n_171), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI22xp33_ASAP7_75t_SL g394 ( .A1(n_172), .A2(n_395), .B1(n_399), .B2(n_401), .Y(n_394) );
AND2x2_ASAP7_75t_L g431 ( .A(n_172), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_210), .Y(n_172) );
INVx1_ASAP7_75t_L g328 ( .A(n_173), .Y(n_328) );
AND2x4_ASAP7_75t_L g345 ( .A(n_173), .B(n_326), .Y(n_345) );
INVx2_ASAP7_75t_L g367 ( .A(n_173), .Y(n_367) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_173), .Y(n_450) );
AND2x2_ASAP7_75t_L g521 ( .A(n_173), .B(n_278), .Y(n_521) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_190), .Y(n_173) );
NOR3xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_180), .C(n_184), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x4_ASAP7_75t_L g231 ( .A(n_177), .B(n_181), .Y(n_231) );
OR2x6_ASAP7_75t_L g205 ( .A(n_178), .B(n_194), .Y(n_205) );
INVxp33_ASAP7_75t_L g271 ( .A(n_178), .Y(n_271) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x4_ASAP7_75t_L g223 ( .A(n_179), .B(n_201), .Y(n_223) );
INVxp67_ASAP7_75t_L g554 ( .A(n_180), .Y(n_554) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x6_ASAP7_75t_L g537 ( .A(n_182), .B(n_195), .Y(n_537) );
INVx2_ASAP7_75t_L g194 ( .A(n_183), .Y(n_194) );
AND2x6_ASAP7_75t_L g220 ( .A(n_183), .B(n_199), .Y(n_220) );
INVx4_ASAP7_75t_L g238 ( .A(n_185), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_185), .B(n_248), .Y(n_247) );
INVx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
BUFx4f_ASAP7_75t_L g209 ( .A(n_186), .Y(n_209) );
AND2x4_ASAP7_75t_L g188 ( .A(n_187), .B(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_SL g264 ( .A(n_187), .B(n_189), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_188), .B(n_206), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_188), .A2(n_281), .B(n_285), .Y(n_280) );
INVxp67_ASAP7_75t_L g250 ( .A(n_191), .Y(n_250) );
AND2x4_ASAP7_75t_L g191 ( .A(n_192), .B(n_195), .Y(n_191) );
INVx1_ASAP7_75t_L g272 ( .A(n_193), .Y(n_272) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_203), .B(n_206), .Y(n_196) );
INVx1_ASAP7_75t_L g216 ( .A(n_198), .Y(n_216) );
AND2x4_ASAP7_75t_L g198 ( .A(n_199), .B(n_201), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_205), .A2(n_214), .B1(n_215), .B2(n_216), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_SL g232 ( .A1(n_205), .A2(n_206), .B(n_233), .C(n_234), .Y(n_232) );
INVxp67_ASAP7_75t_L g240 ( .A(n_205), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_205), .A2(n_206), .B(n_260), .C(n_261), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g282 ( .A1(n_205), .A2(n_206), .B(n_283), .C(n_284), .Y(n_282) );
O2A1O1Ixp33_ASAP7_75t_SL g292 ( .A1(n_205), .A2(n_206), .B(n_293), .C(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g268 ( .A(n_206), .Y(n_268) );
INVx5_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_207), .Y(n_243) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_208), .A2(n_266), .B(n_274), .Y(n_265) );
AO21x2_ASAP7_75t_L g310 ( .A1(n_208), .A2(n_266), .B(n_274), .Y(n_310) );
INVx2_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_209), .A2(n_230), .B(n_235), .Y(n_229) );
AND2x2_ASAP7_75t_L g286 ( .A(n_210), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g315 ( .A(n_210), .Y(n_315) );
INVx3_ASAP7_75t_L g326 ( .A(n_210), .Y(n_326) );
AND2x4_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_217), .B(n_224), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_216), .B(n_242), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B1(n_221), .B2(n_222), .Y(n_217) );
INVxp67_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVxp67_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_225), .A2(n_516), .B1(n_518), .B2(n_520), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_225), .B(n_527), .Y(n_526) );
INVx2_ASAP7_75t_SL g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_253), .Y(n_226) );
INVx3_ASAP7_75t_L g299 ( .A(n_227), .Y(n_299) );
AND2x2_ASAP7_75t_L g307 ( .A(n_227), .B(n_308), .Y(n_307) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_227), .Y(n_337) );
NAND2x1_ASAP7_75t_SL g531 ( .A(n_227), .B(n_298), .Y(n_531) );
AND2x4_ASAP7_75t_L g227 ( .A(n_228), .B(n_236), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g304 ( .A(n_229), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_229), .B(n_310), .Y(n_322) );
AND2x2_ASAP7_75t_L g335 ( .A(n_229), .B(n_236), .Y(n_335) );
AND2x4_ASAP7_75t_L g342 ( .A(n_229), .B(n_343), .Y(n_342) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_229), .Y(n_391) );
INVxp67_ASAP7_75t_L g398 ( .A(n_229), .Y(n_398) );
INVx1_ASAP7_75t_L g403 ( .A(n_229), .Y(n_403) );
INVx1_ASAP7_75t_L g252 ( .A(n_231), .Y(n_252) );
INVx1_ASAP7_75t_L g302 ( .A(n_236), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_236), .B(n_312), .Y(n_321) );
INVx2_ASAP7_75t_L g389 ( .A(n_236), .Y(n_389) );
INVx1_ASAP7_75t_L g428 ( .A(n_236), .Y(n_428) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_246), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B1(n_244), .B2(n_245), .Y(n_237) );
INVx3_ASAP7_75t_L g245 ( .A(n_238), .Y(n_245) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_245), .A2(n_256), .B(n_262), .Y(n_255) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_245), .A2(n_256), .B(n_262), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_250), .B1(n_251), .B2(n_252), .Y(n_246) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g358 ( .A(n_253), .B(n_335), .Y(n_358) );
AND2x2_ASAP7_75t_L g426 ( .A(n_253), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g440 ( .A(n_253), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_253), .B(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_L g253 ( .A(n_254), .B(n_265), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2x1_ASAP7_75t_L g303 ( .A(n_255), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g396 ( .A(n_255), .B(n_389), .Y(n_396) );
AND2x2_ASAP7_75t_L g487 ( .A(n_255), .B(n_309), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_263), .Y(n_288) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g298 ( .A(n_265), .Y(n_298) );
INVx2_ASAP7_75t_L g343 ( .A(n_265), .Y(n_343) );
AND2x2_ASAP7_75t_L g388 ( .A(n_265), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_267), .B(n_273), .Y(n_266) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_286), .Y(n_276) );
AND2x2_ASAP7_75t_L g430 ( .A(n_277), .B(n_431), .Y(n_430) );
OR2x6_ASAP7_75t_L g489 ( .A(n_277), .B(n_490), .Y(n_489) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx4_ASAP7_75t_L g319 ( .A(n_278), .Y(n_319) );
AND2x4_ASAP7_75t_L g327 ( .A(n_278), .B(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g362 ( .A(n_278), .B(n_287), .Y(n_362) );
INVx2_ASAP7_75t_L g411 ( .A(n_278), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_278), .B(n_385), .Y(n_460) );
AND2x2_ASAP7_75t_L g497 ( .A(n_278), .B(n_315), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_278), .B(n_380), .Y(n_505) );
OR2x6_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g338 ( .A(n_286), .B(n_327), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_286), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_SL g477 ( .A(n_286), .B(n_365), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_286), .B(n_378), .Y(n_499) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_287), .Y(n_317) );
AND2x2_ASAP7_75t_L g325 ( .A(n_287), .B(n_326), .Y(n_325) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_287), .Y(n_348) );
INVx2_ASAP7_75t_L g351 ( .A(n_287), .Y(n_351) );
INVx1_ASAP7_75t_L g384 ( .A(n_287), .Y(n_384) );
INVx1_ASAP7_75t_L g432 ( .A(n_287), .Y(n_432) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_289), .B(n_295), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
NAND2xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_300), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_298), .B(n_301), .Y(n_374) );
OR2x2_ASAP7_75t_L g446 ( .A(n_298), .B(n_447), .Y(n_446) );
AND4x1_ASAP7_75t_SL g492 ( .A(n_298), .B(n_474), .C(n_493), .D(n_494), .Y(n_492) );
OR2x2_ASAP7_75t_L g516 ( .A(n_299), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AND2x2_ASAP7_75t_L g353 ( .A(n_302), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_302), .B(n_311), .Y(n_503) );
AND2x2_ASAP7_75t_L g528 ( .A(n_303), .B(n_388), .Y(n_528) );
OAI32xp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_313), .A3(n_318), .B1(n_320), .B2(n_323), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g401 ( .A(n_308), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g501 ( .A(n_308), .B(n_455), .Y(n_501) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
AND2x2_ASAP7_75t_L g397 ( .A(n_309), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g483 ( .A(n_309), .Y(n_483) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_310), .B(n_312), .Y(n_517) );
INVx3_ASAP7_75t_L g334 ( .A(n_311), .Y(n_334) );
NAND2x1p5_ASAP7_75t_L g512 ( .A(n_311), .B(n_439), .Y(n_512) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_312), .Y(n_371) );
AND2x2_ASAP7_75t_L g390 ( .A(n_312), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g524 ( .A(n_314), .Y(n_524) );
NAND2x1_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g364 ( .A(n_315), .Y(n_364) );
NOR2x1_ASAP7_75t_L g465 ( .A(n_315), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_318), .B(n_424), .Y(n_423) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g356 ( .A(n_319), .B(n_324), .Y(n_356) );
AND2x4_ASAP7_75t_L g378 ( .A(n_319), .B(n_328), .Y(n_378) );
AND2x4_ASAP7_75t_SL g449 ( .A(n_319), .B(n_450), .Y(n_449) );
NOR2x1_ASAP7_75t_L g475 ( .A(n_319), .B(n_400), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_320), .A2(n_443), .B1(n_446), .B2(n_448), .Y(n_442) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx2_ASAP7_75t_SL g462 ( .A(n_321), .Y(n_462) );
INVx2_ASAP7_75t_L g354 ( .A(n_322), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_325), .B(n_331), .Y(n_330) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_325), .A2(n_461), .B1(n_464), .B2(n_467), .Y(n_463) );
INVx1_ASAP7_75t_L g385 ( .A(n_326), .Y(n_385) );
AND2x2_ASAP7_75t_L g408 ( .A(n_326), .B(n_367), .Y(n_408) );
INVx2_ASAP7_75t_L g331 ( .A(n_327), .Y(n_331) );
OAI21xp5_ASAP7_75t_SL g329 ( .A1(n_330), .A2(n_332), .B(n_336), .Y(n_329) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_333), .A2(n_405), .B1(n_409), .B2(n_410), .Y(n_404) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_334), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_334), .B(n_402), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_334), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NOR3xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_355), .C(n_359), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_344), .B1(n_349), .B2(n_352), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g369 ( .A(n_342), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g409 ( .A(n_342), .B(n_396), .Y(n_409) );
AND2x2_ASAP7_75t_L g461 ( .A(n_342), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g478 ( .A(n_342), .B(n_428), .Y(n_478) );
AND2x2_ASAP7_75t_L g533 ( .A(n_342), .B(n_427), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx4_ASAP7_75t_L g400 ( .A(n_345), .Y(n_400) );
AND2x2_ASAP7_75t_L g410 ( .A(n_345), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx2_ASAP7_75t_L g415 ( .A(n_348), .Y(n_415) );
AND2x2_ASAP7_75t_L g424 ( .A(n_348), .B(n_408), .Y(n_424) );
INVx1_ASAP7_75t_L g459 ( .A(n_350), .Y(n_459) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g380 ( .A(n_351), .Y(n_380) );
INVxp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_353), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_354), .B(n_422), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_363), .B(n_368), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_361), .B(n_400), .Y(n_509) );
INVx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
AOI21xp33_ASAP7_75t_SL g372 ( .A1(n_364), .A2(n_373), .B(n_375), .Y(n_372) );
AND2x2_ASAP7_75t_L g519 ( .A(n_364), .B(n_378), .Y(n_519) );
AND2x4_ASAP7_75t_L g382 ( .A(n_365), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_SL g416 ( .A(n_365), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_365), .B(n_432), .Y(n_498) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI21xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_381), .B(n_386), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_378), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_378), .B(n_383), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_379), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g441 ( .A(n_379), .Y(n_441) );
INVx1_ASAP7_75t_L g445 ( .A(n_379), .Y(n_445) );
AND2x2_ASAP7_75t_L g529 ( .A(n_379), .B(n_497), .Y(n_529) );
AND2x2_ASAP7_75t_L g532 ( .A(n_379), .B(n_449), .Y(n_532) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_SL g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_384), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVx1_ASAP7_75t_L g511 ( .A(n_388), .Y(n_511) );
AND2x2_ASAP7_75t_L g402 ( .A(n_389), .B(n_403), .Y(n_402) );
NAND4xp75_ASAP7_75t_L g392 ( .A(n_393), .B(n_412), .C(n_433), .D(n_451), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_404), .Y(n_393) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g482 ( .A(n_396), .B(n_483), .Y(n_482) );
NAND2x1p5_ASAP7_75t_L g468 ( .A(n_397), .B(n_462), .Y(n_468) );
NAND2xp5_ASAP7_75t_R g484 ( .A(n_400), .B(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g534 ( .A(n_400), .Y(n_534) );
INVx2_ASAP7_75t_L g447 ( .A(n_402), .Y(n_447) );
BUFx3_ASAP7_75t_L g439 ( .A(n_403), .Y(n_439) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g490 ( .A(n_408), .Y(n_490) );
AND2x2_ASAP7_75t_L g444 ( .A(n_410), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g466 ( .A(n_411), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_417), .B(n_419), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_415), .B(n_449), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_416), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_418), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_423), .B1(n_425), .B2(n_429), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
OA21x2_ASAP7_75t_L g434 ( .A1(n_427), .A2(n_435), .B(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g455 ( .A(n_427), .Y(n_455) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g486 ( .A(n_428), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g494 ( .A(n_428), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_429), .B(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g464 ( .A(n_432), .B(n_465), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_440), .B(n_442), .Y(n_433) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g481 ( .A(n_438), .B(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_445), .Y(n_493) );
INVx2_ASAP7_75t_SL g485 ( .A(n_449), .Y(n_485) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_463), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_456), .B1(n_458), .B2(n_461), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g514 ( .A(n_458), .Y(n_514) );
NOR2x1_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_506), .Y(n_469) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_479), .C(n_491), .Y(n_470) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_472), .B(n_476), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
AOI22xp33_ASAP7_75t_SL g479 ( .A1(n_480), .A2(n_484), .B1(n_486), .B2(n_488), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NOR3xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_495), .C(n_502), .Y(n_491) );
AOI21xp33_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_499), .B(n_500), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_525), .Y(n_506) );
NOR3xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_515), .C(n_522), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B1(n_513), .B2(n_514), .Y(n_508) );
OR2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
NOR3xp33_ASAP7_75t_L g522 ( .A(n_516), .B(n_521), .C(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVxp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AOI222xp33_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_529), .B1(n_530), .B2(n_532), .C1(n_533), .C2(n_534), .Y(n_525) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OAI222xp33_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B1(n_546), .B2(n_549), .C1(n_552), .C2(n_555), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_547), .Y(n_546) );
CKINVDCx16_ASAP7_75t_R g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
CKINVDCx16_ASAP7_75t_R g552 ( .A(n_553), .Y(n_552) );
endmodule