module real_jpeg_11914_n_16 (n_5, n_4, n_8, n_0, n_12, n_318, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_318;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g102 ( 
.A(n_0),
.Y(n_102)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_4),
.A2(n_39),
.B1(n_40),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_4),
.A2(n_24),
.B1(n_26),
.B2(n_62),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_62),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_4),
.A2(n_62),
.B1(n_67),
.B2(n_71),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_5),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_163),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_5),
.A2(n_24),
.B1(n_26),
.B2(n_163),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_5),
.A2(n_67),
.B1(n_71),
.B2(n_163),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_6),
.A2(n_24),
.B1(n_26),
.B2(n_47),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_6),
.A2(n_47),
.B1(n_67),
.B2(n_71),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_7),
.A2(n_24),
.B1(n_26),
.B2(n_33),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_7),
.A2(n_33),
.B1(n_67),
.B2(n_71),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_7),
.A2(n_33),
.B1(n_39),
.B2(n_40),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_10),
.A2(n_38),
.B(n_39),
.C(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_10),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_177),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_10),
.B(n_49),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_10),
.A2(n_24),
.B1(n_26),
.B2(n_177),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_10),
.A2(n_134),
.B1(n_135),
.B2(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_10),
.B(n_31),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_11),
.A2(n_39),
.B1(n_40),
.B2(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_11),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_184),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_11),
.A2(n_24),
.B1(n_26),
.B2(n_184),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_11),
.A2(n_67),
.B1(n_71),
.B2(n_184),
.Y(n_263)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_13),
.A2(n_39),
.B1(n_40),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_13),
.A2(n_51),
.B1(n_67),
.B2(n_71),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_13),
.A2(n_24),
.B1(n_26),
.B2(n_51),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_14),
.A2(n_39),
.B1(n_40),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_14),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_118),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_14),
.A2(n_24),
.B1(n_26),
.B2(n_118),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_14),
.A2(n_67),
.B1(n_71),
.B2(n_118),
.Y(n_257)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_91),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_89),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_75),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_19),
.B(n_75),
.Y(n_90)
);

BUFx24_ASAP7_75t_SL g315 ( 
.A(n_19),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_34),
.CI(n_52),
.CON(n_19),
.SN(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_31),
.B(n_32),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_21),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_21),
.A2(n_31),
.B1(n_85),
.B2(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_21),
.A2(n_32),
.B(n_88),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_21),
.A2(n_31),
.B1(n_180),
.B2(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_21),
.A2(n_31),
.B1(n_213),
.B2(n_226),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_22),
.B(n_58),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_22),
.A2(n_56),
.B(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_22),
.A2(n_86),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

OA22x2_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_22)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_23),
.A2(n_26),
.B(n_225),
.C(n_227),
.Y(n_224)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_24),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_24),
.A2(n_26),
.B1(n_69),
.B2(n_70),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g227 ( 
.A(n_24),
.B(n_27),
.C(n_29),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_26),
.B(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_30),
.B1(n_38),
.B2(n_43),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g176 ( 
.A1(n_29),
.A2(n_43),
.B(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g226 ( 
.A(n_30),
.B(n_177),
.CON(n_226),
.SN(n_226)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_32),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_45),
.B(n_48),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_35),
.A2(n_116),
.B(n_119),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_35),
.A2(n_48),
.B(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_35),
.A2(n_44),
.B1(n_182),
.B2(n_185),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_46),
.B1(n_49),
.B2(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_36),
.B(n_50),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_36),
.A2(n_49),
.B1(n_117),
.B2(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_36),
.A2(n_49),
.B1(n_183),
.B2(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_44),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_37)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_61),
.B(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_49),
.B(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.C(n_63),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_64),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_55),
.A2(n_86),
.B(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_63),
.A2(n_64),
.B1(n_82),
.B2(n_83),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_79),
.C(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_72),
.B(n_74),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_65),
.A2(n_72),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_65),
.B(n_74),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_65),
.A2(n_72),
.B1(n_232),
.B2(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_65),
.A2(n_72),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_65),
.A2(n_72),
.B1(n_240),
.B2(n_250),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_66),
.B(n_129),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_66),
.A2(n_111),
.B(n_127),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_66),
.B(n_177),
.Y(n_266)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_66)
);

CKINVDCx6p67_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_69),
.B(n_71),
.C(n_177),
.Y(n_247)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_102),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_71),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_72),
.B(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_72),
.A2(n_112),
.B(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_72),
.A2(n_74),
.B(n_139),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_72),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.C(n_81),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_76),
.A2(n_77),
.B1(n_79),
.B2(n_305),
.Y(n_308)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_79),
.A2(n_303),
.B1(n_304),
.B2(n_305),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_79),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_81),
.B(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B(n_87),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_299),
.B(n_312),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_164),
.B(n_298),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_146),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_94),
.B(n_146),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_121),
.B2(n_145),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_95),
.B(n_122),
.C(n_131),
.Y(n_310)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_113),
.C(n_115),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_97),
.A2(n_98),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_108),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_99),
.A2(n_100),
.B1(n_108),
.B2(n_109),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_101),
.A2(n_134),
.B(n_257),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_102),
.A2(n_107),
.B1(n_156),
.B2(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_102),
.A2(n_107),
.B1(n_254),
.B2(n_256),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_103),
.A2(n_107),
.B(n_158),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_104),
.A2(n_135),
.B(n_174),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_106),
.B(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_115),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_114),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_131),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_125),
.B(n_130),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_123),
.B(n_125),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_126),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_130),
.B(n_302),
.C(n_306),
.Y(n_301)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_130),
.B(n_302),
.CI(n_306),
.CON(n_311),
.SN(n_311)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_140),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g306 ( 
.A1(n_132),
.A2(n_133),
.B(n_142),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_133),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_137),
.B1(n_138),
.B2(n_141),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B(n_136),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_155),
.B(n_157),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_134),
.A2(n_135),
.B1(n_255),
.B2(n_263),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_135),
.B(n_177),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.C(n_152),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_151),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_152),
.B(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_160),
.C(n_161),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_159),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_159),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_161),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_162),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_292),
.B(n_297),
.Y(n_164)
);

AOI221xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_201),
.B1(n_217),
.B2(n_291),
.C(n_318),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_190),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_167),
.B(n_190),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_186),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_168),
.B(n_187),
.C(n_188),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_178),
.C(n_181),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_170),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_178),
.B(n_181),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.C(n_200),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_200),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.C(n_198),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_196),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_197),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_215),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_202),
.B(n_215),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.C(n_207),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_203),
.B(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_205),
.B(n_207),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.C(n_211),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_211),
.B(n_234),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_290),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_285),
.B(n_289),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_241),
.B(n_284),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_236),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_221),
.B(n_236),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_233),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_229),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_223),
.B(n_229),
.C(n_233),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_224),
.B(n_228),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.C(n_239),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_237),
.B(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_238),
.B(n_239),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_279),
.B(n_283),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_269),
.B(n_278),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_258),
.B(n_268),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_253),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_253),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_248),
.B1(n_251),
.B2(n_252),
.Y(n_245)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_246),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_251),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_264),
.B(n_267),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_266),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_271),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_274),
.C(n_277),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_276),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_282),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_288),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_294),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_309),
.Y(n_299)
);

AOI21xp33_ASAP7_75t_L g312 ( 
.A1(n_300),
.A2(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_307),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_307),
.Y(n_314)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_311),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_311),
.Y(n_316)
);


endmodule