module fake_aes_632_n_712 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_712);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_712;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_415;
wire n_235;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g80 ( .A(n_46), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_9), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_9), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_26), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_71), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_11), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_2), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_36), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_76), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_15), .Y(n_89) );
INVxp33_ASAP7_75t_L g90 ( .A(n_14), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_49), .Y(n_91) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_25), .Y(n_92) );
CKINVDCx14_ASAP7_75t_R g93 ( .A(n_17), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_30), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_40), .Y(n_95) );
INVx2_ASAP7_75t_SL g96 ( .A(n_45), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_18), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_13), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_21), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_55), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_75), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_65), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_34), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_78), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_35), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_50), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_3), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_38), .Y(n_108) );
OR2x2_ASAP7_75t_L g109 ( .A(n_43), .B(n_47), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_44), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_11), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_23), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_12), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_79), .Y(n_114) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_56), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_1), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_62), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_42), .Y(n_118) );
INVxp33_ASAP7_75t_L g119 ( .A(n_63), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_10), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_77), .Y(n_121) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_52), .Y(n_122) );
INVxp33_ASAP7_75t_L g123 ( .A(n_13), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_53), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_27), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_33), .Y(n_126) );
INVxp33_ASAP7_75t_SL g127 ( .A(n_58), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_114), .B(n_0), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_101), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_99), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_111), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_114), .B(n_0), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_113), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_111), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_101), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_111), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_88), .Y(n_137) );
AND2x2_ASAP7_75t_SL g138 ( .A(n_109), .B(n_31), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_88), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_91), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_101), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_113), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g143 ( .A(n_93), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_91), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_99), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_84), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_94), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_87), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_94), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_95), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_95), .Y(n_151) );
BUFx8_ASAP7_75t_L g152 ( .A(n_109), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_90), .B(n_1), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_102), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_102), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_92), .B(n_2), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_81), .Y(n_157) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_82), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_105), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_86), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_105), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_122), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_103), .B(n_3), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_85), .B(n_4), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_96), .Y(n_165) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_85), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_123), .B(n_4), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_106), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_106), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_108), .Y(n_170) );
INVxp33_ASAP7_75t_L g171 ( .A(n_89), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_127), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_130), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_164), .Y(n_174) );
INVxp67_ASAP7_75t_L g175 ( .A(n_158), .Y(n_175) );
NOR2xp33_ASAP7_75t_R g176 ( .A(n_143), .B(n_83), .Y(n_176) );
OA22x2_ASAP7_75t_L g177 ( .A1(n_158), .A2(n_120), .B1(n_89), .B2(n_97), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_129), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_145), .Y(n_179) );
NAND2x1p5_ASAP7_75t_L g180 ( .A(n_132), .B(n_97), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_132), .B(n_98), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_132), .B(n_98), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_171), .B(n_119), .Y(n_183) );
AO22x1_ASAP7_75t_L g184 ( .A1(n_152), .A2(n_80), .B1(n_100), .B2(n_115), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_164), .A2(n_116), .B1(n_107), .B2(n_120), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_137), .B(n_96), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_164), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_129), .Y(n_188) );
OR2x2_ASAP7_75t_L g189 ( .A(n_166), .B(n_107), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_129), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_129), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_137), .B(n_104), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_166), .B(n_116), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_138), .A2(n_153), .B1(n_167), .B2(n_152), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_139), .B(n_104), .Y(n_195) );
INVx5_ASAP7_75t_L g196 ( .A(n_165), .Y(n_196) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_157), .Y(n_197) );
NOR2xp33_ASAP7_75t_SL g198 ( .A(n_152), .B(n_80), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_139), .B(n_110), .Y(n_199) );
INVx3_ASAP7_75t_L g200 ( .A(n_164), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_147), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_140), .B(n_117), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_147), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_153), .B(n_124), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_147), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_129), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_140), .B(n_126), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_129), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_147), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_154), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_144), .B(n_149), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_154), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_153), .B(n_126), .Y(n_214) );
INVx1_ASAP7_75t_SL g215 ( .A(n_160), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_144), .B(n_125), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_129), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_165), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_148), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_149), .B(n_125), .Y(n_220) );
OR2x6_ASAP7_75t_L g221 ( .A(n_128), .B(n_121), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_165), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_150), .B(n_121), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_165), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_167), .B(n_118), .Y(n_225) );
INVx4_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
NAND2x1p5_ASAP7_75t_L g227 ( .A(n_167), .B(n_118), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_154), .Y(n_228) );
OR2x2_ASAP7_75t_L g229 ( .A(n_128), .B(n_112), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_154), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_161), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_176), .Y(n_232) );
BUFx3_ASAP7_75t_L g233 ( .A(n_211), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_211), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_209), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_219), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_209), .Y(n_237) );
BUFx4f_ASAP7_75t_L g238 ( .A(n_221), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_209), .Y(n_239) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_175), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_228), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_183), .B(n_152), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_228), .Y(n_243) );
BUFx2_ASAP7_75t_L g244 ( .A(n_221), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_183), .B(n_150), .Y(n_245) );
BUFx2_ASAP7_75t_L g246 ( .A(n_221), .Y(n_246) );
BUFx3_ASAP7_75t_L g247 ( .A(n_211), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_228), .Y(n_248) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_215), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_201), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_229), .B(n_151), .Y(n_251) );
NOR2x1_ASAP7_75t_L g252 ( .A(n_221), .B(n_156), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_193), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_203), .Y(n_254) );
OR2x6_ASAP7_75t_L g255 ( .A(n_180), .B(n_156), .Y(n_255) );
NOR2xp33_ASAP7_75t_R g256 ( .A(n_173), .B(n_179), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_214), .B(n_151), .Y(n_257) );
BUFx12f_ASAP7_75t_L g258 ( .A(n_173), .Y(n_258) );
INVxp33_ASAP7_75t_SL g259 ( .A(n_198), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_219), .Y(n_260) );
NOR3xp33_ASAP7_75t_L g261 ( .A(n_184), .B(n_146), .C(n_163), .Y(n_261) );
INVx4_ASAP7_75t_L g262 ( .A(n_200), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_176), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_193), .B(n_138), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_205), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_204), .B(n_172), .Y(n_266) );
INVx5_ASAP7_75t_L g267 ( .A(n_212), .Y(n_267) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_222), .Y(n_268) );
AND2x6_ASAP7_75t_SL g269 ( .A(n_193), .B(n_163), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_212), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_180), .B(n_181), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_225), .B(n_162), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_212), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_210), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_181), .B(n_169), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_181), .B(n_169), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_226), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_213), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_227), .Y(n_279) );
BUFx4f_ASAP7_75t_L g280 ( .A(n_227), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_226), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_230), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_200), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_182), .B(n_168), .Y(n_284) );
NOR3xp33_ASAP7_75t_SL g285 ( .A(n_179), .B(n_168), .C(n_112), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_226), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_177), .A2(n_138), .B1(n_161), .B2(n_165), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_231), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_222), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_182), .B(n_161), .Y(n_290) );
INVx3_ASAP7_75t_L g291 ( .A(n_200), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_174), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_187), .Y(n_293) );
NAND2xp33_ASAP7_75t_SL g294 ( .A(n_185), .B(n_142), .Y(n_294) );
NOR2xp67_ASAP7_75t_L g295 ( .A(n_194), .B(n_161), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_182), .B(n_133), .Y(n_296) );
NOR2xp33_ASAP7_75t_SL g297 ( .A(n_197), .B(n_170), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_267), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_276), .B(n_195), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_264), .A2(n_177), .B1(n_216), .B2(n_195), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_283), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_276), .B(n_251), .Y(n_302) );
AO32x2_ASAP7_75t_L g303 ( .A1(n_262), .A2(n_223), .A3(n_220), .B1(n_141), .B2(n_135), .Y(n_303) );
BUFx12f_ASAP7_75t_L g304 ( .A(n_258), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_253), .Y(n_305) );
OAI22xp33_ASAP7_75t_L g306 ( .A1(n_238), .A2(n_189), .B1(n_192), .B2(n_207), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_249), .B(n_216), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_240), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_283), .Y(n_309) );
NOR3xp33_ASAP7_75t_L g310 ( .A(n_294), .B(n_199), .C(n_202), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_267), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_247), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_280), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_276), .B(n_216), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_247), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_256), .Y(n_316) );
OR2x6_ASAP7_75t_L g317 ( .A(n_255), .B(n_170), .Y(n_317) );
AND2x2_ASAP7_75t_SL g318 ( .A(n_238), .B(n_223), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_271), .Y(n_319) );
INVx4_ASAP7_75t_L g320 ( .A(n_238), .Y(n_320) );
OR2x6_ASAP7_75t_L g321 ( .A(n_255), .B(n_170), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_279), .B(n_186), .Y(n_322) );
A2O1A1Ixp33_ASAP7_75t_L g323 ( .A1(n_295), .A2(n_220), .B(n_186), .C(n_159), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_247), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_242), .B(n_159), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_271), .B(n_159), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_233), .Y(n_327) );
AOI22xp33_ASAP7_75t_SL g328 ( .A1(n_297), .A2(n_155), .B1(n_108), .B2(n_136), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_255), .B(n_155), .Y(n_329) );
CKINVDCx11_ASAP7_75t_R g330 ( .A(n_258), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_233), .Y(n_331) );
BUFx4_ASAP7_75t_SL g332 ( .A(n_236), .Y(n_332) );
BUFx2_ASAP7_75t_L g333 ( .A(n_255), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_234), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_234), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_244), .A2(n_155), .B1(n_141), .B2(n_135), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_276), .B(n_131), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_262), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_283), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_279), .B(n_131), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_291), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_255), .B(n_134), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_245), .A2(n_218), .B(n_224), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_296), .B(n_134), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_244), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_246), .Y(n_346) );
NOR2xp33_ASAP7_75t_SL g347 ( .A(n_280), .B(n_135), .Y(n_347) );
INVx2_ASAP7_75t_SL g348 ( .A(n_280), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_272), .B(n_246), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_275), .B(n_136), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_287), .A2(n_141), .B1(n_196), .B2(n_218), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_267), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_252), .B(n_196), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_301), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_302), .B(n_279), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_308), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_317), .A2(n_295), .B1(n_252), .B2(n_292), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_301), .Y(n_358) );
OAI211xp5_ASAP7_75t_SL g359 ( .A1(n_300), .A2(n_285), .B(n_266), .C(n_261), .Y(n_359) );
CKINVDCx8_ASAP7_75t_R g360 ( .A(n_317), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_309), .Y(n_361) );
CKINVDCx16_ASAP7_75t_R g362 ( .A(n_304), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_330), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_298), .Y(n_364) );
OAI211xp5_ASAP7_75t_L g365 ( .A1(n_300), .A2(n_263), .B(n_232), .C(n_260), .Y(n_365) );
CKINVDCx11_ASAP7_75t_R g366 ( .A(n_304), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_298), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_309), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_343), .A2(n_293), .B(n_292), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_317), .A2(n_293), .B1(n_259), .B2(n_284), .Y(n_370) );
INVx3_ASAP7_75t_L g371 ( .A(n_311), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_326), .B(n_257), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_306), .A2(n_290), .B1(n_265), .B2(n_250), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_349), .A2(n_262), .B1(n_291), .B2(n_232), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_306), .B(n_269), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_311), .Y(n_376) );
AOI21xp33_ASAP7_75t_L g377 ( .A1(n_349), .A2(n_263), .B(n_262), .Y(n_377) );
NOR2xp67_ASAP7_75t_L g378 ( .A(n_320), .B(n_267), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_338), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_307), .B(n_248), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_345), .A2(n_291), .B1(n_248), .B2(n_250), .Y(n_381) );
BUFx2_ASAP7_75t_SL g382 ( .A(n_320), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_321), .A2(n_278), .B1(n_265), .B2(n_282), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_319), .B(n_269), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_346), .A2(n_248), .B1(n_274), .B2(n_254), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_299), .B(n_254), .Y(n_386) );
OA21x2_ASAP7_75t_L g387 ( .A1(n_323), .A2(n_325), .B(n_191), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_352), .Y(n_388) );
AOI22xp33_ASAP7_75t_SL g389 ( .A1(n_375), .A2(n_333), .B1(n_318), .B2(n_321), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_359), .A2(n_310), .B1(n_318), .B2(n_321), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_370), .A2(n_329), .B1(n_322), .B2(n_346), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_372), .B(n_323), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_368), .Y(n_393) );
INVx2_ASAP7_75t_SL g394 ( .A(n_364), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_356), .B(n_342), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_372), .B(n_325), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_354), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g398 ( .A1(n_370), .A2(n_316), .B1(n_347), .B2(n_322), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_386), .B(n_314), .Y(n_399) );
INVx4_ASAP7_75t_L g400 ( .A(n_364), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_384), .A2(n_322), .B1(n_344), .B2(n_340), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_357), .A2(n_340), .B1(n_331), .B2(n_305), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_356), .B(n_337), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_355), .B(n_303), .Y(n_404) );
OAI21x1_ASAP7_75t_L g405 ( .A1(n_369), .A2(n_351), .B(n_336), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_382), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_357), .A2(n_331), .B1(n_315), .B2(n_328), .Y(n_407) );
AO21x2_ASAP7_75t_L g408 ( .A1(n_373), .A2(n_350), .B(n_303), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_373), .B(n_274), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_365), .A2(n_334), .B1(n_335), .B2(n_348), .C(n_313), .Y(n_410) );
OA21x2_ASAP7_75t_L g411 ( .A1(n_383), .A2(n_178), .B(n_206), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_383), .A2(n_353), .B1(n_278), .B2(n_282), .C(n_315), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_362), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_362), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_380), .B(n_312), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_377), .A2(n_353), .B1(n_341), .B2(n_339), .C(n_239), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_360), .A2(n_324), .B1(n_312), .B2(n_327), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_392), .B(n_387), .Y(n_418) );
NAND2x1_ASAP7_75t_L g419 ( .A(n_393), .B(n_387), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_395), .B(n_387), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_397), .B(n_354), .Y(n_421) );
NAND3xp33_ASAP7_75t_L g422 ( .A(n_390), .B(n_387), .C(n_385), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_393), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_392), .B(n_358), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_389), .A2(n_382), .B1(n_374), .B2(n_312), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_393), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_400), .Y(n_427) );
INVx4_ASAP7_75t_L g428 ( .A(n_400), .Y(n_428) );
INVx5_ASAP7_75t_L g429 ( .A(n_400), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_391), .A2(n_312), .B1(n_324), .B2(n_381), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_397), .B(n_368), .Y(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_400), .B(n_367), .Y(n_432) );
OAI211xp5_ASAP7_75t_SL g433 ( .A1(n_401), .A2(n_330), .B(n_366), .C(n_360), .Y(n_433) );
OAI22xp33_ASAP7_75t_L g434 ( .A1(n_396), .A2(n_380), .B1(n_358), .B2(n_361), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_398), .A2(n_324), .B1(n_327), .B2(n_388), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_406), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_411), .Y(n_437) );
AO21x2_ASAP7_75t_L g438 ( .A1(n_409), .A2(n_361), .B(n_379), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_394), .B(n_367), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_395), .B(n_368), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_411), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_409), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_406), .Y(n_443) );
NOR4xp25_ASAP7_75t_SL g444 ( .A(n_410), .B(n_363), .C(n_332), .D(n_303), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_394), .Y(n_445) );
OR2x6_ASAP7_75t_L g446 ( .A(n_417), .B(n_364), .Y(n_446) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_396), .A2(n_378), .B1(n_388), .B2(n_379), .C(n_338), .Y(n_447) );
NOR2x1_ASAP7_75t_L g448 ( .A(n_417), .B(n_388), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_411), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_415), .B(n_367), .Y(n_450) );
NAND4xp25_ASAP7_75t_SL g451 ( .A(n_410), .B(n_332), .C(n_379), .D(n_7), .Y(n_451) );
BUFx2_ASAP7_75t_L g452 ( .A(n_427), .Y(n_452) );
NAND4xp25_ASAP7_75t_SL g453 ( .A(n_425), .B(n_412), .C(n_402), .D(n_407), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_431), .B(n_404), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_431), .B(n_404), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_433), .B(n_413), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_420), .B(n_403), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_429), .B(n_412), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_420), .B(n_403), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_428), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_431), .B(n_408), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_442), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_423), .B(n_426), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_442), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_440), .Y(n_465) );
AO31x2_ASAP7_75t_L g466 ( .A1(n_437), .A2(n_399), .A3(n_408), .B(n_411), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_438), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_427), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_438), .Y(n_469) );
AOI211xp5_ASAP7_75t_L g470 ( .A1(n_451), .A2(n_414), .B(n_378), .C(n_399), .Y(n_470) );
OAI31xp33_ASAP7_75t_L g471 ( .A1(n_451), .A2(n_415), .A3(n_352), .B(n_367), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_440), .B(n_408), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_421), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_438), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_418), .B(n_408), .Y(n_475) );
INVx1_ASAP7_75t_SL g476 ( .A(n_427), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_418), .B(n_371), .Y(n_477) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_428), .A2(n_376), .B1(n_371), .B2(n_405), .Y(n_478) );
OAI221xp5_ASAP7_75t_L g479 ( .A1(n_433), .A2(n_416), .B1(n_376), .B2(n_371), .C(n_327), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_423), .B(n_371), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_421), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_434), .A2(n_416), .B1(n_376), .B2(n_324), .Y(n_482) );
NAND4xp25_ASAP7_75t_L g483 ( .A(n_422), .B(n_178), .C(n_191), .D(n_206), .Y(n_483) );
OAI221xp5_ASAP7_75t_L g484 ( .A1(n_435), .A2(n_376), .B1(n_327), .B2(n_235), .C(n_239), .Y(n_484) );
OAI31xp33_ASAP7_75t_L g485 ( .A1(n_434), .A2(n_235), .A3(n_237), .B(n_241), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_436), .Y(n_486) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_447), .A2(n_237), .B1(n_303), .B2(n_243), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_423), .Y(n_488) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_426), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_426), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_438), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_424), .B(n_5), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_450), .B(n_405), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_437), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_429), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_437), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_441), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_450), .B(n_5), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_447), .A2(n_241), .B1(n_243), .B2(n_288), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_481), .B(n_424), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_461), .B(n_441), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_461), .B(n_441), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_473), .B(n_450), .Y(n_503) );
NOR2xp67_ASAP7_75t_L g504 ( .A(n_460), .B(n_429), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_454), .B(n_449), .Y(n_505) );
NOR2xp33_ASAP7_75t_R g506 ( .A(n_460), .B(n_429), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_494), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_457), .B(n_419), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_462), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_454), .B(n_449), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_455), .B(n_449), .Y(n_511) );
NOR2xp33_ASAP7_75t_R g512 ( .A(n_460), .B(n_429), .Y(n_512) );
NAND2xp33_ASAP7_75t_R g513 ( .A(n_452), .B(n_444), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_462), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_453), .A2(n_422), .B1(n_446), .B2(n_450), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_465), .B(n_436), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_457), .B(n_436), .Y(n_517) );
INVxp67_ASAP7_75t_L g518 ( .A(n_452), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_464), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_455), .B(n_419), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_494), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_496), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_493), .B(n_464), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_497), .Y(n_524) );
NOR4xp25_ASAP7_75t_SL g525 ( .A(n_458), .B(n_444), .C(n_429), .D(n_428), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_493), .B(n_446), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_459), .B(n_443), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_496), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_497), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_463), .B(n_446), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_463), .B(n_446), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_456), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_459), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_475), .B(n_446), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_488), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_475), .B(n_446), .Y(n_536) );
NAND2xp33_ASAP7_75t_SL g537 ( .A(n_498), .B(n_428), .Y(n_537) );
INVx3_ASAP7_75t_SL g538 ( .A(n_468), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_476), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_488), .Y(n_540) );
AND2x4_ASAP7_75t_L g541 ( .A(n_477), .B(n_429), .Y(n_541) );
NAND2xp33_ASAP7_75t_L g542 ( .A(n_495), .B(n_448), .Y(n_542) );
OAI322xp33_ASAP7_75t_L g543 ( .A1(n_492), .A2(n_436), .A3(n_443), .B1(n_8), .B2(n_10), .C1(n_12), .C2(n_14), .Y(n_543) );
AND2x2_ASAP7_75t_SL g544 ( .A(n_498), .B(n_432), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_490), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_472), .B(n_477), .Y(n_546) );
NOR2x1_ASAP7_75t_L g547 ( .A(n_483), .B(n_443), .Y(n_547) );
NAND2x1p5_ASAP7_75t_L g548 ( .A(n_480), .B(n_448), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_489), .B(n_443), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_472), .B(n_432), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_490), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_480), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_466), .B(n_445), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_470), .B(n_445), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_466), .B(n_445), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_467), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_467), .Y(n_557) );
INVxp33_ASAP7_75t_L g558 ( .A(n_506), .Y(n_558) );
INVx2_ASAP7_75t_SL g559 ( .A(n_538), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_532), .B(n_479), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_533), .B(n_469), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_500), .B(n_469), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_532), .A2(n_482), .B1(n_471), .B2(n_485), .Y(n_563) );
INVxp67_ASAP7_75t_SL g564 ( .A(n_504), .Y(n_564) );
AND2x4_ASAP7_75t_SL g565 ( .A(n_541), .B(n_432), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_507), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_514), .Y(n_567) );
OAI21xp33_ASAP7_75t_L g568 ( .A1(n_515), .A2(n_478), .B(n_491), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_505), .B(n_474), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_514), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_537), .A2(n_487), .B1(n_430), .B2(n_499), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_505), .B(n_491), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_510), .B(n_474), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_544), .A2(n_439), .B1(n_486), .B2(n_432), .Y(n_574) );
OAI31xp33_ASAP7_75t_L g575 ( .A1(n_554), .A2(n_484), .A3(n_439), .B(n_8), .Y(n_575) );
OAI32xp33_ASAP7_75t_L g576 ( .A1(n_539), .A2(n_6), .A3(n_7), .B1(n_15), .B2(n_16), .Y(n_576) );
INVxp67_ASAP7_75t_SL g577 ( .A(n_553), .Y(n_577) );
AOI21xp33_ASAP7_75t_SL g578 ( .A1(n_538), .A2(n_6), .B(n_16), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_519), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_510), .B(n_466), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_543), .B(n_17), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_507), .Y(n_582) );
OAI21xp5_ASAP7_75t_SL g583 ( .A1(n_547), .A2(n_439), .B(n_19), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_519), .Y(n_584) );
AOI322xp5_ASAP7_75t_L g585 ( .A1(n_544), .A2(n_439), .A3(n_18), .B1(n_19), .B2(n_20), .C1(n_466), .C2(n_208), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_525), .A2(n_466), .B(n_288), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g587 ( .A1(n_518), .A2(n_208), .B(n_217), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_513), .A2(n_224), .B1(n_222), .B2(n_190), .Y(n_588) );
NAND3x1_ASAP7_75t_L g589 ( .A(n_512), .B(n_20), .C(n_22), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_511), .B(n_217), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_509), .Y(n_591) );
OAI221xp5_ASAP7_75t_SL g592 ( .A1(n_553), .A2(n_555), .B1(n_508), .B2(n_546), .C(n_534), .Y(n_592) );
NOR4xp25_ASAP7_75t_L g593 ( .A(n_542), .B(n_24), .C(n_28), .D(n_29), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_511), .B(n_190), .Y(n_594) );
OAI21xp5_ASAP7_75t_SL g595 ( .A1(n_541), .A2(n_190), .B(n_188), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_503), .B(n_32), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_524), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_552), .B(n_190), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_523), .B(n_517), .Y(n_599) );
NAND2xp33_ASAP7_75t_SL g600 ( .A(n_555), .B(n_188), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_541), .A2(n_196), .B1(n_222), .B2(n_224), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_521), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_508), .B(n_188), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_501), .B(n_502), .Y(n_604) );
AOI22xp5_ASAP7_75t_SL g605 ( .A1(n_520), .A2(n_37), .B1(n_39), .B2(n_41), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_534), .A2(n_224), .B1(n_188), .B2(n_196), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_523), .A2(n_289), .B1(n_268), .B2(n_281), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_521), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_524), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_529), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_529), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_600), .B(n_528), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_591), .Y(n_613) );
NOR2x1_ASAP7_75t_L g614 ( .A(n_583), .B(n_542), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_604), .B(n_546), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_566), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_559), .Y(n_617) );
INVx1_ASAP7_75t_SL g618 ( .A(n_565), .Y(n_618) );
XOR2x2_ASAP7_75t_L g619 ( .A(n_589), .B(n_550), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_580), .B(n_520), .Y(n_620) );
OAI221xp5_ASAP7_75t_SL g621 ( .A1(n_575), .A2(n_526), .B1(n_536), .B2(n_527), .C(n_531), .Y(n_621) );
AO21x1_ASAP7_75t_L g622 ( .A1(n_564), .A2(n_557), .B(n_548), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_569), .B(n_501), .Y(n_623) );
NOR4xp25_ASAP7_75t_SL g624 ( .A(n_595), .B(n_557), .C(n_535), .D(n_551), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_582), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_560), .B(n_523), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_562), .B(n_502), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_572), .B(n_527), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_560), .B(n_556), .C(n_516), .Y(n_629) );
BUFx3_ASAP7_75t_L g630 ( .A(n_602), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_567), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_561), .B(n_536), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_608), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_573), .B(n_550), .Y(n_634) );
INVx1_ASAP7_75t_SL g635 ( .A(n_558), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_570), .Y(n_636) );
OAI221xp5_ASAP7_75t_L g637 ( .A1(n_581), .A2(n_548), .B1(n_556), .B2(n_526), .C(n_535), .Y(n_637) );
NOR3x1_ASAP7_75t_L g638 ( .A(n_564), .B(n_540), .C(n_551), .Y(n_638) );
CKINVDCx16_ASAP7_75t_R g639 ( .A(n_605), .Y(n_639) );
INVxp67_ASAP7_75t_SL g640 ( .A(n_577), .Y(n_640) );
OAI21xp5_ASAP7_75t_L g641 ( .A1(n_578), .A2(n_548), .B(n_540), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_599), .B(n_531), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_579), .Y(n_643) );
NOR4xp25_ASAP7_75t_SL g644 ( .A(n_592), .B(n_530), .C(n_549), .D(n_528), .Y(n_644) );
AOI211x1_ASAP7_75t_L g645 ( .A1(n_568), .A2(n_530), .B(n_549), .C(n_522), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_584), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_577), .B(n_522), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_597), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_592), .B(n_545), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_611), .B(n_545), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_613), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_643), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_643), .Y(n_653) );
AOI322xp5_ASAP7_75t_L g654 ( .A1(n_639), .A2(n_581), .A3(n_563), .B1(n_574), .B2(n_610), .C1(n_609), .C2(n_571), .Y(n_654) );
INVxp67_ASAP7_75t_L g655 ( .A(n_626), .Y(n_655) );
XNOR2xp5_ASAP7_75t_L g656 ( .A(n_619), .B(n_563), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_631), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_649), .A2(n_596), .B1(n_603), .B2(n_588), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_649), .B(n_594), .Y(n_659) );
AOI22xp5_ASAP7_75t_SL g660 ( .A1(n_617), .A2(n_586), .B1(n_585), .B2(n_593), .Y(n_660) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_614), .A2(n_576), .B(n_587), .Y(n_661) );
NAND3x1_ASAP7_75t_L g662 ( .A(n_626), .B(n_607), .C(n_598), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_612), .A2(n_601), .B(n_590), .Y(n_663) );
AOI211x1_ASAP7_75t_L g664 ( .A1(n_637), .A2(n_606), .B(n_51), .C(n_54), .Y(n_664) );
OAI22xp5_ASAP7_75t_SL g665 ( .A1(n_635), .A2(n_606), .B1(n_57), .B2(n_59), .Y(n_665) );
NAND3xp33_ASAP7_75t_L g666 ( .A(n_629), .B(n_267), .C(n_289), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_618), .Y(n_667) );
OR2x2_ASAP7_75t_L g668 ( .A(n_623), .B(n_48), .Y(n_668) );
INVx2_ASAP7_75t_SL g669 ( .A(n_630), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_636), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_620), .B(n_60), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_620), .B(n_61), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_646), .Y(n_673) );
INVx2_ASAP7_75t_SL g674 ( .A(n_630), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_667), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g676 ( .A1(n_656), .A2(n_621), .B1(n_641), .B2(n_640), .C(n_619), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_659), .A2(n_622), .B1(n_632), .B2(n_642), .Y(n_677) );
NOR2xp33_ASAP7_75t_R g678 ( .A(n_669), .B(n_615), .Y(n_678) );
NOR2x1p5_ASAP7_75t_L g679 ( .A(n_666), .B(n_654), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_655), .B(n_645), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_657), .Y(n_681) );
NOR2xp33_ASAP7_75t_R g682 ( .A(n_674), .B(n_638), .Y(n_682) );
OAI322xp33_ASAP7_75t_L g683 ( .A1(n_660), .A2(n_628), .A3(n_627), .B1(n_634), .B2(n_648), .C1(n_650), .C2(n_647), .Y(n_683) );
AOI222xp33_ASAP7_75t_L g684 ( .A1(n_661), .A2(n_647), .B1(n_625), .B2(n_616), .C1(n_633), .C2(n_612), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_652), .B(n_644), .Y(n_685) );
NOR2xp67_ASAP7_75t_L g686 ( .A(n_666), .B(n_633), .Y(n_686) );
OAI221xp5_ASAP7_75t_L g687 ( .A1(n_661), .A2(n_650), .B1(n_625), .B2(n_616), .C(n_622), .Y(n_687) );
NOR2x1_ASAP7_75t_L g688 ( .A(n_668), .B(n_624), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_670), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_L g690 ( .A1(n_671), .A2(n_64), .B(n_66), .C(n_67), .Y(n_690) );
OAI22xp33_ASAP7_75t_SL g691 ( .A1(n_651), .A2(n_68), .B1(n_69), .B2(n_70), .Y(n_691) );
INVx1_ASAP7_75t_SL g692 ( .A(n_662), .Y(n_692) );
OAI211xp5_ASAP7_75t_SL g693 ( .A1(n_658), .A2(n_270), .B(n_286), .C(n_281), .Y(n_693) );
AOI31xp33_ASAP7_75t_L g694 ( .A1(n_663), .A2(n_72), .A3(n_73), .B(n_74), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_673), .A2(n_289), .B1(n_268), .B2(n_270), .C(n_273), .Y(n_695) );
NOR4xp25_ASAP7_75t_L g696 ( .A(n_672), .B(n_273), .C(n_277), .D(n_286), .Y(n_696) );
OA22x2_ASAP7_75t_L g697 ( .A1(n_665), .A2(n_277), .B1(n_267), .B2(n_268), .Y(n_697) );
OR3x2_ASAP7_75t_L g698 ( .A(n_664), .B(n_268), .C(n_289), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_676), .A2(n_679), .B1(n_692), .B2(n_684), .Y(n_699) );
AOI22xp5_ASAP7_75t_SL g700 ( .A1(n_675), .A2(n_697), .B1(n_685), .B2(n_680), .Y(n_700) );
CKINVDCx5p33_ASAP7_75t_R g701 ( .A(n_678), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_677), .B(n_689), .Y(n_702) );
OAI221xp5_ASAP7_75t_L g703 ( .A1(n_687), .A2(n_688), .B1(n_696), .B2(n_686), .C(n_694), .Y(n_703) );
AND2x2_ASAP7_75t_SL g704 ( .A(n_699), .B(n_698), .Y(n_704) );
AO22x2_ASAP7_75t_L g705 ( .A1(n_702), .A2(n_681), .B1(n_683), .B2(n_682), .Y(n_705) );
AOI221xp5_ASAP7_75t_SL g706 ( .A1(n_703), .A2(n_691), .B1(n_690), .B2(n_682), .C(n_695), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_704), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_705), .A2(n_701), .B1(n_700), .B2(n_693), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_707), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_708), .B(n_705), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_709), .A2(n_706), .B1(n_653), .B2(n_289), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_711), .A2(n_710), .B(n_268), .Y(n_712) );
endmodule