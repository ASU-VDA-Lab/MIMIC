module fake_jpeg_869_n_65 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_65);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_65;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

BUFx12_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_18),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_22),
.Y(n_33)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_32),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_34),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_26),
.B1(n_28),
.B2(n_23),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_37),
.B(n_38),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_26),
.B1(n_23),
.B2(n_20),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_20),
.B(n_19),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_1),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_19),
.C(n_15),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_1),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_SL g49 ( 
.A1(n_44),
.A2(n_39),
.B(n_36),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_13),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_2),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_55),
.B(n_56),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

A2O1A1O1Ixp25_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_51),
.B(n_14),
.C(n_12),
.D(n_10),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_58),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_61)
);

NOR3xp33_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_4),
.C(n_5),
.Y(n_62)
);

OAI31xp33_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_60),
.A3(n_7),
.B(n_8),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_7),
.B(n_8),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);


endmodule