module fake_jpeg_1792_n_201 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_201);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_47),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_22),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_26),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_74),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_46),
.B1(n_41),
.B2(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_0),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_37),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_76),
.Y(n_87)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_58),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_86),
.Y(n_102)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_53),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_63),
.B(n_50),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_57),
.C(n_70),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_49),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_92),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_74),
.B1(n_77),
.B2(n_71),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_97),
.B1(n_100),
.B2(n_106),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_73),
.B1(n_61),
.B2(n_51),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_101),
.C(n_65),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_74),
.B1(n_77),
.B2(n_61),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_77),
.B1(n_59),
.B2(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_69),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_104),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_66),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_63),
.B1(n_60),
.B2(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_79),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_68),
.B1(n_56),
.B2(n_75),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_1),
.B(n_3),
.Y(n_126)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_65),
.C(n_68),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_56),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_75),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_110),
.B(n_4),
.Y(n_128)
);

XNOR2x1_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_115),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_90),
.B(n_84),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_123),
.B(n_33),
.Y(n_138)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

AOI32xp33_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_56),
.A3(n_65),
.B1(n_3),
.B2(n_4),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_127),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_93),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_126),
.C(n_128),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_125),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_83),
.B(n_2),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_1),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_5),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_129),
.B(n_5),
.Y(n_136)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_118),
.A2(n_108),
.B1(n_100),
.B2(n_36),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_138),
.B(n_139),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_115),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_149),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_34),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_150),
.C(n_27),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_136),
.B(n_141),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_114),
.A2(n_6),
.B(n_7),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_13),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_10),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_142)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_11),
.B(n_12),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_143),
.A2(n_14),
.B(n_15),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_144),
.A2(n_19),
.B(n_20),
.C(n_29),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_121),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_121),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_156),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_158),
.A2(n_169),
.B1(n_140),
.B2(n_131),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_139),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_159),
.B(n_160),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_137),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_165),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_16),
.Y(n_164)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_17),
.B(n_18),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_134),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_30),
.B(n_24),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_145),
.B1(n_144),
.B2(n_143),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_25),
.C(n_28),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_135),
.C(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_177),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_170),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_161),
.C(n_157),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

OAI322xp33_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_165),
.A3(n_166),
.B1(n_168),
.B2(n_167),
.C1(n_171),
.C2(n_162),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_185),
.Y(n_193)
);

NAND2xp33_ASAP7_75t_SL g194 ( 
.A(n_186),
.B(n_184),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_SL g187 ( 
.A1(n_182),
.A2(n_158),
.B(n_161),
.C(n_169),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_187),
.A2(n_179),
.B(n_169),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_163),
.C(n_169),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_177),
.B1(n_182),
.B2(n_178),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_190),
.A2(n_191),
.B(n_194),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_189),
.A2(n_174),
.B1(n_176),
.B2(n_20),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_192),
.B(n_187),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_197),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_183),
.Y(n_197)
);

AO21x1_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_191),
.B(n_196),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_199),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_200),
.B(n_192),
.Y(n_201)
);


endmodule