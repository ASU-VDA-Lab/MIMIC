module fake_jpeg_14274_n_155 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_155);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_13),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_9),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_3),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_36),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_69),
.B(n_72),
.Y(n_86)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_1),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_73),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_76),
.B(n_77),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_26),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_78),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_80),
.B(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_83),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_53),
.B(n_65),
.C(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_50),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_65),
.B(n_62),
.C(n_61),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_2),
.B(n_4),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_56),
.B1(n_55),
.B2(n_60),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_22),
.B(n_41),
.C(n_40),
.Y(n_103)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_54),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_98),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_59),
.Y(n_98)
);

AO21x2_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_29),
.B(n_42),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_110),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_31),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_93),
.B(n_4),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_103),
.B(n_99),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_32),
.Y(n_127)
);

OAI22x1_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_111),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_30),
.C(n_39),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_129),
.C(n_45),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_112),
.B(n_108),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_117),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_17),
.C(n_38),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_118),
.B(n_130),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_108),
.B(n_7),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_123),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_8),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_128),
.Y(n_141)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_10),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_99),
.C(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_112),
.B(n_11),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_133),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

NOR2xp67_ASAP7_75t_SL g142 ( 
.A(n_135),
.B(n_138),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_139),
.C(n_116),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_129),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_122),
.C(n_119),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_146),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_140),
.C(n_136),
.Y(n_149)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_141),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_149),
.C(n_144),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_150),
.A2(n_151),
.B(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_146),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_134),
.C(n_143),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_126),
.Y(n_155)
);


endmodule