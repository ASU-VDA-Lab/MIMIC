module fake_jpeg_286_n_265 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_49),
.Y(n_68)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_56),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_18),
.B(n_14),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_55),
.Y(n_77)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_12),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_29),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_12),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_10),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_63),
.Y(n_102)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_28),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_66),
.B(n_30),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_37),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_23),
.B1(n_33),
.B2(n_38),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_91),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_66),
.A2(n_26),
.B1(n_31),
.B2(n_40),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_70),
.A2(n_89),
.B1(n_53),
.B2(n_42),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_93),
.Y(n_127)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

CKINVDCx9p33_ASAP7_75t_R g80 ( 
.A(n_48),
.Y(n_80)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_98),
.Y(n_109)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_43),
.A2(n_38),
.B1(n_33),
.B2(n_30),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_88),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_31),
.B1(n_26),
.B2(n_40),
.Y(n_89)
);

HAxp5_ASAP7_75t_SL g91 ( 
.A(n_61),
.B(n_40),
.CON(n_91),
.SN(n_91)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_56),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_62),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_41),
.B(n_23),
.Y(n_98)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_60),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_102),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_104),
.B(n_103),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_50),
.C(n_54),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_105),
.B(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_106),
.Y(n_139)
);

OA21x2_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_47),
.B(n_52),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_SL g143 ( 
.A1(n_108),
.A2(n_124),
.B(n_126),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_70),
.A2(n_65),
.B(n_57),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_119),
.B(n_122),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_114),
.Y(n_144)
);

FAx1_ASAP7_75t_SL g114 ( 
.A(n_68),
.B(n_61),
.CI(n_64),
.CON(n_114),
.SN(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_31),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_26),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_39),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_133),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_87),
.A2(n_39),
.B1(n_4),
.B2(n_5),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_83),
.B(n_2),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_6),
.Y(n_154)
);

AO22x1_ASAP7_75t_SL g137 ( 
.A1(n_129),
.A2(n_73),
.B1(n_87),
.B2(n_85),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_2),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_101),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_78),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_103),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_153),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_107),
.A2(n_73),
.B1(n_94),
.B2(n_85),
.Y(n_138)
);

AO22x1_ASAP7_75t_SL g183 ( 
.A1(n_138),
.A2(n_151),
.B1(n_133),
.B2(n_123),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_136),
.Y(n_172)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_150),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_101),
.B1(n_97),
.B2(n_86),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_77),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_155),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_97),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_154),
.B(n_156),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_6),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_109),
.B(n_7),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_117),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_161),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_105),
.B(n_7),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_8),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_8),
.Y(n_182)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_131),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_170),
.C(n_186),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_122),
.B(n_110),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_167),
.A2(n_173),
.B(n_174),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_140),
.A2(n_122),
.B1(n_114),
.B2(n_119),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_106),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_108),
.B(n_114),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_108),
.B(n_135),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_176),
.B(n_157),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_140),
.B(n_129),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_166),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_141),
.B(n_121),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_181),
.B(n_185),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_157),
.Y(n_188)
);

OA21x2_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_187),
.B(n_184),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_120),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_111),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_111),
.C(n_115),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_191),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_187),
.A2(n_167),
.B1(n_173),
.B2(n_177),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_194),
.A2(n_189),
.B1(n_197),
.B2(n_201),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_180),
.B1(n_160),
.B2(n_113),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_158),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_203),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_202),
.B(n_79),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_138),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_184),
.A2(n_168),
.B(n_171),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_204),
.A2(n_139),
.B(n_149),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_149),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_150),
.Y(n_216)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_145),
.Y(n_210)
);

FAx1_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_183),
.CI(n_143),
.CON(n_207),
.SN(n_207)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_207),
.A2(n_209),
.B(n_196),
.Y(n_228)
);

AOI321xp33_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_170),
.A3(n_178),
.B1(n_183),
.B2(n_137),
.C(n_139),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_222),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_198),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_137),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_212),
.C(n_213),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_145),
.C(n_179),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_179),
.C(n_180),
.Y(n_213)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_217),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_221),
.C(n_192),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_79),
.C(n_99),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_212),
.C(n_218),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_226),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_220),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_228),
.A2(n_215),
.B(n_207),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_210),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_233),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_232),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_201),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_227),
.A2(n_215),
.B(n_189),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_234),
.A2(n_228),
.B(n_231),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_238),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_236),
.B(n_241),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_229),
.A2(n_190),
.B1(n_219),
.B2(n_207),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_SL g239 ( 
.A(n_224),
.B(n_194),
.C(n_221),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_223),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_211),
.C(n_195),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_245),
.B(n_244),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_190),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_246),
.B(n_249),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_237),
.A2(n_229),
.B1(n_192),
.B2(n_203),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_235),
.B1(n_236),
.B2(n_240),
.Y(n_251)
);

FAx1_ASAP7_75t_SL g249 ( 
.A(n_241),
.B(n_225),
.CI(n_198),
.CON(n_249),
.SN(n_249)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_251),
.B(n_79),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_8),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_252),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_132),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_253),
.B(n_247),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_258),
.Y(n_259)
);

NOR3xp33_ASAP7_75t_SL g257 ( 
.A(n_254),
.B(n_249),
.C(n_132),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_253),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_255),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_260),
.Y(n_262)
);

NOR3xp33_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_9),
.C(n_259),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_9),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_262),
.Y(n_265)
);


endmodule