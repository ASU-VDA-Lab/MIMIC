module real_jpeg_6958_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

BUFx10_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_1),
.B(n_5),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_13),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_3),
.B(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_19),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_4),
.B(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g6 ( 
.A(n_7),
.B(n_31),
.Y(n_6)
);

OAI211xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_11),
.B(n_23),
.C(n_28),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_10),
.Y(n_8)
);

AND2x2_ASAP7_75t_SL g16 ( 
.A(n_10),
.B(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_10),
.A2(n_18),
.B1(n_22),
.B2(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_10),
.B(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_10),
.B(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_15),
.Y(n_11)
);

AND2x2_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_14),
.Y(n_12)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

OR2x4_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_16),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_21),
.B(n_22),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_27),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);


endmodule