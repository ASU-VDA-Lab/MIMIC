module fake_jpeg_30992_n_90 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_90);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_90;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx3_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_43),
.Y(n_47)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2x1_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_1),
.Y(n_50)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_0),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_29),
.B1(n_35),
.B2(n_33),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_51),
.B1(n_2),
.B2(n_4),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_37),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_6),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_31),
.B1(n_34),
.B2(n_4),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_54),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_20),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_2),
.C(n_3),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_34),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_66),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_56),
.A2(n_47),
.B1(n_53),
.B2(n_55),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_58),
.B(n_62),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_61),
.Y(n_73)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_5),
.B(n_28),
.C(n_9),
.Y(n_62)
);

FAx1_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_65),
.CI(n_25),
.CON(n_76),
.SN(n_76)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_64),
.B(n_22),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_16),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_71),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_23),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_75),
.B(n_77),
.Y(n_80)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_26),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_74),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_82),
.Y(n_83)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_80),
.Y(n_85)
);

AOI31xp33_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_70),
.A3(n_72),
.B(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_86),
.B(n_70),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_88),
.A2(n_71),
.B1(n_61),
.B2(n_68),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_73),
.Y(n_90)
);


endmodule