module fake_netlist_5_1572_n_1226 (n_137, n_294, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_204, n_250, n_260, n_298, n_286, n_122, n_282, n_10, n_24, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_9, n_195, n_42, n_227, n_45, n_271, n_94, n_123, n_167, n_234, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_95, n_183, n_185, n_243, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_72, n_104, n_41, n_56, n_141, n_15, n_145, n_48, n_50, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_149, n_309, n_30, n_14, n_84, n_130, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_207, n_37, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_175, n_262, n_238, n_99, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_199, n_187, n_32, n_103, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1226);

input n_137;
input n_294;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_204;
input n_250;
input n_260;
input n_298;
input n_286;
input n_122;
input n_282;
input n_10;
input n_24;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_9;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_123;
input n_167;
input n_234;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_95;
input n_183;
input n_185;
input n_243;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_145;
input n_48;
input n_50;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_149;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_207;
input n_37;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_175;
input n_262;
input n_238;
input n_99;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_199;
input n_187;
input n_32;
input n_103;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1226;

wire n_924;
wire n_676;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_1194;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_1166;
wire n_615;
wire n_469;
wire n_851;
wire n_1060;
wire n_1141;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_1178;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_913;
wire n_865;
wire n_1161;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_1150;
wire n_1222;
wire n_605;
wire n_776;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_525;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1085;
wire n_1066;
wire n_1191;
wire n_1198;
wire n_721;
wire n_998;
wire n_1157;
wire n_841;
wire n_1099;
wire n_1050;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_1128;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_372;
wire n_443;
wire n_677;
wire n_859;
wire n_864;
wire n_1110;
wire n_951;
wire n_1121;
wire n_1203;
wire n_821;
wire n_714;
wire n_447;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_909;
wire n_625;
wire n_949;
wire n_854;
wire n_1179;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_640;
wire n_968;
wire n_624;
wire n_825;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_1195;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_1090;
wire n_1200;
wire n_633;
wire n_1192;
wire n_530;
wire n_439;
wire n_1024;
wire n_556;
wire n_1107;
wire n_1063;
wire n_448;
wire n_758;
wire n_999;
wire n_1185;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_1032;
wire n_981;
wire n_1143;
wire n_804;
wire n_867;
wire n_1124;
wire n_537;
wire n_1158;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_1182;
wire n_756;
wire n_1145;
wire n_943;
wire n_524;
wire n_878;
wire n_399;
wire n_579;
wire n_341;
wire n_394;
wire n_1049;
wire n_992;
wire n_1153;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_812;
wire n_842;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_1154;
wire n_883;
wire n_1135;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_1163;
wire n_519;
wire n_406;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1207;
wire n_1100;
wire n_1214;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_918;
wire n_942;
wire n_381;
wire n_1147;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_592;
wire n_1169;
wire n_920;
wire n_894;
wire n_1046;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_1221;
wire n_654;
wire n_370;
wire n_1172;
wire n_976;
wire n_1095;
wire n_1096;
wire n_343;
wire n_379;
wire n_428;
wire n_833;
wire n_570;
wire n_514;
wire n_457;
wire n_1045;
wire n_1079;
wire n_1208;
wire n_853;
wire n_603;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_1168;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_1201;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_1148;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_995;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_1176;
wire n_374;
wire n_339;
wire n_1149;
wire n_882;
wire n_398;
wire n_1146;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_1225;
wire n_522;
wire n_550;
wire n_696;
wire n_1020;
wire n_798;
wire n_350;
wire n_662;
wire n_459;
wire n_897;
wire n_646;
wire n_1062;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_1219;
wire n_1204;
wire n_1215;
wire n_1216;
wire n_580;
wire n_622;
wire n_1171;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_1218;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1188;
wire n_1030;
wire n_1223;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_1165;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_673;
wire n_631;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_1177;
wire n_680;
wire n_974;
wire n_432;
wire n_553;
wire n_395;
wire n_727;
wire n_839;
wire n_901;
wire n_813;
wire n_1159;
wire n_1210;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_369;
wire n_675;
wire n_888;
wire n_613;
wire n_871;
wire n_1119;
wire n_1167;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_928;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_482;
wire n_517;
wire n_342;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_1173;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_969;
wire n_866;
wire n_1069;
wire n_1132;
wire n_1075;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_903;
wire n_1006;
wire n_740;
wire n_329;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_1061;
wire n_338;
wire n_477;
wire n_571;
wire n_333;
wire n_693;
wire n_461;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_1193;
wire n_567;
wire n_1113;
wire n_652;
wire n_778;
wire n_1122;
wire n_1111;
wire n_1197;
wire n_1211;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_770;
wire n_844;
wire n_1031;
wire n_471;
wire n_609;
wire n_852;
wire n_1041;
wire n_989;
wire n_1039;
wire n_1102;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1187;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_466;
wire n_1164;
wire n_420;
wire n_630;
wire n_1202;
wire n_489;
wire n_632;
wire n_699;
wire n_1174;
wire n_979;
wire n_1002;
wire n_617;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_585;
wire n_349;
wire n_1106;
wire n_1190;
wire n_1224;
wire n_616;
wire n_953;
wire n_601;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_1212;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1183;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_1091;
wire n_494;
wire n_1217;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_1059;
wire n_1131;
wire n_1084;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_607;
wire n_425;
wire n_513;
wire n_710;
wire n_407;
wire n_527;
wire n_707;
wire n_679;
wire n_832;
wire n_795;
wire n_695;
wire n_857;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_561;
wire n_1220;
wire n_1044;
wire n_1205;
wire n_346;
wire n_937;
wire n_1209;
wire n_393;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_1027;
wire n_490;
wire n_805;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_596;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_529;
wire n_735;
wire n_702;
wire n_822;
wire n_412;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1160;
wire n_1080;
wire n_1162;
wire n_491;
wire n_1074;
wire n_427;
wire n_1199;
wire n_791;
wire n_732;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_1181;
wire n_1196;
wire n_651;
wire n_435;
wire n_809;
wire n_952;
wire n_870;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_803;
wire n_868;
wire n_1092;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_1213;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_1186;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1175;
wire n_960;
wire n_1056;
wire n_759;
wire n_1018;
wire n_1155;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_1184;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_1189;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_1180;
wire n_1206;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_950;
wire n_533;
wire n_1170;
wire n_747;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_57),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_182),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_1),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_114),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_149),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_307),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_301),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_314),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_37),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_210),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_145),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_201),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_298),
.B(n_312),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_30),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_141),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_251),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_102),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_50),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_126),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_161),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_129),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_270),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_234),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_51),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_170),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_171),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_258),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_139),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_9),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_39),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_159),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_147),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_124),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_68),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_137),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_223),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_303),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_253),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_134),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_221),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_265),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_157),
.Y(n_358)
);

BUFx10_ASAP7_75t_L g359 ( 
.A(n_144),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_75),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_29),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_254),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_156),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_173),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_50),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_205),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_269),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_34),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_38),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_315),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_19),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_278),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_175),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_200),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_45),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_155),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_116),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_46),
.Y(n_378)
);

BUFx2_ASAP7_75t_SL g379 ( 
.A(n_154),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_272),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_216),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_158),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_115),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_34),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_L g385 ( 
.A(n_125),
.B(n_261),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_49),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_255),
.B(n_104),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_8),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_59),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_48),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_101),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_56),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_218),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_99),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_211),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_63),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_165),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_90),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_61),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_133),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_4),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_110),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_204),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_94),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_10),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_279),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_109),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_316),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_263),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_18),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_190),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_233),
.Y(n_412)
);

BUFx10_ASAP7_75t_L g413 ( 
.A(n_117),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_163),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_297),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_276),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_131),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_285),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_42),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_30),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_291),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_239),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_256),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_32),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_299),
.Y(n_425)
);

BUFx10_ASAP7_75t_L g426 ( 
.A(n_67),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_186),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_107),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_5),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_86),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_277),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_4),
.Y(n_432)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_106),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_260),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_148),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_9),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_271),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_208),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_197),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_274),
.Y(n_440)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_95),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_309),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_93),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_135),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_180),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_41),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_188),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_119),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_244),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_167),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_267),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_105),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_11),
.Y(n_453)
);

BUFx2_ASAP7_75t_SL g454 ( 
.A(n_259),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_118),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_252),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_194),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_202),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_281),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_287),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_264),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_169),
.Y(n_462)
);

BUFx5_ASAP7_75t_L g463 ( 
.A(n_168),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_24),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_203),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_191),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_113),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_41),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_112),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_122),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_31),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_66),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_178),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_275),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_330),
.Y(n_475)
);

OAI22x1_ASAP7_75t_SL g476 ( 
.A1(n_429),
.A2(n_3),
.B1(n_0),
.B2(n_2),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_368),
.Y(n_477)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_391),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_391),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_325),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_356),
.B(n_0),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_325),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_350),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_325),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_325),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_320),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_399),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_391),
.Y(n_488)
);

BUFx12f_ASAP7_75t_L g489 ( 
.A(n_350),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_432),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_420),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_417),
.B(n_2),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_391),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_356),
.B(n_5),
.Y(n_494)
);

INVx5_ASAP7_75t_L g495 ( 
.A(n_459),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_471),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_447),
.B(n_6),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_459),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_417),
.B(n_6),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_459),
.Y(n_500)
);

CKINVDCx6p67_ASAP7_75t_R g501 ( 
.A(n_426),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_459),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_447),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_331),
.A2(n_89),
.B(n_88),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_472),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_472),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_472),
.Y(n_507)
);

BUFx12f_ASAP7_75t_L g508 ( 
.A(n_426),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_422),
.B(n_7),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_333),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_345),
.Y(n_511)
);

INVx5_ASAP7_75t_L g512 ( 
.A(n_359),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_360),
.Y(n_513)
);

AOI22x1_ASAP7_75t_SL g514 ( 
.A1(n_317),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_338),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_343),
.B(n_12),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_473),
.B(n_337),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_367),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_359),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_382),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_365),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_339),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_377),
.A2(n_92),
.B(n_91),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_424),
.Y(n_524)
);

INVx5_ASAP7_75t_L g525 ( 
.A(n_413),
.Y(n_525)
);

BUFx8_ASAP7_75t_SL g526 ( 
.A(n_372),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_413),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_415),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_427),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_323),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_324),
.Y(n_531)
);

OA21x2_ASAP7_75t_L g532 ( 
.A1(n_318),
.A2(n_12),
.B(n_13),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_436),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_453),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_319),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_326),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_464),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_343),
.B(n_14),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_435),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_408),
.B(n_14),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_433),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_541)
);

BUFx12f_ASAP7_75t_L g542 ( 
.A(n_334),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_468),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_445),
.B(n_15),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_463),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_460),
.B(n_16),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_470),
.Y(n_547)
);

NOR2x1_ASAP7_75t_L g548 ( 
.A(n_385),
.B(n_96),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_371),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_526),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_480),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_482),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_486),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_536),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_484),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_485),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_515),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_530),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_505),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_531),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_542),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_507),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_506),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_R g564 ( 
.A(n_489),
.B(n_433),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_503),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_508),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_501),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_503),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_496),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_527),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_510),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_512),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_475),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_479),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_477),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_487),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_522),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_509),
.B(n_444),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_488),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_519),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_490),
.Y(n_581)
);

NAND2xp33_ASAP7_75t_SL g582 ( 
.A(n_516),
.B(n_340),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_538),
.A2(n_441),
.B1(n_397),
.B2(n_418),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_525),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_525),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_510),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_525),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_535),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_488),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_517),
.B(n_441),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_522),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_510),
.B(n_322),
.Y(n_592)
);

NOR2xp67_ASAP7_75t_L g593 ( 
.A(n_554),
.B(n_478),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_L g594 ( 
.A(n_590),
.B(n_499),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_578),
.A2(n_492),
.B1(n_439),
.B2(n_449),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_558),
.Y(n_596)
);

AO21x2_ASAP7_75t_L g597 ( 
.A1(n_583),
.A2(n_523),
.B(n_504),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_577),
.B(n_478),
.Y(n_598)
);

AND2x6_ASAP7_75t_SL g599 ( 
.A(n_573),
.B(n_481),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_575),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_564),
.B(n_570),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_576),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_591),
.B(n_495),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_560),
.B(n_549),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_R g605 ( 
.A(n_550),
.B(n_393),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_579),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_579),
.B(n_495),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_564),
.B(n_483),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_572),
.B(n_491),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_571),
.B(n_481),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_571),
.B(n_518),
.Y(n_611)
);

NAND3xp33_ASAP7_75t_L g612 ( 
.A(n_582),
.B(n_541),
.C(n_546),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_574),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_586),
.Y(n_614)
);

AO221x1_ASAP7_75t_L g615 ( 
.A1(n_565),
.A2(n_336),
.B1(n_342),
.B2(n_335),
.C(n_327),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_586),
.B(n_520),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_580),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_574),
.B(n_495),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_589),
.B(n_540),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_589),
.B(n_540),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_592),
.B(n_520),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_568),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_551),
.B(n_528),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_553),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_585),
.B(n_494),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_551),
.B(n_562),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_563),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_581),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_552),
.B(n_528),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_555),
.B(n_528),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_584),
.B(n_534),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_587),
.B(n_497),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_556),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_559),
.B(n_497),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_561),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_569),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_L g637 ( 
.A(n_567),
.B(n_548),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_566),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_557),
.B(n_529),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_590),
.B(n_539),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_588),
.Y(n_641)
);

BUFx5_ASAP7_75t_L g642 ( 
.A(n_552),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_588),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_578),
.A2(n_456),
.B1(n_370),
.B2(n_412),
.Y(n_644)
);

BUFx5_ASAP7_75t_L g645 ( 
.A(n_552),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_590),
.B(n_544),
.Y(n_646)
);

CKINVDCx14_ASAP7_75t_R g647 ( 
.A(n_564),
.Y(n_647)
);

OR2x6_ASAP7_75t_L g648 ( 
.A(n_624),
.B(n_379),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_610),
.B(n_511),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_594),
.A2(n_321),
.B1(n_332),
.B2(n_328),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_627),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_633),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_605),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_644),
.B(n_341),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_640),
.B(n_547),
.Y(n_655)
);

CKINVDCx11_ASAP7_75t_R g656 ( 
.A(n_599),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_626),
.Y(n_657)
);

INVxp33_ASAP7_75t_L g658 ( 
.A(n_628),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_635),
.B(n_454),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_614),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_634),
.B(n_544),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_639),
.B(n_346),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_610),
.B(n_513),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_606),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_635),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_612),
.A2(n_344),
.B1(n_349),
.B2(n_348),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_593),
.B(n_596),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_635),
.B(n_387),
.Y(n_668)
);

BUFx4f_ASAP7_75t_L g669 ( 
.A(n_636),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_595),
.A2(n_329),
.B1(n_351),
.B2(n_347),
.Y(n_670)
);

NOR2x1p5_ASAP7_75t_L g671 ( 
.A(n_596),
.B(n_361),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_609),
.B(n_369),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_602),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_622),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_632),
.A2(n_354),
.B1(n_355),
.B2(n_353),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_623),
.Y(n_676)
);

NOR2x2_ASAP7_75t_L g677 ( 
.A(n_631),
.B(n_476),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_647),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_631),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_611),
.B(n_521),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_619),
.B(n_620),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_641),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_613),
.B(n_352),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_597),
.A2(n_545),
.B(n_498),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_643),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_617),
.B(n_357),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_622),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_616),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_622),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_642),
.B(n_358),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_629),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_630),
.Y(n_692)
);

NAND3xp33_ASAP7_75t_SL g693 ( 
.A(n_608),
.B(n_378),
.C(n_375),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_625),
.B(n_524),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_601),
.B(n_363),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_638),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_607),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_642),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_645),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_637),
.A2(n_374),
.B1(n_376),
.B2(n_373),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_598),
.B(n_537),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_645),
.Y(n_702)
);

BUFx12f_ASAP7_75t_L g703 ( 
.A(n_615),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_618),
.Y(n_704)
);

NOR3xp33_ASAP7_75t_SL g705 ( 
.A(n_603),
.B(n_386),
.C(n_384),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_605),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_646),
.B(n_362),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_621),
.Y(n_708)
);

HB1xp67_ASAP7_75t_SL g709 ( 
.A(n_624),
.Y(n_709)
);

INVxp67_ASAP7_75t_SL g710 ( 
.A(n_611),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_604),
.B(n_380),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_602),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_604),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_610),
.B(n_533),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_604),
.B(n_381),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_646),
.B(n_364),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_646),
.B(n_366),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_604),
.B(n_383),
.Y(n_718)
);

INVx5_ASAP7_75t_L g719 ( 
.A(n_631),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_604),
.B(n_388),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_600),
.Y(n_721)
);

OR2x6_ASAP7_75t_L g722 ( 
.A(n_624),
.B(n_533),
.Y(n_722)
);

BUFx4f_ASAP7_75t_L g723 ( 
.A(n_635),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_604),
.B(n_543),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_614),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_713),
.B(n_514),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_681),
.A2(n_498),
.B(n_493),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_651),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_724),
.B(n_404),
.Y(n_729)
);

AO32x2_ASAP7_75t_L g730 ( 
.A1(n_670),
.A2(n_532),
.A3(n_514),
.B1(n_19),
.B2(n_17),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_657),
.B(n_414),
.Y(n_731)
);

OAI21xp5_ASAP7_75t_L g732 ( 
.A1(n_698),
.A2(n_423),
.B(n_421),
.Y(n_732)
);

O2A1O1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_661),
.A2(n_434),
.B(n_437),
.C(n_431),
.Y(n_733)
);

CKINVDCx11_ASAP7_75t_R g734 ( 
.A(n_656),
.Y(n_734)
);

O2A1O1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_707),
.A2(n_443),
.B(n_448),
.C(n_440),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_676),
.B(n_692),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_696),
.B(n_389),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_673),
.B(n_390),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_721),
.Y(n_739)
);

HAxp5_ASAP7_75t_L g740 ( 
.A(n_671),
.B(n_392),
.CON(n_740),
.SN(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_723),
.B(n_394),
.Y(n_741)
);

NOR3xp33_ASAP7_75t_SL g742 ( 
.A(n_693),
.B(n_401),
.C(n_396),
.Y(n_742)
);

A2O1A1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_716),
.A2(n_398),
.B(n_400),
.C(n_395),
.Y(n_743)
);

OR2x6_ASAP7_75t_L g744 ( 
.A(n_665),
.B(n_682),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_714),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_717),
.A2(n_403),
.B1(n_406),
.B2(n_402),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_702),
.A2(n_463),
.B(n_98),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_685),
.B(n_407),
.Y(n_748)
);

NAND3xp33_ASAP7_75t_L g749 ( 
.A(n_672),
.B(n_410),
.C(n_405),
.Y(n_749)
);

BUFx8_ASAP7_75t_SL g750 ( 
.A(n_678),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_655),
.A2(n_502),
.B(n_500),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_694),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_SL g753 ( 
.A(n_712),
.B(n_430),
.C(n_419),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_658),
.B(n_688),
.Y(n_754)
);

O2A1O1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_654),
.A2(n_411),
.B(n_416),
.C(n_409),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_R g756 ( 
.A(n_653),
.B(n_425),
.Y(n_756)
);

O2A1O1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_652),
.A2(n_438),
.B(n_442),
.C(n_428),
.Y(n_757)
);

OR2x6_ASAP7_75t_SL g758 ( 
.A(n_706),
.B(n_446),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_699),
.A2(n_451),
.B(n_450),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_660),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_710),
.B(n_452),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_714),
.A2(n_457),
.B(n_458),
.C(n_455),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_683),
.A2(n_461),
.B(n_465),
.C(n_462),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_725),
.Y(n_764)
);

NOR2x1_ASAP7_75t_L g765 ( 
.A(n_659),
.B(n_466),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_691),
.B(n_467),
.Y(n_766)
);

BUFx4f_ASAP7_75t_L g767 ( 
.A(n_659),
.Y(n_767)
);

NAND2x1p5_ASAP7_75t_L g768 ( 
.A(n_687),
.B(n_97),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_697),
.A2(n_474),
.B(n_469),
.Y(n_769)
);

AO32x2_ASAP7_75t_L g770 ( 
.A1(n_708),
.A2(n_21),
.A3(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_649),
.B(n_100),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_669),
.Y(n_772)
);

AND2x6_ASAP7_75t_L g773 ( 
.A(n_704),
.B(n_103),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_711),
.B(n_715),
.Y(n_774)
);

A2O1A1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_650),
.A2(n_23),
.B(n_20),
.C(n_22),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_664),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_722),
.B(n_24),
.Y(n_777)
);

A2O1A1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_666),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_649),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_779)
);

OR2x2_ASAP7_75t_SL g780 ( 
.A(n_677),
.B(n_28),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_680),
.B(n_31),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_718),
.B(n_32),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_663),
.Y(n_783)
);

NAND2x1p5_ASAP7_75t_L g784 ( 
.A(n_689),
.B(n_108),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_722),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_680),
.B(n_33),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_709),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_695),
.A2(n_36),
.B(n_33),
.C(n_35),
.Y(n_788)
);

BUFx8_ASAP7_75t_L g789 ( 
.A(n_703),
.Y(n_789)
);

O2A1O1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_690),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_790)
);

AND2x2_ASAP7_75t_SL g791 ( 
.A(n_701),
.B(n_39),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_719),
.B(n_111),
.Y(n_792)
);

OAI22x1_ASAP7_75t_L g793 ( 
.A1(n_719),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_719),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_674),
.B(n_40),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_679),
.B(n_44),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_667),
.A2(n_121),
.B(n_120),
.Y(n_797)
);

CKINVDCx14_ASAP7_75t_R g798 ( 
.A(n_648),
.Y(n_798)
);

CKINVDCx14_ASAP7_75t_R g799 ( 
.A(n_648),
.Y(n_799)
);

OR2x4_ASAP7_75t_L g800 ( 
.A(n_705),
.B(n_668),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_675),
.B(n_47),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_668),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_R g803 ( 
.A(n_686),
.B(n_123),
.Y(n_803)
);

NAND3xp33_ASAP7_75t_L g804 ( 
.A(n_700),
.B(n_48),
.C(n_49),
.Y(n_804)
);

BUFx12f_ASAP7_75t_L g805 ( 
.A(n_656),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_651),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_665),
.B(n_127),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_681),
.A2(n_130),
.B(n_128),
.Y(n_808)
);

CKINVDCx8_ASAP7_75t_R g809 ( 
.A(n_678),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_713),
.B(n_51),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_713),
.B(n_132),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_723),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_723),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_681),
.B(n_52),
.Y(n_814)
);

INVx4_ASAP7_75t_L g815 ( 
.A(n_723),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_681),
.B(n_53),
.Y(n_816)
);

NAND3xp33_ASAP7_75t_SL g817 ( 
.A(n_720),
.B(n_53),
.C(n_54),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_681),
.A2(n_138),
.B(n_136),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_651),
.Y(n_819)
);

O2A1O1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_670),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_820)
);

INVx8_ASAP7_75t_L g821 ( 
.A(n_659),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_651),
.Y(n_822)
);

NAND2x1p5_ASAP7_75t_L g823 ( 
.A(n_665),
.B(n_140),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_713),
.A2(n_143),
.B1(n_146),
.B2(n_142),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_SL g825 ( 
.A(n_720),
.B(n_58),
.C(n_59),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_SL g826 ( 
.A1(n_662),
.A2(n_151),
.B(n_152),
.C(n_150),
.Y(n_826)
);

O2A1O1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_670),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_827)
);

NOR2xp67_ASAP7_75t_L g828 ( 
.A(n_713),
.B(n_153),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_723),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_681),
.A2(n_162),
.B(n_160),
.Y(n_830)
);

AOI221xp5_ASAP7_75t_L g831 ( 
.A1(n_670),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.C(n_64),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_665),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_651),
.Y(n_833)
);

A2O1A1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_720),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_653),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_653),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_713),
.B(n_65),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_713),
.B(n_164),
.Y(n_838)
);

AO31x2_ASAP7_75t_L g839 ( 
.A1(n_684),
.A2(n_69),
.A3(n_67),
.B(n_68),
.Y(n_839)
);

INVx8_ASAP7_75t_L g840 ( 
.A(n_821),
.Y(n_840)
);

CKINVDCx16_ASAP7_75t_R g841 ( 
.A(n_772),
.Y(n_841)
);

INVx8_ASAP7_75t_L g842 ( 
.A(n_821),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_760),
.B(n_166),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_739),
.Y(n_844)
);

INVx6_ASAP7_75t_L g845 ( 
.A(n_812),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_728),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_794),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_744),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_744),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_813),
.Y(n_850)
);

NOR2x1_ASAP7_75t_L g851 ( 
.A(n_815),
.B(n_832),
.Y(n_851)
);

CKINVDCx11_ASAP7_75t_R g852 ( 
.A(n_805),
.Y(n_852)
);

AO21x2_ASAP7_75t_L g853 ( 
.A1(n_732),
.A2(n_174),
.B(n_172),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_794),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_813),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_806),
.Y(n_856)
);

OAI21x1_ASAP7_75t_L g857 ( 
.A1(n_747),
.A2(n_177),
.B(n_176),
.Y(n_857)
);

AOI22x1_ASAP7_75t_L g858 ( 
.A1(n_727),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_819),
.Y(n_859)
);

INVx8_ASAP7_75t_L g860 ( 
.A(n_829),
.Y(n_860)
);

BUFx2_ASAP7_75t_SL g861 ( 
.A(n_829),
.Y(n_861)
);

AND2x6_ASAP7_75t_L g862 ( 
.A(n_771),
.B(n_179),
.Y(n_862)
);

CKINVDCx14_ASAP7_75t_R g863 ( 
.A(n_798),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_745),
.Y(n_864)
);

BUFx2_ASAP7_75t_SL g865 ( 
.A(n_764),
.Y(n_865)
);

INVx1_ASAP7_75t_SL g866 ( 
.A(n_787),
.Y(n_866)
);

OR2x6_ASAP7_75t_L g867 ( 
.A(n_783),
.B(n_72),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_814),
.A2(n_183),
.B(n_181),
.Y(n_868)
);

OAI21x1_ASAP7_75t_SL g869 ( 
.A1(n_788),
.A2(n_185),
.B(n_184),
.Y(n_869)
);

INVx1_ASAP7_75t_SL g870 ( 
.A(n_777),
.Y(n_870)
);

CKINVDCx16_ASAP7_75t_R g871 ( 
.A(n_799),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_737),
.B(n_73),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_750),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_SL g874 ( 
.A(n_831),
.B(n_73),
.C(n_74),
.Y(n_874)
);

AO21x2_ASAP7_75t_L g875 ( 
.A1(n_816),
.A2(n_189),
.B(n_187),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_754),
.B(n_74),
.Y(n_876)
);

CKINVDCx14_ASAP7_75t_R g877 ( 
.A(n_734),
.Y(n_877)
);

AOI21xp33_ASAP7_75t_L g878 ( 
.A1(n_774),
.A2(n_75),
.B(n_76),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_822),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_783),
.Y(n_880)
);

BUFx4f_ASAP7_75t_SL g881 ( 
.A(n_800),
.Y(n_881)
);

CKINVDCx16_ASAP7_75t_R g882 ( 
.A(n_802),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_833),
.Y(n_883)
);

AO21x2_ASAP7_75t_L g884 ( 
.A1(n_731),
.A2(n_826),
.B(n_729),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_752),
.B(n_76),
.Y(n_885)
);

AOI22x1_ASAP7_75t_L g886 ( 
.A1(n_808),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_736),
.A2(n_193),
.B(n_192),
.Y(n_887)
);

BUFx12f_ASAP7_75t_L g888 ( 
.A(n_835),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_785),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_795),
.Y(n_890)
);

INVx5_ASAP7_75t_L g891 ( 
.A(n_773),
.Y(n_891)
);

INVxp67_ASAP7_75t_SL g892 ( 
.A(n_776),
.Y(n_892)
);

AO21x2_ASAP7_75t_L g893 ( 
.A1(n_743),
.A2(n_196),
.B(n_195),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_809),
.Y(n_894)
);

INVx6_ASAP7_75t_L g895 ( 
.A(n_789),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_836),
.Y(n_896)
);

AO21x2_ASAP7_75t_L g897 ( 
.A1(n_828),
.A2(n_199),
.B(n_198),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_767),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_807),
.Y(n_899)
);

BUFx2_ASAP7_75t_SL g900 ( 
.A(n_773),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_781),
.Y(n_901)
);

INVx5_ASAP7_75t_L g902 ( 
.A(n_773),
.Y(n_902)
);

INVx1_ASAP7_75t_SL g903 ( 
.A(n_756),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_738),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_768),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_765),
.B(n_206),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_786),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_758),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_766),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_796),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_823),
.Y(n_911)
);

INVx8_ASAP7_75t_L g912 ( 
.A(n_740),
.Y(n_912)
);

INVx4_ASAP7_75t_L g913 ( 
.A(n_784),
.Y(n_913)
);

NAND2x1p5_ASAP7_75t_L g914 ( 
.A(n_792),
.B(n_207),
.Y(n_914)
);

BUFx2_ASAP7_75t_R g915 ( 
.A(n_801),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_791),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_818),
.A2(n_266),
.B(n_311),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_742),
.B(n_209),
.Y(n_918)
);

INVxp67_ASAP7_75t_SL g919 ( 
.A(n_810),
.Y(n_919)
);

BUFx4f_ASAP7_75t_L g920 ( 
.A(n_803),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_839),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_726),
.B(n_80),
.Y(n_922)
);

NAND2x1p5_ASAP7_75t_L g923 ( 
.A(n_811),
.B(n_212),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_761),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_770),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_780),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_770),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_748),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_749),
.B(n_81),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_753),
.Y(n_930)
);

BUFx2_ASAP7_75t_SL g931 ( 
.A(n_838),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_804),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_741),
.B(n_213),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_779),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_837),
.Y(n_935)
);

BUFx12f_ASAP7_75t_L g936 ( 
.A(n_793),
.Y(n_936)
);

INVx5_ASAP7_75t_L g937 ( 
.A(n_824),
.Y(n_937)
);

INVxp67_ASAP7_75t_L g938 ( 
.A(n_782),
.Y(n_938)
);

NOR2x1_ASAP7_75t_R g939 ( 
.A(n_730),
.B(n_81),
.Y(n_939)
);

AOI22x1_ASAP7_75t_L g940 ( 
.A1(n_830),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_940)
);

INVx8_ASAP7_75t_L g941 ( 
.A(n_762),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_775),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_746),
.B(n_82),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_817),
.Y(n_944)
);

NOR2x1_ASAP7_75t_R g945 ( 
.A(n_730),
.B(n_825),
.Y(n_945)
);

OAI21x1_ASAP7_75t_SL g946 ( 
.A1(n_820),
.A2(n_262),
.B(n_310),
.Y(n_946)
);

BUFx2_ASAP7_75t_SL g947 ( 
.A(n_797),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_755),
.A2(n_257),
.B(n_308),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_827),
.Y(n_949)
);

INVxp67_ASAP7_75t_SL g950 ( 
.A(n_790),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_834),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_778),
.B(n_769),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_757),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_751),
.Y(n_954)
);

BUFx4f_ASAP7_75t_SL g955 ( 
.A(n_888),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_859),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_860),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_860),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_859),
.Y(n_959)
);

BUFx2_ASAP7_75t_SL g960 ( 
.A(n_896),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_846),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_904),
.B(n_759),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_856),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_SL g964 ( 
.A1(n_916),
.A2(n_733),
.B1(n_735),
.B2(n_763),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_844),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_879),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_883),
.Y(n_967)
);

INVx4_ASAP7_75t_SL g968 ( 
.A(n_845),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_873),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_845),
.Y(n_970)
);

AO21x2_ASAP7_75t_L g971 ( 
.A1(n_921),
.A2(n_268),
.B(n_306),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_938),
.B(n_85),
.Y(n_972)
);

OAI22xp33_ASAP7_75t_L g973 ( 
.A1(n_916),
.A2(n_949),
.B1(n_935),
.B2(n_944),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_847),
.Y(n_974)
);

OAI22xp33_ASAP7_75t_L g975 ( 
.A1(n_920),
.A2(n_910),
.B1(n_922),
.B2(n_919),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_SL g976 ( 
.A1(n_936),
.A2(n_87),
.B1(n_214),
.B2(n_215),
.Y(n_976)
);

INVx1_ASAP7_75t_SL g977 ( 
.A(n_861),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_909),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_978)
);

INVx5_ASAP7_75t_SL g979 ( 
.A(n_847),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_892),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_937),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_899),
.B(n_313),
.Y(n_982)
);

BUFx8_ASAP7_75t_L g983 ( 
.A(n_850),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_901),
.A2(n_226),
.B(n_227),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_951),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_891),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_907),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_851),
.B(n_228),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_934),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_924),
.B(n_229),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_937),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_943),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_954),
.Y(n_993)
);

NAND2x1p5_ASAP7_75t_L g994 ( 
.A(n_850),
.B(n_238),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_932),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_840),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_942),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_954),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_952),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_870),
.B(n_240),
.Y(n_1000)
);

OAI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_874),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_857),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_927),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_890),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_890),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_872),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_SL g1007 ( 
.A1(n_876),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_1007)
);

CKINVDCx20_ASAP7_75t_R g1008 ( 
.A(n_852),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_854),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_950),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_840),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_885),
.B(n_273),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_889),
.Y(n_1013)
);

BUFx2_ASAP7_75t_R g1014 ( 
.A(n_861),
.Y(n_1014)
);

INVx6_ASAP7_75t_L g1015 ( 
.A(n_842),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_911),
.Y(n_1016)
);

AO21x2_ASAP7_75t_L g1017 ( 
.A1(n_948),
.A2(n_884),
.B(n_868),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_880),
.B(n_280),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_841),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_843),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_848),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_855),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_905),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_877),
.Y(n_1024)
);

BUFx2_ASAP7_75t_R g1025 ( 
.A(n_898),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_903),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_937),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_1027)
);

INVx6_ASAP7_75t_L g1028 ( 
.A(n_854),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_905),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_880),
.B(n_305),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_SL g1031 ( 
.A1(n_878),
.A2(n_286),
.B(n_288),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_905),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_931),
.A2(n_902),
.B1(n_953),
.B2(n_928),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_887),
.A2(n_289),
.B(n_290),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_917),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_933),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_923),
.A2(n_295),
.B(n_296),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_933),
.A2(n_941),
.B1(n_912),
.B2(n_930),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_925),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_925),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_849),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_900),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_900),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_941),
.A2(n_300),
.B1(n_302),
.B2(n_304),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_965),
.Y(n_1045)
);

NOR3xp33_ASAP7_75t_SL g1046 ( 
.A(n_975),
.B(n_882),
.C(n_871),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_R g1047 ( 
.A(n_1019),
.B(n_863),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_1026),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_1004),
.B(n_929),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_R g1050 ( 
.A(n_969),
.B(n_894),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_956),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_973),
.A2(n_1038),
.B1(n_1010),
.B2(n_962),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_956),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_1008),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_970),
.Y(n_1055)
);

CKINVDCx16_ASAP7_75t_R g1056 ( 
.A(n_1024),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_1005),
.B(n_926),
.Y(n_1057)
);

NOR3xp33_ASAP7_75t_L g1058 ( 
.A(n_976),
.B(n_1031),
.C(n_1033),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_987),
.B(n_945),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1020),
.A2(n_915),
.B1(n_902),
.B2(n_913),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_957),
.Y(n_1061)
);

AO31x2_ASAP7_75t_L g1062 ( 
.A1(n_1002),
.A2(n_947),
.A3(n_940),
.B(n_886),
.Y(n_1062)
);

CKINVDCx11_ASAP7_75t_R g1063 ( 
.A(n_968),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_1013),
.B(n_866),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_SL g1065 ( 
.A1(n_1007),
.A2(n_906),
.B1(n_886),
.B2(n_940),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_955),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_999),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_R g1068 ( 
.A(n_958),
.B(n_881),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1012),
.B(n_918),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_960),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_1001),
.A2(n_972),
.B(n_1034),
.C(n_946),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_995),
.B(n_939),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_959),
.Y(n_1073)
);

AO31x2_ASAP7_75t_L g1074 ( 
.A1(n_1002),
.A2(n_947),
.A3(n_869),
.B(n_853),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_R g1075 ( 
.A(n_1015),
.B(n_880),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_983),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_1021),
.Y(n_1077)
);

CKINVDCx16_ASAP7_75t_R g1078 ( 
.A(n_996),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_983),
.Y(n_1079)
);

NAND2xp33_ASAP7_75t_R g1080 ( 
.A(n_986),
.B(n_867),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_968),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_1015),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_1041),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_1035),
.A2(n_869),
.A3(n_893),
.B(n_875),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_1025),
.Y(n_1085)
);

OR2x6_ASAP7_75t_L g1086 ( 
.A(n_994),
.B(n_865),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_R g1087 ( 
.A(n_1011),
.B(n_864),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_980),
.B(n_862),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_SL g1089 ( 
.A1(n_1037),
.A2(n_858),
.B1(n_908),
.B2(n_914),
.Y(n_1089)
);

CKINVDCx8_ASAP7_75t_R g1090 ( 
.A(n_1018),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_961),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_1028),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_1030),
.B(n_897),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_1028),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_1000),
.B(n_895),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_979),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_1014),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_963),
.B(n_966),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_967),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_1022),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1023),
.B(n_1029),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_982),
.B(n_1032),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_993),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_989),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_989),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_998),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_SL g1107 ( 
.A1(n_984),
.A2(n_981),
.B1(n_991),
.B2(n_1027),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_985),
.B(n_997),
.Y(n_1108)
);

CKINVDCx16_ASAP7_75t_R g1109 ( 
.A(n_977),
.Y(n_1109)
);

OR2x2_ASAP7_75t_L g1110 ( 
.A(n_1049),
.B(n_1039),
.Y(n_1110)
);

OR2x2_ASAP7_75t_L g1111 ( 
.A(n_1045),
.B(n_1039),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1091),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1058),
.A2(n_1036),
.B1(n_992),
.B2(n_1017),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1104),
.Y(n_1114)
);

INVxp67_ASAP7_75t_L g1115 ( 
.A(n_1083),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1067),
.B(n_1040),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1051),
.Y(n_1117)
);

INVx2_ASAP7_75t_R g1118 ( 
.A(n_1105),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1053),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1073),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1067),
.B(n_1003),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_1103),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_1090),
.Y(n_1123)
);

NAND2x1_ASAP7_75t_L g1124 ( 
.A(n_1086),
.B(n_1042),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1103),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_1086),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1069),
.B(n_1043),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1072),
.B(n_988),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1098),
.Y(n_1129)
);

OR2x2_ASAP7_75t_L g1130 ( 
.A(n_1077),
.B(n_990),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_1106),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_1064),
.B(n_1016),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1102),
.B(n_964),
.Y(n_1133)
);

OAI211xp5_ASAP7_75t_L g1134 ( 
.A1(n_1065),
.A2(n_1006),
.B(n_1044),
.C(n_978),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_1099),
.B(n_971),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1108),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1052),
.B(n_979),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1059),
.B(n_974),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1057),
.B(n_1009),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_1109),
.B(n_971),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1129),
.B(n_1136),
.Y(n_1141)
);

NOR3xp33_ASAP7_75t_L g1142 ( 
.A(n_1134),
.B(n_1089),
.C(n_1071),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1127),
.B(n_1046),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1114),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1117),
.Y(n_1145)
);

OR2x2_ASAP7_75t_L g1146 ( 
.A(n_1125),
.B(n_1088),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1119),
.Y(n_1147)
);

INVx4_ASAP7_75t_L g1148 ( 
.A(n_1126),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1120),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1115),
.B(n_1093),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_1133),
.B(n_1107),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1110),
.B(n_1101),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1112),
.B(n_1062),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_1131),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1122),
.B(n_1125),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1121),
.B(n_1074),
.Y(n_1156)
);

BUFx2_ASAP7_75t_SL g1157 ( 
.A(n_1123),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1122),
.B(n_1101),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1135),
.B(n_1074),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1121),
.B(n_1084),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1159),
.B(n_1135),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1159),
.B(n_1116),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1144),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_1155),
.B(n_1150),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_1154),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1149),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1149),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1156),
.B(n_1118),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1153),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1145),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1141),
.B(n_1146),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1147),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1152),
.B(n_1111),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1166),
.Y(n_1174)
);

OAI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1173),
.A2(n_1151),
.B1(n_1137),
.B2(n_1140),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1167),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1170),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1172),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1164),
.B(n_1151),
.Y(n_1179)
);

NOR2xp67_ASAP7_75t_L g1180 ( 
.A(n_1163),
.B(n_1148),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1165),
.A2(n_1142),
.B1(n_1113),
.B2(n_1128),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1161),
.A2(n_1113),
.B(n_1060),
.C(n_1124),
.Y(n_1182)
);

OAI32xp33_ASAP7_75t_L g1183 ( 
.A1(n_1169),
.A2(n_1080),
.A3(n_1143),
.B1(n_1158),
.B2(n_1130),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1162),
.B(n_1160),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1174),
.Y(n_1185)
);

CKINVDCx16_ASAP7_75t_R g1186 ( 
.A(n_1179),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1182),
.A2(n_1171),
.B(n_1168),
.Y(n_1187)
);

AOI31xp33_ASAP7_75t_L g1188 ( 
.A1(n_1181),
.A2(n_1085),
.A3(n_1070),
.B(n_1097),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1184),
.B(n_1161),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1176),
.Y(n_1190)
);

AOI21xp33_ASAP7_75t_SL g1191 ( 
.A1(n_1175),
.A2(n_1056),
.B(n_1054),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1177),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1186),
.B(n_1175),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1192),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_SL g1195 ( 
.A(n_1187),
.B(n_1183),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1191),
.B(n_1076),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1185),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1194),
.Y(n_1198)
);

NAND2x1p5_ASAP7_75t_L g1199 ( 
.A(n_1193),
.B(n_1180),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1197),
.Y(n_1200)
);

AOI221xp5_ASAP7_75t_L g1201 ( 
.A1(n_1195),
.A2(n_1188),
.B1(n_1181),
.B2(n_1190),
.C(n_1178),
.Y(n_1201)
);

NOR3xp33_ASAP7_75t_SL g1202 ( 
.A(n_1196),
.B(n_1079),
.C(n_1078),
.Y(n_1202)
);

AOI211xp5_ASAP7_75t_L g1203 ( 
.A1(n_1195),
.A2(n_1095),
.B(n_1188),
.C(n_1123),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1201),
.B(n_1189),
.Y(n_1204)
);

OAI211xp5_ASAP7_75t_SL g1205 ( 
.A1(n_1203),
.A2(n_1132),
.B(n_1055),
.C(n_1063),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1199),
.A2(n_1048),
.B(n_1066),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1204),
.Y(n_1207)
);

NAND2xp33_ASAP7_75t_SL g1208 ( 
.A(n_1205),
.B(n_1202),
.Y(n_1208)
);

NOR2x1_ASAP7_75t_L g1209 ( 
.A(n_1207),
.B(n_1206),
.Y(n_1209)
);

NAND3xp33_ASAP7_75t_L g1210 ( 
.A(n_1209),
.B(n_1208),
.C(n_1200),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_1210),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_R g1212 ( 
.A(n_1210),
.B(n_1096),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1212),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1211),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1214),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1213),
.A2(n_1198),
.B1(n_1123),
.B2(n_1157),
.Y(n_1216)
);

AO22x2_ASAP7_75t_L g1217 ( 
.A1(n_1215),
.A2(n_1081),
.B1(n_1082),
.B2(n_1047),
.Y(n_1217)
);

NOR2xp67_ASAP7_75t_L g1218 ( 
.A(n_1216),
.B(n_1061),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1217),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1218),
.Y(n_1220)
);

OR2x6_ASAP7_75t_L g1221 ( 
.A(n_1219),
.B(n_1061),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1220),
.B(n_1100),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_R g1223 ( 
.A1(n_1221),
.A2(n_1050),
.B1(n_1068),
.B2(n_1087),
.Y(n_1223)
);

AOI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1222),
.A2(n_1094),
.B1(n_1092),
.B2(n_1138),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1224),
.B(n_1139),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_SL g1226 ( 
.A1(n_1225),
.A2(n_1223),
.B1(n_1092),
.B2(n_1075),
.Y(n_1226)
);


endmodule