module fake_jpeg_5611_n_294 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_294);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_219;
wire n_70;
wire n_130;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_107;
wire n_39;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx8_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_43),
.B(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_0),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_22),
.B(n_1),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_25),
.B(n_2),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_47),
.B(n_57),
.Y(n_84)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_58),
.B1(n_59),
.B2(n_64),
.Y(n_70)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_55),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_22),
.B(n_2),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g85 ( 
.A(n_54),
.Y(n_85)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_28),
.B(n_2),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_33),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_3),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_61),
.B(n_63),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_5),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_68),
.Y(n_91)
);

BUFx4f_ASAP7_75t_SL g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_74),
.B(n_80),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_27),
.B1(n_26),
.B2(n_18),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_79),
.B1(n_83),
.B2(n_87),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_107),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_58),
.A2(n_27),
.B1(n_26),
.B2(n_18),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

OA22x2_ASAP7_75t_SL g81 ( 
.A1(n_54),
.A2(n_26),
.B1(n_24),
.B2(n_27),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g116 ( 
.A(n_81),
.B(n_24),
.Y(n_116)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_82),
.B(n_86),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_59),
.A2(n_18),
.B1(n_31),
.B2(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_31),
.B1(n_49),
.B2(n_55),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_94),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_45),
.A2(n_31),
.B1(n_35),
.B2(n_40),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_90),
.A2(n_93),
.B1(n_106),
.B2(n_108),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_61),
.A2(n_35),
.B1(n_36),
.B2(n_28),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_102),
.Y(n_137)
);

CKINVDCx6p67_ASAP7_75t_R g96 ( 
.A(n_50),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_96),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_51),
.A2(n_36),
.B1(n_29),
.B2(n_33),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_41),
.B1(n_42),
.B2(n_9),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_29),
.B1(n_38),
.B2(n_30),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_39),
.B1(n_32),
.B2(n_24),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_38),
.Y(n_101)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_50),
.A2(n_30),
.B1(n_37),
.B2(n_24),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_5),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_114),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_93),
.B(n_90),
.C(n_85),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_111),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_39),
.B1(n_32),
.B2(n_24),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_138),
.B1(n_144),
.B2(n_108),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_83),
.B(n_79),
.C(n_75),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_53),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_122),
.Y(n_149)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_85),
.Y(n_119)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_89),
.B(n_5),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_120),
.B(n_126),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_53),
.Y(n_122)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_125),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_80),
.A2(n_39),
.B1(n_41),
.B2(n_9),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_76),
.B(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_127),
.B(n_140),
.Y(n_164)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_134),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_53),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_133),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_69),
.B(n_52),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_7),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_95),
.A2(n_41),
.B1(n_42),
.B2(n_9),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_91),
.A2(n_41),
.B(n_42),
.C(n_10),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_139),
.A2(n_141),
.B1(n_104),
.B2(n_71),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_96),
.B(n_6),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_87),
.A2(n_41),
.B1(n_7),
.B2(n_10),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_6),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_98),
.B(n_11),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_69),
.B(n_6),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_98),
.Y(n_162)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_152),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_153),
.B1(n_110),
.B2(n_139),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_148),
.B(n_143),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_151),
.A2(n_169),
.B1(n_172),
.B2(n_141),
.Y(n_194)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

OAI22x1_ASAP7_75t_SL g153 ( 
.A1(n_116),
.A2(n_70),
.B1(n_100),
.B2(n_77),
.Y(n_153)
);

BUFx8_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_154),
.Y(n_179)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_157),
.Y(n_191)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_70),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_163),
.C(n_121),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_162),
.B(n_118),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_103),
.C(n_104),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_103),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_166),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_98),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_173),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_71),
.B1(n_100),
.B2(n_13),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_7),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_177),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_181),
.Y(n_207)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_170),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_182),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_151),
.B1(n_169),
.B2(n_161),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_111),
.Y(n_185)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_192),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_177),
.B(n_127),
.Y(n_188)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_165),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_197),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_143),
.B(n_115),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_195),
.B(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_193),
.B(n_198),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_153),
.B1(n_164),
.B2(n_166),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_145),
.B(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_121),
.Y(n_199)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_154),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_202),
.B(n_204),
.Y(n_217)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_159),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_223),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_163),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_227),
.C(n_197),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_216),
.A2(n_221),
.B1(n_224),
.B2(n_215),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_204),
.B(n_168),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_178),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_194),
.A2(n_139),
.B1(n_152),
.B2(n_167),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_188),
.B1(n_195),
.B2(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_184),
.A2(n_146),
.B1(n_158),
.B2(n_171),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_183),
.A2(n_154),
.B(n_173),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_187),
.A2(n_180),
.B1(n_181),
.B2(n_183),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_199),
.B(n_139),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_206),
.B(n_200),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_235),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_236),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_231),
.A2(n_201),
.B1(n_178),
.B2(n_158),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_192),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_238),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g235 ( 
.A(n_206),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_186),
.C(n_205),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_205),
.Y(n_237)
);

AOI321xp33_ASAP7_75t_L g258 ( 
.A1(n_237),
.A2(n_239),
.A3(n_179),
.B1(n_155),
.B2(n_191),
.C(n_113),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_182),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_L g239 ( 
.A1(n_212),
.A2(n_214),
.B(n_215),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_193),
.C(n_200),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_242),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_208),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_201),
.C(n_202),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_196),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_212),
.A2(n_198),
.B1(n_196),
.B2(n_179),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_217),
.B(n_210),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_245),
.B(n_207),
.Y(n_246)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_247),
.B(n_257),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_228),
.A2(n_216),
.B1(n_221),
.B2(n_211),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_251),
.B1(n_134),
.B2(n_124),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_232),
.A2(n_219),
.B1(n_224),
.B2(n_227),
.Y(n_251)
);

AOI322xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_233),
.A3(n_228),
.B1(n_237),
.B2(n_230),
.C1(n_231),
.C2(n_236),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_258),
.Y(n_269)
);

OAI21x1_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_223),
.B(n_154),
.Y(n_255)
);

O2A1O1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_255),
.A2(n_234),
.B(n_243),
.C(n_244),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_226),
.B1(n_113),
.B2(n_203),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_262),
.B1(n_248),
.B2(n_247),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_240),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_269),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_191),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_261),
.A2(n_266),
.B(n_251),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_246),
.B(n_130),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_268),
.C(n_256),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_226),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_255),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_254),
.B(n_11),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_249),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_270),
.B(n_277),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_271),
.A2(n_267),
.B1(n_263),
.B2(n_259),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_272),
.B(n_276),
.Y(n_282)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_273),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_274),
.A2(n_275),
.B(n_266),
.Y(n_281)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_265),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_258),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_280),
.A2(n_281),
.B(n_283),
.Y(n_287)
);

XOR2x2_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_261),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_280),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_285),
.B(n_286),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_250),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_283),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_282),
.B(n_272),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_288),
.A2(n_279),
.B(n_15),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_291),
.B(n_14),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_114),
.C(n_16),
.Y(n_291)
);

AO21x2_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_14),
.B(n_17),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_292),
.B(n_293),
.Y(n_294)
);


endmodule