module fake_jpeg_21525_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_16),
.B(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_15),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_17),
.B1(n_25),
.B2(n_21),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_45),
.A2(n_56),
.B1(n_63),
.B2(n_26),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_17),
.B1(n_25),
.B2(n_21),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_46),
.A2(n_33),
.B1(n_29),
.B2(n_16),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g88 ( 
.A(n_50),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_28),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_17),
.B1(n_25),
.B2(n_20),
.Y(n_56)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_21),
.B1(n_42),
.B2(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_70),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_68),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_53),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_72),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_53),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_75),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_44),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_76),
.B(n_18),
.C(n_1),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_47),
.B(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_85),
.Y(n_106)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_36),
.B1(n_20),
.B2(n_23),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_82),
.B1(n_103),
.B2(n_105),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_35),
.B(n_16),
.C(n_28),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_38),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_84),
.A2(n_38),
.B(n_19),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_34),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_87),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_24),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_48),
.A2(n_34),
.B1(n_22),
.B2(n_24),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_90),
.A2(n_100),
.B1(n_102),
.B2(n_19),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_93),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_95),
.Y(n_115)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_48),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_98),
.B1(n_35),
.B2(n_38),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_24),
.B1(n_22),
.B2(n_27),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_36),
.B1(n_20),
.B2(n_23),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_26),
.B1(n_19),
.B2(n_30),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_53),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_57),
.B(n_31),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_52),
.A2(n_36),
.B1(n_23),
.B2(n_27),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_109),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_84),
.A2(n_27),
.B1(n_33),
.B2(n_26),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_35),
.B1(n_29),
.B2(n_32),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_118),
.B1(n_120),
.B2(n_122),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_71),
.A2(n_35),
.B1(n_29),
.B2(n_32),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_65),
.A2(n_35),
.B1(n_28),
.B2(n_32),
.Y(n_120)
);

AO21x2_ASAP7_75t_L g122 ( 
.A1(n_76),
.A2(n_38),
.B(n_19),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_67),
.B(n_89),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_80),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_70),
.A2(n_19),
.B1(n_38),
.B2(n_30),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_99),
.B1(n_96),
.B2(n_93),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_19),
.B1(n_18),
.B2(n_38),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_133),
.A2(n_135),
.B1(n_73),
.B2(n_64),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_92),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_84),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_137),
.B(n_157),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_139),
.B(n_142),
.Y(n_195)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_146),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_136),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_150),
.B1(n_159),
.B2(n_127),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_109),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_91),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_108),
.A2(n_76),
.B(n_102),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_148),
.A2(n_156),
.B(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_108),
.A2(n_101),
.B1(n_82),
.B2(n_68),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_151),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_136),
.B(n_69),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_155),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_158),
.B1(n_163),
.B2(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_154),
.Y(n_199)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_121),
.Y(n_157)
);

OAI22x1_ASAP7_75t_SL g158 ( 
.A1(n_112),
.A2(n_88),
.B1(n_92),
.B2(n_75),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_112),
.A2(n_78),
.B1(n_64),
.B2(n_79),
.Y(n_159)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_165),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_121),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_120),
.Y(n_175)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_117),
.B(n_88),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_167),
.Y(n_190)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_117),
.C(n_125),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_170),
.C(n_180),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_164),
.C(n_156),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_134),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_173),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_160),
.B(n_138),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_174),
.A2(n_181),
.B1(n_198),
.B2(n_0),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_177),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_118),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_111),
.Y(n_178)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_132),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_122),
.B1(n_113),
.B2(n_115),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_122),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_186),
.C(n_192),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_163),
.A2(n_122),
.B1(n_119),
.B2(n_115),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_184),
.A2(n_126),
.B1(n_110),
.B2(n_80),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_122),
.Y(n_185)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_122),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_119),
.Y(n_191)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_107),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_78),
.C(n_74),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_154),
.B(n_143),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_162),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_145),
.A2(n_126),
.B1(n_110),
.B2(n_123),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g201 ( 
.A1(n_185),
.A2(n_146),
.B(n_161),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_194),
.B(n_193),
.Y(n_238)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_196),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_212),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_196),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_211),
.B(n_214),
.Y(n_242)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_220),
.Y(n_244)
);

NAND3xp33_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_151),
.C(n_149),
.Y(n_214)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_218),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_234)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_7),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_176),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_223),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_177),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_178),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_199),
.Y(n_227)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_220),
.A2(n_174),
.B1(n_183),
.B2(n_186),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_229),
.A2(n_245),
.B1(n_226),
.B2(n_201),
.Y(n_268)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_204),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_171),
.C(n_170),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_241),
.C(n_246),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_189),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_247),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_209),
.A2(n_192),
.B1(n_175),
.B2(n_179),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_237),
.A2(n_240),
.B1(n_221),
.B2(n_208),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_242),
.B(n_239),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_209),
.A2(n_180),
.B1(n_193),
.B2(n_189),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_168),
.C(n_172),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_203),
.A2(n_172),
.B1(n_3),
.B2(n_4),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_8),
.C(n_13),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_8),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_228),
.A2(n_202),
.B(n_203),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_253),
.B(n_257),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_252),
.A2(n_266),
.B1(n_245),
.B2(n_229),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_202),
.B(n_219),
.Y(n_253)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_264),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_233),
.B(n_212),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_256),
.B(n_260),
.Y(n_270)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_210),
.C(n_206),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_261),
.C(n_267),
.Y(n_271)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_259),
.B(n_263),
.Y(n_274)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_205),
.C(n_216),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_241),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_200),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_265),
.Y(n_278)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_231),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_200),
.C(n_201),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_269),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_9),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_244),
.B(n_232),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_273),
.A2(n_268),
.B1(n_253),
.B2(n_269),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_275),
.Y(n_289)
);

NAND3xp33_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_246),
.C(n_249),
.Y(n_277)
);

AOI21x1_ASAP7_75t_L g295 ( 
.A1(n_277),
.A2(n_15),
.B(n_11),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_280),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_237),
.C(n_234),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_258),
.C(n_267),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_234),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_264),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_287),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_292),
.C(n_293),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_281),
.A2(n_251),
.B1(n_250),
.B2(n_230),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_282),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_250),
.C(n_9),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_9),
.C(n_13),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_294),
.A2(n_278),
.B(n_276),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_270),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_298),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_272),
.C(n_284),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_300),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_289),
.A2(n_275),
.B(n_283),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_282),
.C(n_279),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_285),
.C(n_287),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_293),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_305),
.A2(n_300),
.B(n_15),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_306),
.A2(n_310),
.B(n_303),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_304),
.C(n_291),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_SL g310 ( 
.A(n_302),
.B(n_294),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_311),
.A2(n_313),
.B(n_308),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_312),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_315),
.A2(n_309),
.B(n_11),
.Y(n_316)
);

AOI321xp33_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_11),
.A3(n_10),
.B1(n_314),
.B2(n_5),
.C(n_2),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_317),
.Y(n_318)
);

AOI21x1_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_10),
.B(n_4),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_3),
.Y(n_320)
);


endmodule