module fake_ariane_1642_n_1854 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1854);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1854;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1429;
wire n_1324;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_133),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_123),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_100),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_91),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_90),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_101),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_137),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_105),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_78),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_117),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_83),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_56),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_170),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_174),
.Y(n_198)
);

BUFx2_ASAP7_75t_R g199 ( 
.A(n_4),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_53),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_160),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_27),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_125),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_152),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_52),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_140),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_1),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_41),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_30),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_67),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_18),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_14),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_72),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_36),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_156),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_43),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_45),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_39),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_5),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_40),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_26),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_168),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_182),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_44),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_47),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_47),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_179),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_63),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_122),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_89),
.Y(n_232)
);

BUFx8_ASAP7_75t_SL g233 ( 
.A(n_164),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_108),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_24),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_70),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_159),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_161),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_103),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_98),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_145),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_53),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_141),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_111),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_13),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_96),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_36),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_114),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_2),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_95),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_21),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_104),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_21),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_50),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_87),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_4),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_3),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_39),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_135),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_76),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_148),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_146),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_69),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_33),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_180),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_44),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_2),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_54),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_30),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_11),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_99),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_5),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_106),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_175),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_27),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_64),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_56),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_81),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_54),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_121),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_29),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_126),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_124),
.Y(n_283)
);

BUFx5_ASAP7_75t_L g284 ( 
.A(n_1),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_171),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_15),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_113),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_38),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_153),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_110),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_41),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_9),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_19),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_23),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_94),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_130),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_9),
.Y(n_297)
);

BUFx5_ASAP7_75t_L g298 ( 
.A(n_149),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_102),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_10),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_131),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_166),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_32),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_183),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_86),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_29),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_8),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_80),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_62),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_107),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_75),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_37),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_61),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_34),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_154),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_138),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_19),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_150),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_60),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_13),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_181),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_85),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_93),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_147),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_162),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_59),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_0),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_42),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_116),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_176),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_43),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_12),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_24),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_23),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_163),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_127),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_49),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_169),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_84),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_33),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_115),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_71),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_15),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_31),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_6),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_151),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_97),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_34),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_10),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_112),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_17),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_20),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_73),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_58),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_178),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_120),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_3),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_40),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_12),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_61),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_136),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_0),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_48),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_59),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_143),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_16),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_184),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_233),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_213),
.B(n_6),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_245),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_213),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_213),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_218),
.B(n_7),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_213),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_207),
.B(n_7),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_233),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_207),
.B(n_8),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_286),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_328),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_210),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_209),
.Y(n_381)
);

INVxp33_ASAP7_75t_SL g382 ( 
.A(n_209),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_184),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_213),
.B(n_11),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_213),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_214),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_216),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_213),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_226),
.B(n_14),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_220),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_221),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_223),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_284),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_203),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_196),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_226),
.B(n_16),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_203),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_284),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_263),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_228),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_284),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_242),
.Y(n_402)
);

NOR2xp67_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_17),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_251),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_253),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_254),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_248),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_284),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_284),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_203),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_257),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_264),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_269),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_270),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_272),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_196),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_284),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_284),
.Y(n_419)
);

NOR2xp67_ASAP7_75t_L g420 ( 
.A(n_332),
.B(n_18),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_333),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_333),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_344),
.Y(n_423)
);

INVxp33_ASAP7_75t_L g424 ( 
.A(n_195),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_255),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_255),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_277),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_333),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_344),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_203),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_265),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_249),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_351),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_249),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_351),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_186),
.B(n_20),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_333),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_265),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_279),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_333),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_333),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_333),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_352),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_187),
.B(n_22),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_281),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_249),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_290),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_288),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_249),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_194),
.B(n_22),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_197),
.B(n_25),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_235),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_352),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_320),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_320),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_200),
.B(n_25),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_292),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_293),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_320),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_320),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_294),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_368),
.Y(n_462)
);

AND2x2_ASAP7_75t_SL g463 ( 
.A(n_369),
.B(n_205),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_419),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_419),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_376),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_419),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_378),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_424),
.B(n_416),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_367),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_422),
.Y(n_471)
);

BUFx10_ASAP7_75t_L g472 ( 
.A(n_461),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_383),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_371),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_395),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_422),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_422),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_371),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_372),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_417),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_425),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_327),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_372),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_426),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_431),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_374),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_453),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_416),
.B(n_235),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_399),
.B(n_225),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_438),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_407),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_394),
.B(n_397),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_437),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_437),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_447),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_447),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_374),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_380),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_370),
.B(n_345),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_423),
.B(n_235),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_385),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_410),
.B(n_229),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_386),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_437),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_388),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_387),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_388),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_393),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_390),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_393),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_407),
.B(n_263),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_398),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_398),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_379),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_401),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_423),
.B(n_354),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_391),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_392),
.Y(n_518)
);

AND2x6_ASAP7_75t_L g519 ( 
.A(n_401),
.B(n_205),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_408),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_408),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_409),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_400),
.B(n_263),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_409),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_402),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_418),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_418),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_404),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_R g529 ( 
.A(n_405),
.B(n_290),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_421),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_406),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_421),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_411),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_412),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_413),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_428),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_430),
.B(n_432),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_428),
.Y(n_538)
);

CKINVDCx16_ASAP7_75t_R g539 ( 
.A(n_381),
.Y(n_539)
);

OAI22x1_ASAP7_75t_L g540 ( 
.A1(n_499),
.A2(n_452),
.B1(n_373),
.B2(n_199),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_499),
.B(n_433),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_477),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_464),
.Y(n_543)
);

AND2x6_ASAP7_75t_L g544 ( 
.A(n_488),
.B(n_232),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_505),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_537),
.B(n_375),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_489),
.B(n_382),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_537),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_529),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_469),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_463),
.B(n_537),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_495),
.Y(n_552)
);

AND2x2_ASAP7_75t_SL g553 ( 
.A(n_463),
.B(n_451),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_L g554 ( 
.A(n_505),
.B(n_298),
.Y(n_554)
);

BUFx4f_ASAP7_75t_L g555 ( 
.A(n_463),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_537),
.B(n_434),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_501),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_505),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_505),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_512),
.B(n_414),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_469),
.B(n_429),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_512),
.B(n_415),
.Y(n_562)
);

BUFx10_ASAP7_75t_L g563 ( 
.A(n_498),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_492),
.B(n_427),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_501),
.B(n_439),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_488),
.B(n_429),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_523),
.B(n_445),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_505),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_534),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_501),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_474),
.B(n_478),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_496),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_505),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_464),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_474),
.Y(n_575)
);

AO21x2_ASAP7_75t_L g576 ( 
.A1(n_508),
.A2(n_530),
.B(n_479),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_500),
.B(n_435),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_478),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_477),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_472),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_479),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_500),
.B(n_443),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_512),
.B(n_448),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_483),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_464),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_491),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_483),
.B(n_457),
.Y(n_587)
);

OAI22xp33_ASAP7_75t_SL g588 ( 
.A1(n_482),
.A2(n_451),
.B1(n_389),
.B2(n_396),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_472),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_511),
.B(n_458),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_486),
.B(n_440),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_465),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_486),
.B(n_440),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_512),
.B(n_231),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_497),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_472),
.B(n_237),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_521),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_521),
.Y(n_598)
);

NOR2x1p5_ASAP7_75t_L g599 ( 
.A(n_503),
.B(n_297),
.Y(n_599)
);

BUFx6f_ASAP7_75t_SL g600 ( 
.A(n_472),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_507),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_510),
.B(n_238),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_510),
.B(n_441),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_465),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_513),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_465),
.B(n_232),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_482),
.A2(n_444),
.B1(n_450),
.B2(n_436),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_521),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_539),
.B(n_349),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_470),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_475),
.Y(n_611)
);

BUFx10_ASAP7_75t_L g612 ( 
.A(n_506),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_513),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_515),
.B(n_520),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_467),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_515),
.B(n_259),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_520),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_522),
.B(n_441),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_467),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_522),
.B(n_442),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_516),
.B(n_375),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_487),
.B(n_456),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_467),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_524),
.Y(n_624)
);

AND2x2_ASAP7_75t_SL g625 ( 
.A(n_533),
.B(n_369),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_533),
.Y(n_626)
);

BUFx8_ASAP7_75t_SL g627 ( 
.A(n_514),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_480),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_516),
.B(n_420),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_524),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_532),
.B(n_442),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_485),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_532),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_536),
.B(n_377),
.Y(n_634)
);

OAI22xp33_ASAP7_75t_L g635 ( 
.A1(n_509),
.A2(n_247),
.B1(n_303),
.B2(n_201),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_502),
.B(n_384),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_539),
.B(n_211),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_521),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_536),
.B(n_384),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_517),
.A2(n_353),
.B1(n_324),
.B2(n_377),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_538),
.B(n_446),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_494),
.Y(n_642)
);

INVx5_ASAP7_75t_L g643 ( 
.A(n_519),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_521),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_518),
.Y(n_645)
);

BUFx4f_ASAP7_75t_L g646 ( 
.A(n_519),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_SL g647 ( 
.A(n_525),
.B(n_324),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_538),
.B(n_446),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_508),
.B(n_449),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_473),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_528),
.B(n_261),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_514),
.B(n_420),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_530),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_521),
.B(n_271),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_531),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_535),
.B(n_219),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_494),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_468),
.B(n_403),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_471),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_494),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_526),
.B(n_527),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_504),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_SL g663 ( 
.A(n_462),
.B(n_353),
.Y(n_663)
);

NAND2xp33_ASAP7_75t_SL g664 ( 
.A(n_466),
.B(n_201),
.Y(n_664)
);

OR2x2_ASAP7_75t_SL g665 ( 
.A(n_481),
.B(n_227),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_477),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_504),
.B(n_403),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_504),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_519),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_471),
.B(n_449),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_476),
.B(n_454),
.Y(n_671)
);

INVx4_ASAP7_75t_SL g672 ( 
.A(n_519),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_476),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_526),
.B(n_273),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_519),
.A2(n_354),
.B1(n_267),
.B2(n_258),
.Y(n_675)
);

OAI21xp33_ASAP7_75t_SL g676 ( 
.A1(n_519),
.A2(n_256),
.B(n_222),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_484),
.B(n_266),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_526),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_477),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_526),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_526),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_519),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_527),
.B(n_460),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_527),
.B(n_283),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_527),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_552),
.B(n_490),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_575),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_543),
.Y(n_688)
);

NOR2x1p5_ASAP7_75t_L g689 ( 
.A(n_549),
.B(n_300),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_L g690 ( 
.A(n_580),
.B(n_527),
.Y(n_690)
);

NAND2xp33_ASAP7_75t_L g691 ( 
.A(n_580),
.B(n_477),
.Y(n_691)
);

NOR3xp33_ASAP7_75t_L g692 ( 
.A(n_626),
.B(n_275),
.C(n_268),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_636),
.B(n_493),
.Y(n_693)
);

NOR3xp33_ASAP7_75t_L g694 ( 
.A(n_626),
.B(n_569),
.C(n_645),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_639),
.B(n_493),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_574),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_547),
.B(n_493),
.Y(n_697)
);

NOR3xp33_ASAP7_75t_L g698 ( 
.A(n_645),
.B(n_306),
.C(n_291),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_553),
.A2(n_303),
.B1(n_247),
.B2(n_227),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_555),
.B(n_493),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_574),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_578),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_546),
.B(n_493),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_L g704 ( 
.A1(n_555),
.A2(n_331),
.B1(n_319),
.B2(n_326),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_546),
.B(n_493),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_555),
.B(n_185),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_564),
.B(n_307),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_563),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_546),
.B(n_192),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_581),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_553),
.B(n_202),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_544),
.B(n_224),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_584),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_587),
.B(n_309),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_585),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_595),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_625),
.A2(n_244),
.B1(n_289),
.B2(n_287),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_627),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_544),
.B(n_282),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_541),
.B(n_334),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_625),
.A2(n_289),
.B1(n_287),
.B2(n_347),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_544),
.B(n_321),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_610),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_572),
.B(n_357),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_548),
.B(n_198),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_589),
.B(n_360),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_589),
.B(n_198),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_550),
.B(n_312),
.Y(n_728)
);

INVx8_ASAP7_75t_L g729 ( 
.A(n_600),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_551),
.B(n_204),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_646),
.B(n_204),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_592),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_646),
.B(n_206),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_576),
.A2(n_550),
.B1(n_607),
.B2(n_605),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_592),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_566),
.B(n_206),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_622),
.A2(n_347),
.B1(n_350),
.B2(n_301),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_566),
.B(n_350),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_629),
.B(n_621),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_604),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_557),
.B(n_299),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_565),
.B(n_313),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_557),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_629),
.B(n_314),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_621),
.B(n_317),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_588),
.B(n_302),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_563),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_560),
.B(n_337),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_621),
.B(n_340),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_601),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_561),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_651),
.B(n_343),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_563),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_561),
.B(n_358),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_556),
.B(n_362),
.Y(n_755)
);

INVx8_ASAP7_75t_L g756 ( 
.A(n_600),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_542),
.B(n_304),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_576),
.A2(n_363),
.B1(n_366),
.B2(n_208),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_542),
.B(n_310),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_604),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_667),
.B(n_577),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_577),
.B(n_348),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_582),
.B(n_348),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_582),
.B(n_348),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_613),
.B(n_359),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_617),
.B(n_359),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_624),
.B(n_359),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_541),
.B(n_454),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_542),
.B(n_311),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_630),
.B(n_359),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_560),
.B(n_315),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_633),
.B(n_188),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_596),
.A2(n_316),
.B1(n_318),
.B2(n_322),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_562),
.B(n_189),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_562),
.B(n_583),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_655),
.B(n_609),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_671),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_671),
.Y(n_778)
);

OAI22x1_ASAP7_75t_L g779 ( 
.A1(n_640),
.A2(n_234),
.B1(n_236),
.B2(n_252),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_609),
.B(n_455),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_661),
.A2(n_614),
.B(n_571),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_641),
.Y(n_782)
);

INVx6_ASAP7_75t_L g783 ( 
.A(n_612),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_647),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_596),
.A2(n_325),
.B1(n_329),
.B2(n_335),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_542),
.B(n_336),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_655),
.B(n_208),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_579),
.B(n_341),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_576),
.A2(n_355),
.B1(n_361),
.B2(n_234),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_656),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_583),
.B(n_190),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_615),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_579),
.B(n_666),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_675),
.A2(n_361),
.B1(n_355),
.B2(n_252),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_634),
.B(n_191),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_SL g796 ( 
.A(n_549),
.B(n_193),
.Y(n_796)
);

AOI221xp5_ASAP7_75t_L g797 ( 
.A1(n_635),
.A2(n_342),
.B1(n_459),
.B2(n_455),
.C(n_460),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_567),
.B(n_212),
.Y(n_798)
);

BUFx5_ASAP7_75t_L g799 ( 
.A(n_573),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_579),
.B(n_298),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_591),
.A2(n_236),
.B(n_365),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_570),
.B(n_215),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_615),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_652),
.B(n_217),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_590),
.B(n_26),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_652),
.B(n_230),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_658),
.B(n_28),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_612),
.B(n_459),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_648),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_658),
.A2(n_594),
.B1(n_669),
.B2(n_682),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_656),
.B(n_28),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_545),
.B(n_31),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_579),
.B(n_298),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_R g814 ( 
.A(n_612),
.B(n_239),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_683),
.Y(n_815)
);

OR2x6_ASAP7_75t_L g816 ( 
.A(n_586),
.B(n_246),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_653),
.B(n_240),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_619),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_683),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_627),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_637),
.B(n_32),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_666),
.B(n_679),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_666),
.B(n_298),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_649),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_611),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_661),
.A2(n_356),
.B(n_241),
.Y(n_826)
);

NAND3xp33_ASAP7_75t_L g827 ( 
.A(n_663),
.B(n_285),
.C(n_339),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_602),
.B(n_616),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_637),
.B(n_35),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_666),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_619),
.A2(n_346),
.B1(n_246),
.B2(n_298),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_602),
.B(n_280),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_650),
.B(n_35),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_659),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_673),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_628),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_616),
.B(n_295),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_670),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_623),
.B(n_278),
.Y(n_839)
);

NAND3xp33_ASAP7_75t_L g840 ( 
.A(n_677),
.B(n_276),
.C(n_338),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_623),
.Y(n_841)
);

NAND2x1_ASAP7_75t_L g842 ( 
.A(n_545),
.B(n_346),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_642),
.A2(n_346),
.B1(n_246),
.B2(n_298),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_632),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_642),
.B(n_296),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_693),
.A2(n_618),
.B(n_631),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_758),
.A2(n_664),
.B1(n_540),
.B2(n_668),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_686),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_776),
.B(n_677),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_695),
.A2(n_603),
.B(n_620),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_697),
.A2(n_593),
.B(n_685),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_688),
.Y(n_852)
);

BUFx4f_ASAP7_75t_L g853 ( 
.A(n_783),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_707),
.B(n_657),
.Y(n_854)
);

AOI21x1_ASAP7_75t_L g855 ( 
.A1(n_700),
.A2(n_822),
.B(n_793),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_729),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_687),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_775),
.B(n_545),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_830),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_723),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_793),
.A2(n_644),
.B(n_597),
.Y(n_861)
);

AOI21x1_ASAP7_75t_L g862 ( 
.A1(n_700),
.A2(n_594),
.B(n_660),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_SL g863 ( 
.A(n_718),
.B(n_664),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_825),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_702),
.Y(n_865)
);

AO32x1_ASAP7_75t_L g866 ( 
.A1(n_710),
.A2(n_662),
.A3(n_668),
.B1(n_657),
.B2(n_660),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_SL g867 ( 
.A(n_820),
.B(n_669),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_R g868 ( 
.A(n_783),
.B(n_682),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_696),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_690),
.A2(n_608),
.B(n_681),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_713),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_691),
.A2(n_644),
.B(n_681),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_707),
.B(n_678),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_731),
.A2(n_678),
.B(n_558),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_805),
.A2(n_599),
.B1(n_684),
.B2(n_674),
.Y(n_875)
);

AO22x1_ASAP7_75t_L g876 ( 
.A1(n_805),
.A2(n_540),
.B1(n_665),
.B2(n_606),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_830),
.Y(n_877)
);

CKINVDCx10_ASAP7_75t_R g878 ( 
.A(n_816),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_731),
.A2(n_678),
.B(n_559),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_714),
.B(n_558),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_716),
.Y(n_881)
);

BUFx4f_ASAP7_75t_L g882 ( 
.A(n_783),
.Y(n_882)
);

AOI221xp5_ASAP7_75t_L g883 ( 
.A1(n_699),
.A2(n_676),
.B1(n_654),
.B2(n_665),
.C(n_554),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_771),
.A2(n_559),
.B(n_558),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_758),
.A2(n_606),
.B1(n_680),
.B2(n_598),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_SL g886 ( 
.A(n_836),
.B(n_643),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_811),
.A2(n_559),
.B1(n_568),
.B2(n_680),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_775),
.B(n_568),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_790),
.B(n_568),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_739),
.B(n_638),
.Y(n_890)
);

AO21x1_ASAP7_75t_L g891 ( 
.A1(n_771),
.A2(n_554),
.B(n_606),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_714),
.B(n_638),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_742),
.B(n_761),
.Y(n_893)
);

NOR2xp67_ASAP7_75t_L g894 ( 
.A(n_844),
.B(n_643),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_751),
.B(n_679),
.Y(n_895)
);

NOR2x1p5_ASAP7_75t_L g896 ( 
.A(n_708),
.B(n_305),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_784),
.B(n_679),
.Y(n_897)
);

OAI21x1_ASAP7_75t_L g898 ( 
.A1(n_800),
.A2(n_679),
.B(n_672),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_750),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_703),
.A2(n_606),
.B(n_643),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_705),
.A2(n_606),
.B(n_643),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_733),
.A2(n_643),
.B(n_243),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_708),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_811),
.A2(n_308),
.B(n_250),
.C(n_260),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_742),
.B(n_606),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_706),
.A2(n_330),
.B(n_323),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_726),
.B(n_672),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_746),
.A2(n_37),
.B(n_38),
.C(n_42),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_706),
.A2(n_274),
.B(n_262),
.Y(n_909)
);

INVx5_ASAP7_75t_L g910 ( 
.A(n_830),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_743),
.A2(n_346),
.B(n_246),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_746),
.A2(n_45),
.B(n_46),
.C(n_48),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_701),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_726),
.B(n_672),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_782),
.B(n_672),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_830),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_715),
.Y(n_917)
);

INVx11_ASAP7_75t_L g918 ( 
.A(n_747),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_747),
.B(n_46),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_813),
.A2(n_298),
.B(n_92),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_834),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_743),
.A2(n_88),
.B(n_165),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_752),
.B(n_49),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_816),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_734),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_809),
.B(n_51),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_802),
.A2(n_118),
.B(n_158),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_816),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_729),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_807),
.A2(n_55),
.B(n_57),
.C(n_58),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_711),
.B(n_55),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_796),
.B(n_57),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_835),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_734),
.A2(n_60),
.B1(n_62),
.B2(n_65),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_721),
.B(n_66),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_741),
.A2(n_68),
.B(n_74),
.Y(n_936)
);

AOI21x1_ASAP7_75t_L g937 ( 
.A1(n_813),
.A2(n_77),
.B(n_79),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_732),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_753),
.B(n_82),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_807),
.B(n_109),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_741),
.A2(n_119),
.B(n_128),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_774),
.A2(n_129),
.B(n_132),
.Y(n_942)
);

BUFx8_ASAP7_75t_L g943 ( 
.A(n_753),
.Y(n_943)
);

INVx4_ASAP7_75t_L g944 ( 
.A(n_729),
.Y(n_944)
);

NOR2x1_ASAP7_75t_L g945 ( 
.A(n_689),
.B(n_134),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_724),
.B(n_139),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_823),
.A2(n_730),
.B(n_824),
.Y(n_947)
);

AOI21x1_ASAP7_75t_L g948 ( 
.A1(n_765),
.A2(n_142),
.B(n_144),
.Y(n_948)
);

OAI22xp33_ASAP7_75t_L g949 ( 
.A1(n_717),
.A2(n_155),
.B1(n_157),
.B2(n_172),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_791),
.A2(n_772),
.B(n_795),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_756),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_828),
.A2(n_819),
.B(n_815),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_748),
.A2(n_812),
.B(n_728),
.C(n_737),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_799),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_777),
.Y(n_955)
);

AOI22x1_ASAP7_75t_L g956 ( 
.A1(n_801),
.A2(n_826),
.B1(n_838),
.B2(n_841),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_798),
.B(n_748),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_812),
.A2(n_728),
.B(n_810),
.C(n_773),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_727),
.A2(n_845),
.B(n_839),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_766),
.A2(n_767),
.B(n_770),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_727),
.A2(n_763),
.B(n_762),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_799),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_789),
.A2(n_778),
.B1(n_779),
.B2(n_794),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_709),
.B(n_804),
.Y(n_964)
);

AND2x2_ASAP7_75t_SL g965 ( 
.A(n_789),
.B(n_794),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_736),
.B(n_738),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_768),
.B(n_720),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_735),
.A2(n_803),
.B(n_760),
.Y(n_968)
);

O2A1O1Ixp5_ASAP7_75t_L g969 ( 
.A1(n_757),
.A2(n_788),
.B(n_786),
.C(n_769),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_806),
.B(n_754),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_740),
.A2(n_818),
.B(n_792),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_764),
.A2(n_725),
.B(n_817),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_808),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_744),
.A2(n_749),
.B(n_745),
.Y(n_974)
);

NOR3xp33_ASAP7_75t_L g975 ( 
.A(n_704),
.B(n_694),
.C(n_840),
.Y(n_975)
);

BUFx12f_ASAP7_75t_L g976 ( 
.A(n_787),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_712),
.A2(n_719),
.B(n_722),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_755),
.A2(n_842),
.B(n_837),
.Y(n_978)
);

NOR3xp33_ASAP7_75t_L g979 ( 
.A(n_698),
.B(n_692),
.C(n_829),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_821),
.A2(n_832),
.B(n_759),
.C(n_786),
.Y(n_980)
);

O2A1O1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_759),
.A2(n_788),
.B(n_833),
.C(n_780),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_787),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_827),
.A2(n_843),
.B(n_831),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_785),
.A2(n_831),
.B(n_843),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_814),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_799),
.Y(n_986)
);

OAI321xp33_ASAP7_75t_L g987 ( 
.A1(n_797),
.A2(n_805),
.A3(n_635),
.B1(n_811),
.B2(n_607),
.C(n_373),
.Y(n_987)
);

AOI221xp5_ASAP7_75t_L g988 ( 
.A1(n_814),
.A2(n_635),
.B1(n_588),
.B2(n_699),
.C(n_811),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_756),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_688),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_805),
.A2(n_761),
.B(n_588),
.C(n_746),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_SL g992 ( 
.A1(n_699),
.A2(n_383),
.B1(n_395),
.B2(n_367),
.Y(n_992)
);

NOR2xp67_ASAP7_75t_L g993 ( 
.A(n_836),
.B(n_645),
.Y(n_993)
);

NAND3xp33_ASAP7_75t_L g994 ( 
.A(n_805),
.B(n_503),
.C(n_498),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_830),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_805),
.A2(n_707),
.B1(n_811),
.B2(n_775),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_707),
.B(n_636),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_805),
.A2(n_555),
.B1(n_553),
.B2(n_775),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_707),
.B(n_636),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_686),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_693),
.A2(n_695),
.B(n_781),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_707),
.B(n_636),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_729),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_790),
.B(n_610),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_805),
.B(n_626),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_693),
.A2(n_695),
.B(n_781),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_718),
.Y(n_1007)
);

NOR3xp33_ASAP7_75t_L g1008 ( 
.A(n_805),
.B(n_811),
.C(n_588),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_723),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_805),
.B(n_626),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_775),
.B(n_739),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_687),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_688),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_688),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_693),
.A2(n_695),
.B(n_697),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_707),
.B(n_636),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_707),
.B(n_636),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_707),
.B(n_636),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_693),
.A2(n_695),
.B(n_697),
.Y(n_1019)
);

OAI321xp33_ASAP7_75t_L g1020 ( 
.A1(n_805),
.A2(n_635),
.A3(n_811),
.B1(n_607),
.B2(n_373),
.C(n_699),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_775),
.B(n_739),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_910),
.Y(n_1022)
);

BUFx4f_ASAP7_75t_L g1023 ( 
.A(n_929),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_997),
.A2(n_1002),
.B(n_999),
.Y(n_1024)
);

AOI21x1_ASAP7_75t_SL g1025 ( 
.A1(n_1016),
.A2(n_1018),
.B(n_1017),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1011),
.B(n_1021),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_862),
.A2(n_855),
.B(n_898),
.Y(n_1027)
);

BUFx4f_ASAP7_75t_SL g1028 ( 
.A(n_943),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_1011),
.B(n_1021),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_SL g1030 ( 
.A1(n_940),
.A2(n_953),
.B(n_958),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_910),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_910),
.Y(n_1032)
);

AOI21xp33_ASAP7_75t_L g1033 ( 
.A1(n_996),
.A2(n_987),
.B(n_1020),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_856),
.B(n_944),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_SL g1035 ( 
.A1(n_998),
.A2(n_935),
.B(n_888),
.Y(n_1035)
);

O2A1O1Ixp5_ASAP7_75t_L g1036 ( 
.A1(n_957),
.A2(n_961),
.B(n_1015),
.C(n_1019),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_967),
.B(n_893),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_954),
.A2(n_986),
.B(n_962),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_1008),
.A2(n_923),
.B(n_991),
.C(n_935),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_1007),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_849),
.B(n_1004),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_970),
.B(n_966),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_1009),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_1008),
.A2(n_970),
.B1(n_965),
.B2(n_875),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_880),
.A2(n_950),
.B(n_1001),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_SL g1046 ( 
.A(n_985),
.B(n_860),
.Y(n_1046)
);

AOI21x1_ASAP7_75t_SL g1047 ( 
.A1(n_873),
.A2(n_905),
.B(n_892),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_SL g1048 ( 
.A(n_988),
.B(n_979),
.C(n_975),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_858),
.A2(n_888),
.B(n_974),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_857),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_964),
.B(n_973),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_964),
.B(n_931),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_865),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_858),
.A2(n_1006),
.B(n_854),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_962),
.A2(n_986),
.B(n_960),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_965),
.A2(n_847),
.B1(n_963),
.B2(n_925),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_853),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_931),
.B(n_979),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_923),
.A2(n_991),
.B(n_912),
.C(n_908),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_846),
.A2(n_850),
.B(n_972),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1005),
.B(n_1010),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_910),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_959),
.A2(n_884),
.B(n_851),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_994),
.A2(n_871),
.B1(n_1012),
.B2(n_881),
.Y(n_1064)
);

NAND2x1_ASAP7_75t_L g1065 ( 
.A(n_859),
.B(n_995),
.Y(n_1065)
);

CKINVDCx11_ASAP7_75t_R g1066 ( 
.A(n_903),
.Y(n_1066)
);

AOI21x1_ASAP7_75t_SL g1067 ( 
.A1(n_926),
.A2(n_919),
.B(n_915),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_848),
.B(n_1000),
.Y(n_1068)
);

AOI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_980),
.A2(n_981),
.B(n_890),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_861),
.A2(n_879),
.B(n_874),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_872),
.A2(n_870),
.B(n_978),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_SL g1072 ( 
.A1(n_984),
.A2(n_946),
.B(n_981),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_908),
.A2(n_912),
.B(n_930),
.C(n_980),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_SL g1074 ( 
.A1(n_952),
.A2(n_947),
.B(n_891),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_899),
.B(n_955),
.Y(n_1075)
);

AOI21x1_ASAP7_75t_L g1076 ( 
.A1(n_977),
.A2(n_983),
.B(n_948),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1009),
.B(n_864),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_956),
.A2(n_971),
.B(n_968),
.Y(n_1078)
);

OA22x2_ASAP7_75t_L g1079 ( 
.A1(n_992),
.A2(n_982),
.B1(n_933),
.B2(n_921),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_963),
.A2(n_887),
.B1(n_904),
.B2(n_895),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_937),
.A2(n_969),
.B(n_920),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_869),
.Y(n_1082)
);

AO21x2_ASAP7_75t_L g1083 ( 
.A1(n_900),
.A2(n_901),
.B(n_911),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_934),
.A2(n_942),
.A3(n_866),
.B(n_990),
.Y(n_1084)
);

AOI221xp5_ASAP7_75t_L g1085 ( 
.A1(n_876),
.A2(n_949),
.B1(n_847),
.B2(n_863),
.C(n_883),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_975),
.A2(n_932),
.B(n_941),
.C(n_936),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_922),
.A2(n_927),
.B(n_859),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_864),
.B(n_897),
.Y(n_1088)
);

AOI21xp33_ASAP7_75t_L g1089 ( 
.A1(n_907),
.A2(n_897),
.B(n_914),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_945),
.A2(n_919),
.B(n_939),
.C(n_993),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_853),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_882),
.B(n_867),
.Y(n_1092)
);

AOI21x1_ASAP7_75t_L g1093 ( 
.A1(n_902),
.A2(n_889),
.B(n_906),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_SL g1094 ( 
.A1(n_856),
.A2(n_944),
.B(n_1003),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_866),
.A2(n_949),
.B(n_995),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_866),
.A2(n_877),
.B(n_916),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_913),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_877),
.B(n_916),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_877),
.A2(n_916),
.B(n_909),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_882),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_877),
.A2(n_916),
.B(n_885),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_868),
.B(n_924),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_976),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_928),
.B(n_989),
.Y(n_1104)
);

AOI211x1_ASAP7_75t_L g1105 ( 
.A1(n_896),
.A2(n_918),
.B(n_943),
.C(n_878),
.Y(n_1105)
);

NAND2x1p5_ASAP7_75t_L g1106 ( 
.A(n_929),
.B(n_951),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_886),
.A2(n_938),
.B(n_1013),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_917),
.A2(n_1014),
.B(n_894),
.Y(n_1108)
);

BUFx4f_ASAP7_75t_L g1109 ( 
.A(n_929),
.Y(n_1109)
);

OAI22x1_ASAP7_75t_L g1110 ( 
.A1(n_1003),
.A2(n_868),
.B1(n_929),
.B2(n_951),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_951),
.A2(n_1017),
.B(n_1016),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_951),
.B(n_997),
.Y(n_1112)
);

CKINVDCx8_ASAP7_75t_R g1113 ( 
.A(n_878),
.Y(n_1113)
);

BUFx12f_ASAP7_75t_L g1114 ( 
.A(n_943),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_860),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_997),
.A2(n_1017),
.B(n_1016),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_862),
.A2(n_855),
.B(n_898),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_997),
.A2(n_1017),
.B(n_1016),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_997),
.B(n_999),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_862),
.A2(n_855),
.B(n_898),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_856),
.B(n_944),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_997),
.B(n_999),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_996),
.A2(n_647),
.B1(n_805),
.B2(n_663),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_849),
.B(n_967),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_997),
.B(n_999),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_849),
.B(n_967),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_997),
.B(n_999),
.Y(n_1127)
);

AOI21xp33_ASAP7_75t_L g1128 ( 
.A1(n_996),
.A2(n_496),
.B(n_495),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_965),
.A2(n_1008),
.B1(n_988),
.B2(n_996),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_997),
.A2(n_1017),
.B(n_1016),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_862),
.A2(n_855),
.B(n_898),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_SL g1132 ( 
.A1(n_940),
.A2(n_953),
.B(n_958),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_862),
.A2(n_855),
.B(n_898),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_997),
.B(n_999),
.Y(n_1134)
);

INVxp67_ASAP7_75t_L g1135 ( 
.A(n_1009),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_857),
.Y(n_1136)
);

O2A1O1Ixp5_ASAP7_75t_L g1137 ( 
.A1(n_953),
.A2(n_805),
.B(n_998),
.C(n_958),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_997),
.A2(n_1017),
.B(n_1016),
.Y(n_1138)
);

AOI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1015),
.A2(n_1019),
.B(n_961),
.Y(n_1139)
);

O2A1O1Ixp5_ASAP7_75t_L g1140 ( 
.A1(n_953),
.A2(n_805),
.B(n_998),
.C(n_958),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_996),
.A2(n_647),
.B1(n_805),
.B2(n_663),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_997),
.B(n_999),
.Y(n_1142)
);

BUFx8_ASAP7_75t_SL g1143 ( 
.A(n_1007),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_849),
.B(n_967),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_997),
.A2(n_1017),
.B(n_1016),
.Y(n_1145)
);

AOI211x1_ASAP7_75t_L g1146 ( 
.A1(n_997),
.A2(n_999),
.B(n_1002),
.C(n_1016),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_1009),
.Y(n_1147)
);

INVx1_ASAP7_75t_SL g1148 ( 
.A(n_860),
.Y(n_1148)
);

AO31x2_ASAP7_75t_L g1149 ( 
.A1(n_891),
.A2(n_1015),
.A3(n_1019),
.B(n_998),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_997),
.A2(n_1017),
.B(n_1016),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_997),
.B(n_999),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_910),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_849),
.B(n_967),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_996),
.A2(n_997),
.B(n_1002),
.C(n_999),
.Y(n_1154)
);

AOI221xp5_ASAP7_75t_SL g1155 ( 
.A1(n_953),
.A2(n_811),
.B1(n_588),
.B2(n_999),
.C(n_997),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_910),
.Y(n_1156)
);

AOI221xp5_ASAP7_75t_SL g1157 ( 
.A1(n_953),
.A2(n_811),
.B1(n_588),
.B2(n_999),
.C(n_997),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_862),
.A2(n_855),
.B(n_898),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_997),
.B(n_999),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_SL g1160 ( 
.A1(n_996),
.A2(n_952),
.B(n_947),
.Y(n_1160)
);

AO21x1_ASAP7_75t_L g1161 ( 
.A1(n_996),
.A2(n_998),
.B(n_1008),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_852),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_910),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_997),
.A2(n_1017),
.B(n_1016),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_849),
.B(n_610),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_997),
.A2(n_1017),
.B(n_1016),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_997),
.B(n_999),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_849),
.B(n_967),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_996),
.A2(n_997),
.B1(n_1002),
.B2(n_999),
.Y(n_1169)
);

AOI21x1_ASAP7_75t_SL g1170 ( 
.A1(n_997),
.A2(n_1002),
.B(n_999),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_997),
.A2(n_1017),
.B(n_1016),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_910),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1026),
.A2(n_1029),
.B1(n_1129),
.B2(n_1169),
.Y(n_1173)
);

BUFx10_ASAP7_75t_L g1174 ( 
.A(n_1040),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1030),
.A2(n_1132),
.B(n_1035),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1050),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1154),
.B(n_1042),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1154),
.B(n_1042),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1142),
.B(n_1118),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1049),
.A2(n_1060),
.B(n_1137),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1043),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1057),
.B(n_1091),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1124),
.B(n_1126),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1052),
.B(n_1123),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_SL g1185 ( 
.A1(n_1142),
.A2(n_1145),
.B(n_1171),
.C(n_1024),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1116),
.B(n_1130),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1138),
.B(n_1150),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1144),
.B(n_1153),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_1032),
.B(n_1062),
.Y(n_1189)
);

OR2x2_ASAP7_75t_SL g1190 ( 
.A(n_1048),
.B(n_1058),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1119),
.B(n_1122),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1129),
.A2(n_1039),
.B1(n_1141),
.B2(n_1044),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1164),
.B(n_1166),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_1066),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1039),
.A2(n_1033),
.B(n_1059),
.C(n_1085),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1057),
.B(n_1091),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1168),
.B(n_1077),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1100),
.Y(n_1198)
);

BUFx4_ASAP7_75t_SL g1199 ( 
.A(n_1100),
.Y(n_1199)
);

INVx3_ASAP7_75t_R g1200 ( 
.A(n_1103),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_1143),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1125),
.B(n_1127),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1053),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1136),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1134),
.B(n_1151),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1159),
.B(n_1167),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1056),
.B(n_1155),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1023),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1034),
.B(n_1121),
.Y(n_1209)
);

INVx4_ASAP7_75t_L g1210 ( 
.A(n_1023),
.Y(n_1210)
);

CKINVDCx11_ASAP7_75t_R g1211 ( 
.A(n_1113),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1034),
.B(n_1121),
.Y(n_1212)
);

INVx4_ASAP7_75t_L g1213 ( 
.A(n_1109),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1056),
.B(n_1157),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1079),
.A2(n_1128),
.B1(n_1161),
.B2(n_1165),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1135),
.B(n_1051),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1147),
.B(n_1068),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1109),
.Y(n_1218)
);

OR2x6_ASAP7_75t_L g1219 ( 
.A(n_1105),
.B(n_1102),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1059),
.A2(n_1073),
.B1(n_1072),
.B2(n_1146),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_1028),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1068),
.B(n_1104),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1137),
.A2(n_1140),
.B(n_1054),
.Y(n_1223)
);

OR2x6_ASAP7_75t_L g1224 ( 
.A(n_1110),
.B(n_1114),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1111),
.B(n_1112),
.Y(n_1225)
);

INVx3_ASAP7_75t_SL g1226 ( 
.A(n_1115),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1140),
.A2(n_1045),
.B(n_1063),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_1143),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1088),
.B(n_1046),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1071),
.A2(n_1070),
.B(n_1036),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1148),
.B(n_1079),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1075),
.B(n_1066),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1114),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1036),
.A2(n_1086),
.B(n_1096),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1064),
.B(n_1097),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1160),
.B(n_1069),
.Y(n_1236)
);

BUFx10_ASAP7_75t_L g1237 ( 
.A(n_1032),
.Y(n_1237)
);

OR2x6_ASAP7_75t_L g1238 ( 
.A(n_1092),
.B(n_1101),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1022),
.B(n_1152),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1055),
.A2(n_1087),
.B(n_1073),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1080),
.A2(n_1090),
.B1(n_1061),
.B2(n_1089),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1032),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1162),
.B(n_1082),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1106),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1062),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1106),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1090),
.B(n_1028),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1062),
.Y(n_1248)
);

INVx4_ASAP7_75t_L g1249 ( 
.A(n_1062),
.Y(n_1249)
);

BUFx12f_ASAP7_75t_L g1250 ( 
.A(n_1163),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1163),
.Y(n_1251)
);

O2A1O1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1074),
.A2(n_1095),
.B(n_1098),
.C(n_1065),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1076),
.A2(n_1078),
.B(n_1139),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1163),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1022),
.B(n_1031),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1163),
.Y(n_1256)
);

O2A1O1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1094),
.A2(n_1099),
.B(n_1031),
.C(n_1156),
.Y(n_1257)
);

INVx4_ASAP7_75t_L g1258 ( 
.A(n_1172),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1172),
.A2(n_1156),
.B1(n_1107),
.B2(n_1067),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1172),
.B(n_1108),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_SL g1261 ( 
.A(n_1172),
.B(n_1067),
.Y(n_1261)
);

INVx4_ASAP7_75t_L g1262 ( 
.A(n_1083),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1038),
.B(n_1093),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1083),
.B(n_1120),
.Y(n_1264)
);

BUFx4_ASAP7_75t_SL g1265 ( 
.A(n_1025),
.Y(n_1265)
);

O2A1O1Ixp5_ASAP7_75t_SL g1266 ( 
.A1(n_1025),
.A2(n_1170),
.B(n_1047),
.C(n_1149),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1149),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1084),
.B(n_1081),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1027),
.A2(n_1117),
.B(n_1131),
.Y(n_1269)
);

O2A1O1Ixp5_ASAP7_75t_L g1270 ( 
.A1(n_1170),
.A2(n_1047),
.B(n_1084),
.C(n_1133),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1158),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1084),
.A2(n_1132),
.B(n_1030),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1124),
.B(n_1126),
.Y(n_1273)
);

INVx4_ASAP7_75t_L g1274 ( 
.A(n_1057),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1026),
.A2(n_996),
.B1(n_1029),
.B2(n_1129),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1026),
.B(n_1029),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1124),
.B(n_1126),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1057),
.Y(n_1278)
);

NOR2x1_ASAP7_75t_SL g1279 ( 
.A(n_1032),
.B(n_1062),
.Y(n_1279)
);

NAND3xp33_ASAP7_75t_L g1280 ( 
.A(n_1039),
.B(n_996),
.C(n_1008),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1057),
.Y(n_1281)
);

AO21x1_ASAP7_75t_L g1282 ( 
.A1(n_1044),
.A2(n_996),
.B(n_1033),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1124),
.B(n_1126),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1079),
.A2(n_992),
.B1(n_447),
.B2(n_383),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1026),
.B(n_1029),
.Y(n_1285)
);

NAND2x2_ASAP7_75t_L g1286 ( 
.A(n_1119),
.B(n_645),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1057),
.B(n_1091),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1030),
.A2(n_1132),
.B(n_1035),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1041),
.B(n_1037),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1057),
.B(n_1091),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1147),
.Y(n_1291)
);

NAND3xp33_ASAP7_75t_L g1292 ( 
.A(n_1039),
.B(n_996),
.C(n_1008),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1026),
.B(n_1029),
.Y(n_1293)
);

NAND2xp33_ASAP7_75t_L g1294 ( 
.A(n_1154),
.B(n_997),
.Y(n_1294)
);

INVx1_ASAP7_75t_SL g1295 ( 
.A(n_1115),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1026),
.A2(n_996),
.B1(n_1029),
.B2(n_1129),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1030),
.A2(n_1132),
.B(n_1035),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1043),
.Y(n_1298)
);

OR2x6_ASAP7_75t_SL g1299 ( 
.A(n_1040),
.B(n_718),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1057),
.B(n_1091),
.Y(n_1300)
);

INVx3_ASAP7_75t_L g1301 ( 
.A(n_1032),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1042),
.B(n_1142),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1147),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1023),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1032),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1043),
.Y(n_1306)
);

INVxp67_ASAP7_75t_L g1307 ( 
.A(n_1147),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1026),
.B(n_1029),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1057),
.B(n_1091),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1026),
.B(n_1029),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_SL g1311 ( 
.A(n_1113),
.B(n_569),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1026),
.B(n_1029),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1208),
.Y(n_1313)
);

BUFx2_ASAP7_75t_R g1314 ( 
.A(n_1299),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1192),
.B(n_1195),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1302),
.B(n_1191),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1211),
.Y(n_1317)
);

AO21x1_ASAP7_75t_L g1318 ( 
.A1(n_1192),
.A2(n_1220),
.B(n_1173),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1190),
.A2(n_1280),
.B1(n_1292),
.B2(n_1296),
.Y(n_1319)
);

OAI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1275),
.A2(n_1296),
.B1(n_1173),
.B2(n_1178),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1209),
.B(n_1212),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1237),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1231),
.A2(n_1275),
.B1(n_1220),
.B2(n_1207),
.Y(n_1323)
);

BUFx12f_ASAP7_75t_L g1324 ( 
.A(n_1233),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1250),
.Y(n_1325)
);

AOI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1269),
.A2(n_1288),
.B(n_1175),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1291),
.B(n_1303),
.Y(n_1327)
);

INVxp67_ASAP7_75t_L g1328 ( 
.A(n_1183),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1177),
.B(n_1178),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1177),
.B(n_1197),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1182),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1188),
.B(n_1273),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1203),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1254),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1284),
.A2(n_1282),
.B1(n_1184),
.B2(n_1215),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1207),
.A2(n_1214),
.B1(n_1247),
.B2(n_1229),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1204),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1217),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1227),
.A2(n_1234),
.B(n_1180),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1182),
.Y(n_1340)
);

CKINVDCx6p67_ASAP7_75t_R g1341 ( 
.A(n_1201),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1214),
.A2(n_1294),
.B1(n_1206),
.B2(n_1288),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1243),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1179),
.A2(n_1297),
.B1(n_1175),
.B2(n_1285),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1227),
.A2(n_1234),
.B(n_1180),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1239),
.B(n_1242),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1243),
.Y(n_1347)
);

AOI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1297),
.A2(n_1193),
.B(n_1187),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1179),
.A2(n_1312),
.B1(n_1293),
.B2(n_1285),
.Y(n_1349)
);

AND2x4_ASAP7_75t_SL g1350 ( 
.A(n_1210),
.B(n_1213),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1276),
.B(n_1293),
.Y(n_1351)
);

AOI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1186),
.A2(n_1193),
.B(n_1187),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1277),
.B(n_1283),
.Y(n_1353)
);

BUFx2_ASAP7_75t_R g1354 ( 
.A(n_1226),
.Y(n_1354)
);

INVx11_ASAP7_75t_L g1355 ( 
.A(n_1199),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1235),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1276),
.A2(n_1312),
.B1(n_1308),
.B2(n_1310),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1254),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1181),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1307),
.Y(n_1360)
);

OA21x2_ASAP7_75t_L g1361 ( 
.A1(n_1270),
.A2(n_1272),
.B(n_1223),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1272),
.A2(n_1232),
.B1(n_1224),
.B2(n_1216),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1225),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_SL g1364 ( 
.A1(n_1224),
.A2(n_1236),
.B1(n_1311),
.B2(n_1205),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1202),
.A2(n_1205),
.B1(n_1310),
.B2(n_1308),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1186),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1298),
.Y(n_1367)
);

BUFx10_ASAP7_75t_L g1368 ( 
.A(n_1208),
.Y(n_1368)
);

BUFx12f_ASAP7_75t_L g1369 ( 
.A(n_1174),
.Y(n_1369)
);

CKINVDCx14_ASAP7_75t_R g1370 ( 
.A(n_1228),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1222),
.B(n_1289),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_1200),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1306),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1268),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1202),
.B(n_1185),
.Y(n_1375)
);

AOI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1223),
.A2(n_1236),
.B(n_1259),
.Y(n_1376)
);

CKINVDCx11_ASAP7_75t_R g1377 ( 
.A(n_1174),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1255),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1218),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1241),
.A2(n_1224),
.B1(n_1267),
.B2(n_1219),
.Y(n_1380)
);

BUFx4_ASAP7_75t_R g1381 ( 
.A(n_1279),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1255),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1219),
.A2(n_1309),
.B1(n_1290),
.B2(n_1196),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1248),
.Y(n_1384)
);

AO21x1_ASAP7_75t_SL g1385 ( 
.A1(n_1265),
.A2(n_1261),
.B(n_1244),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1238),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1219),
.A2(n_1295),
.B1(n_1286),
.B2(n_1194),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1196),
.A2(n_1309),
.B1(n_1287),
.B2(n_1300),
.Y(n_1388)
);

OAI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1198),
.A2(n_1274),
.B1(n_1281),
.B2(n_1278),
.Y(n_1389)
);

BUFx2_ASAP7_75t_R g1390 ( 
.A(n_1256),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1254),
.Y(n_1391)
);

NAND2x1p5_ASAP7_75t_L g1392 ( 
.A(n_1249),
.B(n_1258),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1246),
.Y(n_1393)
);

BUFx10_ASAP7_75t_L g1394 ( 
.A(n_1218),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1287),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1237),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1242),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1266),
.A2(n_1259),
.B(n_1257),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_SL g1399 ( 
.A1(n_1260),
.A2(n_1300),
.B1(n_1290),
.B2(n_1274),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1262),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1245),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1245),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1249),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1251),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1301),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1221),
.B(n_1304),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1260),
.A2(n_1304),
.B1(n_1262),
.B2(n_1301),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1271),
.A2(n_1253),
.B(n_1252),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1253),
.Y(n_1409)
);

AO21x1_ASAP7_75t_L g1410 ( 
.A1(n_1252),
.A2(n_1264),
.B(n_1257),
.Y(n_1410)
);

NAND2x1p5_ASAP7_75t_L g1411 ( 
.A(n_1258),
.B(n_1305),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1305),
.Y(n_1412)
);

BUFx8_ASAP7_75t_L g1413 ( 
.A(n_1263),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1189),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1263),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1271),
.A2(n_1230),
.B(n_1227),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1176),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1302),
.A2(n_647),
.B1(n_1141),
.B2(n_1123),
.Y(n_1418)
);

INVx8_ASAP7_75t_L g1419 ( 
.A(n_1250),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1226),
.Y(n_1420)
);

INVxp33_ASAP7_75t_L g1421 ( 
.A(n_1229),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1209),
.B(n_1212),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1250),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1176),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_1211),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1230),
.A2(n_1227),
.B(n_1234),
.Y(n_1426)
);

INVx4_ASAP7_75t_L g1427 ( 
.A(n_1209),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1230),
.A2(n_1076),
.B(n_1240),
.Y(n_1428)
);

BUFx12f_ASAP7_75t_L g1429 ( 
.A(n_1211),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1428),
.A2(n_1326),
.B(n_1348),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1413),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1366),
.Y(n_1432)
);

AOI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1352),
.A2(n_1376),
.B(n_1375),
.Y(n_1433)
);

INVx3_ASAP7_75t_L g1434 ( 
.A(n_1413),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1385),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1374),
.B(n_1338),
.Y(n_1436)
);

INVx2_ASAP7_75t_SL g1437 ( 
.A(n_1413),
.Y(n_1437)
);

AO21x2_ASAP7_75t_L g1438 ( 
.A1(n_1398),
.A2(n_1320),
.B(n_1409),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1327),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1415),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1319),
.A2(n_1315),
.B(n_1320),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1365),
.B(n_1316),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1325),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1330),
.B(n_1329),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1363),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_SL g1446 ( 
.A1(n_1315),
.A2(n_1344),
.B1(n_1329),
.B2(n_1335),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1330),
.B(n_1356),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1408),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1335),
.A2(n_1318),
.B1(n_1323),
.B2(n_1418),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1365),
.B(n_1357),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1333),
.B(n_1337),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1343),
.Y(n_1452)
);

BUFx4f_ASAP7_75t_SL g1453 ( 
.A(n_1429),
.Y(n_1453)
);

INVxp67_ASAP7_75t_L g1454 ( 
.A(n_1332),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1347),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1386),
.B(n_1371),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1359),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1346),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1378),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1373),
.Y(n_1460)
);

INVx3_ASAP7_75t_L g1461 ( 
.A(n_1400),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1382),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1351),
.B(n_1349),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1400),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1361),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1361),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1417),
.B(n_1424),
.Y(n_1467)
);

AO21x1_ASAP7_75t_SL g1468 ( 
.A1(n_1342),
.A2(n_1380),
.B(n_1387),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1410),
.Y(n_1469)
);

INVx1_ASAP7_75t_SL g1470 ( 
.A(n_1354),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_1353),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1384),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1397),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1367),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1339),
.B(n_1345),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1361),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1339),
.B(n_1345),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_1355),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1331),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1325),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1342),
.B(n_1339),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1381),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1336),
.B(n_1328),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1360),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_SL g1485 ( 
.A(n_1314),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1345),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1426),
.B(n_1416),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1401),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1402),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1421),
.B(n_1389),
.Y(n_1490)
);

OAI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1421),
.A2(n_1389),
.B(n_1362),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1423),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1404),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1405),
.Y(n_1494)
);

OA21x2_ASAP7_75t_L g1495 ( 
.A1(n_1412),
.A2(n_1414),
.B(n_1393),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1391),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1334),
.B(n_1358),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1407),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1403),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1395),
.B(n_1331),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1358),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1358),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1383),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1411),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1340),
.B(n_1420),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1321),
.B(n_1422),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1381),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1427),
.B(n_1321),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1392),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1481),
.B(n_1387),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1481),
.B(n_1364),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1436),
.B(n_1438),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1444),
.B(n_1422),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1436),
.B(n_1388),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1448),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1495),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1438),
.B(n_1388),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1444),
.B(n_1422),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_1473),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1487),
.B(n_1438),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1487),
.B(n_1406),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1447),
.B(n_1486),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1448),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1447),
.B(n_1399),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1495),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1463),
.B(n_1396),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1439),
.B(n_1322),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1441),
.B(n_1469),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1475),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1431),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1465),
.B(n_1372),
.Y(n_1531)
);

AOI221xp5_ASAP7_75t_L g1532 ( 
.A1(n_1450),
.A2(n_1372),
.B1(n_1317),
.B2(n_1370),
.C(n_1350),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1466),
.B(n_1377),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1495),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1466),
.B(n_1377),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1477),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1469),
.B(n_1313),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1495),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1476),
.B(n_1341),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1476),
.B(n_1341),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1451),
.B(n_1390),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1451),
.B(n_1370),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1473),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1467),
.B(n_1369),
.Y(n_1544)
);

BUFx2_ASAP7_75t_R g1545 ( 
.A(n_1478),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1472),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1430),
.A2(n_1394),
.B(n_1368),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1459),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1459),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1467),
.B(n_1369),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1432),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1448),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1462),
.Y(n_1553)
);

AOI211xp5_ASAP7_75t_L g1554 ( 
.A1(n_1491),
.A2(n_1317),
.B(n_1379),
.C(n_1429),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1528),
.B(n_1546),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1545),
.B(n_1470),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1528),
.B(n_1457),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1545),
.B(n_1453),
.Y(n_1558)
);

NAND3xp33_ASAP7_75t_L g1559 ( 
.A(n_1526),
.B(n_1446),
.C(n_1490),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1546),
.B(n_1484),
.Y(n_1560)
);

NAND3xp33_ASAP7_75t_L g1561 ( 
.A(n_1526),
.B(n_1449),
.C(n_1442),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_R g1562 ( 
.A(n_1541),
.B(n_1425),
.Y(n_1562)
);

NAND3xp33_ASAP7_75t_L g1563 ( 
.A(n_1537),
.B(n_1520),
.C(n_1516),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1521),
.B(n_1440),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1554),
.A2(n_1485),
.B1(n_1482),
.B2(n_1483),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1554),
.B(n_1482),
.Y(n_1566)
);

NOR3xp33_ASAP7_75t_L g1567 ( 
.A(n_1532),
.B(n_1499),
.C(n_1433),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1522),
.B(n_1474),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1511),
.A2(n_1503),
.B1(n_1498),
.B2(n_1435),
.Y(n_1569)
);

NAND2xp33_ASAP7_75t_L g1570 ( 
.A(n_1541),
.B(n_1435),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1511),
.A2(n_1503),
.B1(n_1498),
.B2(n_1435),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1532),
.A2(n_1482),
.B1(n_1507),
.B2(n_1471),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1527),
.A2(n_1507),
.B1(n_1454),
.B2(n_1437),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1551),
.B(n_1519),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1551),
.B(n_1460),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1519),
.B(n_1499),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1519),
.B(n_1462),
.Y(n_1577)
);

AND2x2_ASAP7_75t_SL g1578 ( 
.A(n_1517),
.B(n_1506),
.Y(n_1578)
);

OAI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1537),
.A2(n_1501),
.B(n_1505),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1543),
.B(n_1445),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1543),
.B(n_1452),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1513),
.B(n_1518),
.Y(n_1582)
);

NAND2xp33_ASAP7_75t_R g1583 ( 
.A(n_1541),
.B(n_1478),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1518),
.B(n_1464),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1543),
.B(n_1452),
.Y(n_1585)
);

NAND3xp33_ASAP7_75t_L g1586 ( 
.A(n_1520),
.B(n_1455),
.C(n_1494),
.Y(n_1586)
);

NAND4xp25_ASAP7_75t_L g1587 ( 
.A(n_1542),
.B(n_1494),
.C(n_1493),
.D(n_1488),
.Y(n_1587)
);

AOI221xp5_ASAP7_75t_L g1588 ( 
.A1(n_1520),
.A2(n_1455),
.B1(n_1488),
.B2(n_1493),
.C(n_1496),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1542),
.B(n_1489),
.Y(n_1589)
);

NAND4xp25_ASAP7_75t_L g1590 ( 
.A(n_1542),
.B(n_1501),
.C(n_1480),
.D(n_1443),
.Y(n_1590)
);

OAI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1517),
.A2(n_1505),
.B1(n_1496),
.B2(n_1500),
.C(n_1489),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_SL g1592 ( 
.A1(n_1531),
.A2(n_1434),
.B(n_1508),
.Y(n_1592)
);

OAI21xp33_ASAP7_75t_L g1593 ( 
.A1(n_1510),
.A2(n_1433),
.B(n_1502),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1531),
.B(n_1456),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1533),
.B(n_1458),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1527),
.B(n_1479),
.Y(n_1596)
);

NOR3xp33_ASAP7_75t_L g1597 ( 
.A(n_1533),
.B(n_1509),
.C(n_1504),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1510),
.B(n_1461),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1539),
.B(n_1540),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1553),
.B(n_1497),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1553),
.B(n_1497),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_SL g1602 ( 
.A1(n_1533),
.A2(n_1434),
.B(n_1508),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1582),
.B(n_1515),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1574),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1555),
.B(n_1512),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1568),
.B(n_1512),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1575),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1586),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1588),
.B(n_1529),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1582),
.B(n_1515),
.Y(n_1610)
);

NAND2x1p5_ASAP7_75t_L g1611 ( 
.A(n_1566),
.B(n_1547),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1577),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1598),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1580),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1558),
.B(n_1324),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1581),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1585),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1562),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1560),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1561),
.A2(n_1468),
.B1(n_1517),
.B2(n_1524),
.Y(n_1620)
);

NOR2xp67_ASAP7_75t_L g1621 ( 
.A(n_1563),
.B(n_1516),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1598),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1599),
.B(n_1515),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1599),
.B(n_1523),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1557),
.B(n_1512),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1597),
.B(n_1535),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1600),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1601),
.Y(n_1628)
);

NAND2x1p5_ASAP7_75t_L g1629 ( 
.A(n_1566),
.B(n_1547),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1564),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1589),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1594),
.B(n_1536),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1576),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1579),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1593),
.B(n_1536),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1591),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1587),
.B(n_1514),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1608),
.B(n_1609),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1613),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1612),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1603),
.B(n_1584),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1621),
.B(n_1523),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1613),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1603),
.B(n_1610),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1632),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1608),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1621),
.B(n_1552),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1618),
.B(n_1544),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1609),
.B(n_1559),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1618),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1634),
.B(n_1548),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1612),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1613),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1634),
.B(n_1548),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1610),
.B(n_1552),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1622),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1632),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1614),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1614),
.B(n_1549),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1610),
.B(n_1567),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1611),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1616),
.Y(n_1662)
);

AOI211xp5_ASAP7_75t_L g1663 ( 
.A1(n_1637),
.A2(n_1565),
.B(n_1572),
.C(n_1570),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1623),
.B(n_1624),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1622),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1604),
.Y(n_1666)
);

NOR2x1_ASAP7_75t_L g1667 ( 
.A(n_1615),
.B(n_1570),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1616),
.B(n_1549),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1606),
.B(n_1596),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1617),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1666),
.B(n_1607),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1650),
.B(n_1630),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1646),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1659),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1666),
.B(n_1607),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1648),
.B(n_1556),
.Y(n_1676)
);

INVx2_ASAP7_75t_SL g1677 ( 
.A(n_1650),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_L g1678 ( 
.A(n_1667),
.B(n_1425),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1659),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1650),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1646),
.B(n_1637),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1668),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1667),
.Y(n_1683)
);

NAND2x1p5_ASAP7_75t_L g1684 ( 
.A(n_1642),
.B(n_1530),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1639),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1638),
.B(n_1669),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1668),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1638),
.B(n_1669),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1660),
.B(n_1630),
.Y(n_1689)
);

NAND4xp25_ASAP7_75t_L g1690 ( 
.A(n_1660),
.B(n_1540),
.C(n_1583),
.D(n_1619),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1651),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1651),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1638),
.B(n_1625),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1654),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1654),
.Y(n_1695)
);

OAI21xp5_ASAP7_75t_SL g1696 ( 
.A1(n_1660),
.A2(n_1629),
.B(n_1611),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1640),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1640),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1652),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1649),
.B(n_1619),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1652),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1649),
.B(n_1617),
.Y(n_1702)
);

O2A1O1Ixp33_ASAP7_75t_L g1703 ( 
.A1(n_1649),
.A2(n_1636),
.B(n_1611),
.C(n_1629),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1661),
.A2(n_1636),
.B1(n_1620),
.B2(n_1525),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1669),
.B(n_1606),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1648),
.B(n_1626),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1658),
.Y(n_1707)
);

NAND4xp25_ASAP7_75t_L g1708 ( 
.A(n_1663),
.B(n_1540),
.C(n_1535),
.D(n_1590),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1658),
.B(n_1604),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1639),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1645),
.B(n_1625),
.Y(n_1711)
);

AOI21xp33_ASAP7_75t_L g1712 ( 
.A1(n_1670),
.A2(n_1635),
.B(n_1629),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1645),
.B(n_1605),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1641),
.B(n_1623),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1697),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1678),
.B(n_1644),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1699),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1698),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1700),
.B(n_1662),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1701),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1707),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1673),
.B(n_1662),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1676),
.B(n_1324),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1689),
.B(n_1644),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1686),
.Y(n_1725)
);

NAND3x1_ASAP7_75t_L g1726 ( 
.A(n_1681),
.B(n_1550),
.C(n_1544),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1688),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1689),
.B(n_1644),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1671),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1675),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1704),
.A2(n_1661),
.B1(n_1645),
.B2(n_1657),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1702),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1680),
.B(n_1657),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1709),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1705),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1705),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1693),
.B(n_1657),
.Y(n_1737)
);

AND2x4_ASAP7_75t_SL g1738 ( 
.A(n_1676),
.B(n_1544),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1704),
.A2(n_1661),
.B1(n_1611),
.B2(n_1629),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1674),
.Y(n_1740)
);

INVx1_ASAP7_75t_SL g1741 ( 
.A(n_1672),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1679),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1706),
.B(n_1670),
.Y(n_1743)
);

NAND4xp75_ASAP7_75t_L g1744 ( 
.A(n_1683),
.B(n_1569),
.C(n_1571),
.D(n_1578),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1677),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1682),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1687),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1685),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1684),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1672),
.B(n_1664),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1724),
.B(n_1683),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1718),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1716),
.B(n_1677),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1741),
.B(n_1706),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1735),
.B(n_1695),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1718),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1736),
.B(n_1691),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1737),
.B(n_1692),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1738),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1750),
.Y(n_1760)
);

OAI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1731),
.A2(n_1703),
.B1(n_1696),
.B2(n_1661),
.C(n_1712),
.Y(n_1761)
);

NAND3xp33_ASAP7_75t_L g1762 ( 
.A(n_1745),
.B(n_1694),
.C(n_1663),
.Y(n_1762)
);

INVx1_ASAP7_75t_SL g1763 ( 
.A(n_1738),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1720),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1725),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1726),
.A2(n_1744),
.B1(n_1739),
.B2(n_1716),
.Y(n_1766)
);

AOI221x1_ASAP7_75t_L g1767 ( 
.A1(n_1715),
.A2(n_1717),
.B1(n_1730),
.B2(n_1729),
.C(n_1725),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1720),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1721),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_SL g1770 ( 
.A(n_1723),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1727),
.B(n_1732),
.Y(n_1771)
);

OAI21xp33_ASAP7_75t_L g1772 ( 
.A1(n_1743),
.A2(n_1708),
.B(n_1690),
.Y(n_1772)
);

INVxp67_ASAP7_75t_SL g1773 ( 
.A(n_1726),
.Y(n_1773)
);

AOI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1719),
.A2(n_1647),
.B(n_1642),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1727),
.Y(n_1775)
);

INVxp67_ASAP7_75t_L g1776 ( 
.A(n_1722),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1765),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1775),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1764),
.Y(n_1779)
);

CKINVDCx16_ASAP7_75t_R g1780 ( 
.A(n_1770),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1754),
.B(n_1734),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1771),
.B(n_1715),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1751),
.B(n_1724),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1764),
.Y(n_1784)
);

INVx1_ASAP7_75t_SL g1785 ( 
.A(n_1751),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1771),
.B(n_1740),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1759),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1752),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1766),
.A2(n_1748),
.B1(n_1737),
.B2(n_1685),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1760),
.B(n_1728),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1756),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1760),
.B(n_1728),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1768),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1776),
.B(n_1742),
.Y(n_1794)
);

NAND2x1p5_ASAP7_75t_L g1795 ( 
.A(n_1753),
.B(n_1443),
.Y(n_1795)
);

NAND2xp33_ASAP7_75t_L g1796 ( 
.A(n_1762),
.B(n_1733),
.Y(n_1796)
);

OAI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1796),
.A2(n_1767),
.B(n_1773),
.Y(n_1797)
);

AOI21xp33_ASAP7_75t_SL g1798 ( 
.A1(n_1780),
.A2(n_1753),
.B(n_1761),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1785),
.B(n_1790),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1796),
.A2(n_1767),
.B(n_1772),
.Y(n_1800)
);

NAND3xp33_ASAP7_75t_SL g1801 ( 
.A(n_1789),
.B(n_1763),
.C(n_1774),
.Y(n_1801)
);

OAI31xp33_ASAP7_75t_L g1802 ( 
.A1(n_1786),
.A2(n_1753),
.A3(n_1758),
.B(n_1769),
.Y(n_1802)
);

AOI221xp5_ASAP7_75t_L g1803 ( 
.A1(n_1782),
.A2(n_1757),
.B1(n_1755),
.B2(n_1747),
.C(n_1746),
.Y(n_1803)
);

AOI322xp5_ASAP7_75t_L g1804 ( 
.A1(n_1781),
.A2(n_1748),
.A3(n_1635),
.B1(n_1747),
.B2(n_1710),
.C1(n_1721),
.C2(n_1750),
.Y(n_1804)
);

OAI221xp5_ASAP7_75t_SL g1805 ( 
.A1(n_1783),
.A2(n_1777),
.B1(n_1792),
.B2(n_1790),
.C(n_1787),
.Y(n_1805)
);

OAI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1783),
.A2(n_1744),
.B1(n_1792),
.B2(n_1795),
.Y(n_1806)
);

OAI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1795),
.A2(n_1758),
.B1(n_1749),
.B2(n_1710),
.C(n_1684),
.Y(n_1807)
);

AOI222xp33_ASAP7_75t_L g1808 ( 
.A1(n_1777),
.A2(n_1749),
.B1(n_1538),
.B2(n_1534),
.C1(n_1525),
.C2(n_1642),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_SL g1809 ( 
.A(n_1800),
.B(n_1795),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1799),
.B(n_1778),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1797),
.B(n_1806),
.Y(n_1811)
);

INVx3_ASAP7_75t_L g1812 ( 
.A(n_1805),
.Y(n_1812)
);

NAND3xp33_ASAP7_75t_L g1813 ( 
.A(n_1802),
.B(n_1791),
.C(n_1788),
.Y(n_1813)
);

NOR2x1_ASAP7_75t_L g1814 ( 
.A(n_1801),
.B(n_1779),
.Y(n_1814)
);

NOR2x1_ASAP7_75t_L g1815 ( 
.A(n_1807),
.B(n_1784),
.Y(n_1815)
);

NAND3xp33_ASAP7_75t_SL g1816 ( 
.A(n_1798),
.B(n_1803),
.C(n_1804),
.Y(n_1816)
);

NOR2xp67_ASAP7_75t_SL g1817 ( 
.A(n_1808),
.B(n_1480),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1799),
.Y(n_1818)
);

NOR4xp25_ASAP7_75t_L g1819 ( 
.A(n_1797),
.B(n_1793),
.C(n_1794),
.D(n_1749),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1799),
.B(n_1711),
.Y(n_1820)
);

AOI321xp33_ASAP7_75t_L g1821 ( 
.A1(n_1819),
.A2(n_1811),
.A3(n_1814),
.B1(n_1809),
.B2(n_1815),
.C(n_1812),
.Y(n_1821)
);

NOR3xp33_ASAP7_75t_L g1822 ( 
.A(n_1816),
.B(n_1711),
.C(n_1713),
.Y(n_1822)
);

NOR4xp25_ASAP7_75t_L g1823 ( 
.A(n_1812),
.B(n_1713),
.C(n_1670),
.D(n_1643),
.Y(n_1823)
);

OAI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1813),
.A2(n_1647),
.B(n_1642),
.Y(n_1824)
);

OAI211xp5_ASAP7_75t_SL g1825 ( 
.A1(n_1810),
.A2(n_1592),
.B(n_1602),
.C(n_1643),
.Y(n_1825)
);

NOR3x1_ASAP7_75t_L g1826 ( 
.A(n_1820),
.B(n_1595),
.C(n_1573),
.Y(n_1826)
);

NOR2x1_ASAP7_75t_L g1827 ( 
.A(n_1821),
.B(n_1818),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1822),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1823),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1826),
.Y(n_1830)
);

AOI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1824),
.A2(n_1817),
.B1(n_1647),
.B2(n_1642),
.Y(n_1831)
);

NOR2x1_ASAP7_75t_L g1832 ( 
.A(n_1825),
.B(n_1492),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1821),
.B(n_1647),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1827),
.B(n_1714),
.Y(n_1834)
);

NAND3xp33_ASAP7_75t_L g1835 ( 
.A(n_1829),
.B(n_1492),
.C(n_1647),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1833),
.B(n_1639),
.Y(n_1836)
);

OR5x1_ASAP7_75t_L g1837 ( 
.A(n_1828),
.B(n_1714),
.C(n_1664),
.D(n_1633),
.E(n_1655),
.Y(n_1837)
);

NOR5xp2_ASAP7_75t_L g1838 ( 
.A(n_1830),
.B(n_1633),
.C(n_1628),
.D(n_1627),
.E(n_1631),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1832),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1834),
.Y(n_1840)
);

XNOR2x1_ASAP7_75t_L g1841 ( 
.A(n_1839),
.B(n_1831),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1836),
.Y(n_1842)
);

AOI22x1_ASAP7_75t_L g1843 ( 
.A1(n_1840),
.A2(n_1837),
.B1(n_1835),
.B2(n_1838),
.Y(n_1843)
);

O2A1O1Ixp33_ASAP7_75t_L g1844 ( 
.A1(n_1843),
.A2(n_1842),
.B(n_1841),
.C(n_1643),
.Y(n_1844)
);

OAI22x1_ASAP7_75t_L g1845 ( 
.A1(n_1844),
.A2(n_1656),
.B1(n_1639),
.B2(n_1665),
.Y(n_1845)
);

OAI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1844),
.A2(n_1653),
.B(n_1643),
.Y(n_1846)
);

OAI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1846),
.A2(n_1656),
.B(n_1653),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1845),
.B(n_1653),
.Y(n_1848)
);

AOI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1848),
.A2(n_1656),
.B(n_1653),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1847),
.A2(n_1665),
.B(n_1656),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1849),
.Y(n_1851)
);

AOI22xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1851),
.A2(n_1850),
.B1(n_1550),
.B2(n_1664),
.Y(n_1852)
);

AOI221xp5_ASAP7_75t_L g1853 ( 
.A1(n_1852),
.A2(n_1665),
.B1(n_1550),
.B2(n_1419),
.C(n_1350),
.Y(n_1853)
);

AOI211xp5_ASAP7_75t_L g1854 ( 
.A1(n_1853),
.A2(n_1535),
.B(n_1665),
.C(n_1379),
.Y(n_1854)
);


endmodule