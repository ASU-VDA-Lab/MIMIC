module fake_jpeg_12974_n_102 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_30),
.A2(n_16),
.B1(n_27),
.B2(n_24),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_47),
.B1(n_36),
.B2(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_59),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_2),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_38),
.C(n_31),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_63),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_40),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_41),
.B1(n_34),
.B2(n_18),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_65),
.B1(n_74),
.B2(n_75),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_41),
.B1(n_34),
.B2(n_3),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_1),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_72),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_29),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_8),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_3),
.B(n_4),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_6),
.Y(n_76)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_67),
.C(n_62),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_75),
.B1(n_73),
.B2(n_71),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_20),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_85),
.B(n_9),
.Y(n_92)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_83),
.Y(n_89)
);

INVxp67_ASAP7_75t_SL g94 ( 
.A(n_89),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_82),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_78),
.B(n_87),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_96),
.B(n_82),
.Y(n_97)
);

OAI221xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_85),
.B1(n_88),
.B2(n_79),
.C(n_81),
.Y(n_98)
);

AOI31xp67_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_92),
.A3(n_94),
.B(n_80),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_12),
.B(n_14),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_19),
.Y(n_101)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_101),
.Y(n_102)
);


endmodule