module real_jpeg_7577_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_0),
.A2(n_256),
.B1(n_259),
.B2(n_262),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_0),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_0),
.B(n_275),
.C(n_278),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_0),
.B(n_111),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_0),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_0),
.B(n_163),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_0),
.B(n_239),
.Y(n_348)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_1),
.Y(n_178)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_1),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_1),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_1),
.Y(n_284)
);

INVx8_ASAP7_75t_L g397 ( 
.A(n_1),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_1),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_1),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_2),
.A2(n_126),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_2),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_2),
.A2(n_131),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_2),
.A2(n_131),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_3),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g417 ( 
.A(n_3),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_4),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_5),
.A2(n_148),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_5),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_5),
.A2(n_85),
.B1(n_187),
.B2(n_242),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_5),
.A2(n_160),
.B1(n_242),
.B2(n_338),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g436 ( 
.A1(n_5),
.A2(n_242),
.B1(n_437),
.B2(n_438),
.Y(n_436)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_6),
.Y(n_410)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_7),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_8),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_8),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_8),
.A2(n_124),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_8),
.A2(n_124),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_8),
.A2(n_124),
.B1(n_315),
.B2(n_426),
.Y(n_425)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_9),
.Y(n_277)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_11),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_12),
.A2(n_51),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_12),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_12),
.A2(n_202),
.B1(n_265),
.B2(n_268),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_12),
.A2(n_202),
.B1(n_286),
.B2(n_290),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_12),
.A2(n_202),
.B1(n_351),
.B2(n_353),
.Y(n_350)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_13),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_14),
.A2(n_265),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_14),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_14),
.A2(n_298),
.B1(n_312),
.B2(n_316),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_14),
.A2(n_42),
.B1(n_298),
.B2(n_382),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_14),
.A2(n_33),
.B1(n_59),
.B2(n_298),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_15),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_15),
.A2(n_60),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_15),
.A2(n_60),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_15),
.A2(n_60),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_16),
.A2(n_49),
.B1(n_50),
.B2(n_53),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_16),
.A2(n_49),
.B1(n_234),
.B2(n_238),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_16),
.A2(n_49),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_16),
.A2(n_49),
.B1(n_443),
.B2(n_445),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_17),
.A2(n_66),
.B1(n_89),
.B2(n_93),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_17),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_17),
.A2(n_93),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_17),
.A2(n_93),
.B1(n_183),
.B2(n_187),
.Y(n_182)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_511),
.B(n_513),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_205),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_204),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_150),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_24),
.B(n_150),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_132),
.B2(n_133),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_61),
.C(n_94),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_27),
.A2(n_134),
.B1(n_135),
.B2(n_149),
.Y(n_133)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_27),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_27),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_47),
.B1(n_55),
.B2(n_57),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_28),
.A2(n_55),
.B1(n_57),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_28),
.A2(n_241),
.B(n_244),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_28),
.A2(n_55),
.B1(n_241),
.B2(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_29),
.B(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_29),
.A2(n_414),
.B(n_433),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_37),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_33),
.Y(n_203)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g126 ( 
.A(n_40),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_41),
.Y(n_123)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_41),
.Y(n_130)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_41),
.Y(n_172)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_46),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_48),
.B(n_56),
.Y(n_199)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI32xp33_ASAP7_75t_L g406 ( 
.A1(n_53),
.A2(n_407),
.A3(n_409),
.B1(n_411),
.B2(n_414),
.Y(n_406)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_55),
.B(n_262),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_55),
.A2(n_200),
.B(n_466),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_56),
.B(n_201),
.Y(n_244)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_58),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_61),
.A2(n_62),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_61),
.A2(n_62),
.B1(n_94),
.B2(n_95),
.Y(n_152)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_77),
.B(n_88),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_63),
.A2(n_255),
.B(n_263),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_63),
.A2(n_77),
.B1(n_296),
.B2(n_337),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_63),
.A2(n_263),
.B(n_337),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_63),
.A2(n_77),
.B1(n_442),
.B2(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_64),
.A2(n_156),
.B1(n_163),
.B2(n_164),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_64),
.A2(n_156),
.B1(n_163),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_64),
.A2(n_163),
.B1(n_193),
.B2(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_64),
.B(n_264),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_77),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B1(n_72),
.B2(n_74),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_68),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_68),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_68),
.Y(n_258)
);

INVx6_ASAP7_75t_L g446 ( 
.A(n_68),
.Y(n_446)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_69),
.Y(n_267)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_69),
.Y(n_340)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_75),
.Y(n_159)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_77),
.A2(n_296),
.B(n_299),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_77),
.A2(n_299),
.B(n_442),
.Y(n_441)
);

AOI22x1_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_85),
.B2(n_87),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_83),
.Y(n_179)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_83),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_84),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_84),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_85),
.B(n_306),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_86),
.Y(n_222)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_86),
.Y(n_394)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_92),
.Y(n_261)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_92),
.Y(n_366)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_120),
.B1(n_127),
.B2(n_128),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_96),
.A2(n_127),
.B1(n_128),
.B2(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_96),
.A2(n_127),
.B1(n_168),
.B2(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_96),
.A2(n_127),
.B1(n_381),
.B2(n_436),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_111),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_103),
.B1(n_106),
.B2(n_109),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_102),
.Y(n_368)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_105),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g352 ( 
.A(n_105),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_105),
.Y(n_355)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_105),
.Y(n_413)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g383 ( 
.A(n_110),
.Y(n_383)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_110),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_111),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_111),
.A2(n_121),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_111),
.A2(n_166),
.B1(n_385),
.B2(n_468),
.Y(n_467)
);

AO22x2_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_114),
.Y(n_230)
);

INVx5_ASAP7_75t_L g444 ( 
.A(n_114),
.Y(n_444)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_115),
.Y(n_197)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_118),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_123),
.Y(n_346)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_123),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_127),
.B(n_350),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_127),
.A2(n_381),
.B(n_384),
.Y(n_380)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_130),
.Y(n_239)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_143),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.C(n_173),
.Y(n_150)
);

FAx1_ASAP7_75t_SL g207 ( 
.A(n_151),
.B(n_154),
.CI(n_173),
.CON(n_207),
.SN(n_207)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_154),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_165),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_155),
.Y(n_216)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_159),
.Y(n_273)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp33_ASAP7_75t_SL g369 ( 
.A(n_161),
.B(n_370),
.Y(n_369)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_162),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_163),
.B(n_264),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_166),
.A2(n_343),
.B(n_349),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_166),
.B(n_385),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_166),
.A2(n_349),
.B(n_484),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B(n_198),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_192),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_175),
.A2(n_198),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_175),
.A2(n_192),
.B1(n_213),
.B2(n_455),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_180),
.B(n_182),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_176),
.A2(n_182),
.B1(n_220),
.B2(n_225),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_176),
.A2(n_281),
.B(n_282),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_176),
.A2(n_262),
.B(n_282),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_176),
.A2(n_420),
.B1(n_421),
.B2(n_424),
.Y(n_419)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_177),
.B(n_285),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_177),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_177),
.A2(n_359),
.B1(n_389),
.B2(n_395),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_177),
.A2(n_425),
.B1(n_461),
.B2(n_462),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_179),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_180),
.A2(n_311),
.B(n_319),
.Y(n_310)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_181),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_185),
.Y(n_292)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

BUFx8_ASAP7_75t_L g318 ( 
.A(n_186),
.Y(n_318)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_191),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_192),
.Y(n_455)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_194),
.Y(n_270)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_198),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_245),
.B(n_510),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_207),
.B(n_208),
.Y(n_510)
);

BUFx24_ASAP7_75t_SL g518 ( 
.A(n_207),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_214),
.C(n_217),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_209),
.A2(n_210),
.B1(n_214),
.B2(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_214),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_217),
.B(n_470),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_232),
.C(n_240),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_218),
.B(n_453),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_228),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_219),
.B(n_228),
.Y(n_478)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_220),
.Y(n_461)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_224),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_225),
.A2(n_319),
.B(n_358),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_227),
.Y(n_326)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_229),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_232),
.B(n_240),
.Y(n_453)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_233),
.Y(n_468)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_237),
.Y(n_408)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_244),
.Y(n_433)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI311xp33_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_449),
.A3(n_486),
.B1(n_504),
.C1(n_509),
.Y(n_247)
);

AOI21x1_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_400),
.B(n_448),
.Y(n_248)
);

AO21x2_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_372),
.B(n_399),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_331),
.B(n_371),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_302),
.B(n_330),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_279),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_253),
.B(n_279),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_271),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_254),
.A2(n_271),
.B1(n_272),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_254),
.Y(n_328)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_258),
.Y(n_297)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI21xp33_ASAP7_75t_SL g343 ( 
.A1(n_262),
.A2(n_344),
.B(n_347),
.Y(n_343)
);

HAxp5_ASAP7_75t_SL g414 ( 
.A(n_262),
.B(n_415),
.CON(n_414),
.SN(n_414)
);

INVx4_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_293),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_280),
.B(n_294),
.C(n_301),
.Y(n_332)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_281),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_291),
.Y(n_390)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_300),
.B2(n_301),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_322),
.B(n_329),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_309),
.B(n_321),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_308),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_320),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_320),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx6_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_317),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_327),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_327),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_332),
.B(n_333),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_356),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_336),
.B1(n_341),
.B2(n_342),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_336),
.B(n_341),
.C(n_356),
.Y(n_373)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

AOI32xp33_ASAP7_75t_L g362 ( 
.A1(n_348),
.A2(n_363),
.A3(n_364),
.B1(n_367),
.B2(n_369),
.Y(n_362)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_350),
.Y(n_385)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx6_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_362),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_362),
.Y(n_378)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_363),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx6_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_373),
.B(n_374),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_376),
.B1(n_379),
.B2(n_398),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_377),
.B(n_378),
.C(n_398),
.Y(n_401)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_379),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_386),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_380),
.B(n_387),
.C(n_388),
.Y(n_427)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_389),
.Y(n_420)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_401),
.B(n_402),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_430),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.Y(n_403)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_404),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_406),
.B1(n_418),
.B2(n_419),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_406),
.B(n_418),
.Y(n_482)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx6_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_427),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_427),
.B(n_429),
.C(n_430),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_431),
.A2(n_432),
.B1(n_434),
.B2(n_447),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_431),
.B(n_435),
.C(n_441),
.Y(n_495)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_434),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_435),
.B(n_441),
.Y(n_434)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_436),
.Y(n_484)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx8_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

NAND2xp33_ASAP7_75t_SL g449 ( 
.A(n_450),
.B(n_472),
.Y(n_449)
);

A2O1A1Ixp33_ASAP7_75t_SL g504 ( 
.A1(n_450),
.A2(n_472),
.B(n_505),
.C(n_508),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_469),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_451),
.B(n_469),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_454),
.C(n_456),
.Y(n_451)
);

FAx1_ASAP7_75t_SL g485 ( 
.A(n_452),
.B(n_454),
.CI(n_456),
.CON(n_485),
.SN(n_485)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_464),
.C(n_467),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_458),
.B(n_460),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_458),
.B(n_460),
.Y(n_494)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_464),
.A2(n_465),
.B1(n_467),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_467),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_485),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_473),
.B(n_485),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_478),
.C(n_479),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_474),
.A2(n_475),
.B1(n_478),
.B2(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_478),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_479),
.B(n_497),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_482),
.C(n_483),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_480),
.A2(n_481),
.B1(n_483),
.B2(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_482),
.B(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_483),
.Y(n_492)
);

BUFx24_ASAP7_75t_SL g516 ( 
.A(n_485),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_487),
.B(n_499),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_488),
.A2(n_506),
.B(n_507),
.Y(n_505)
);

NOR2x1_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_496),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_489),
.B(n_496),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_493),
.C(n_495),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_490),
.B(n_502),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_493),
.A2(n_494),
.B1(n_495),
.B2(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_495),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_501),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_500),
.B(n_501),
.Y(n_506)
);

INVx8_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx8_ASAP7_75t_L g514 ( 
.A(n_512),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);


endmodule