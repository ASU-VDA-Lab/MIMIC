module fake_netlist_5_1446_n_653 (n_91, n_82, n_122, n_10, n_24, n_124, n_86, n_83, n_61, n_90, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_105, n_80, n_4, n_35, n_73, n_17, n_92, n_19, n_120, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_653);

input n_91;
input n_82;
input n_122;
input n_10;
input n_24;
input n_124;
input n_86;
input n_83;
input n_61;
input n_90;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_105;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_653;

wire n_137;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_418;
wire n_248;
wire n_136;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_619;
wire n_408;
wire n_376;
wire n_503;
wire n_127;
wire n_235;
wire n_226;
wire n_605;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_483;
wire n_544;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_139;
wire n_280;
wire n_590;
wire n_629;
wire n_378;
wire n_551;
wire n_581;
wire n_382;
wire n_554;
wire n_254;
wire n_583;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_455;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_133;
wire n_330;
wire n_508;
wire n_506;
wire n_610;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_307;
wire n_633;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_134;
wire n_191;
wire n_587;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_132;
wire n_546;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_570;
wire n_457;
wire n_514;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_131;
wire n_192;
wire n_636;
wire n_600;
wire n_223;
wire n_392;
wire n_158;
wire n_138;
wire n_264;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_415;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_584;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_129;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_638;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_309;
wire n_512;
wire n_462;
wire n_130;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_627;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_180;
wire n_560;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_572;
wire n_246;
wire n_596;
wire n_179;
wire n_125;
wire n_410;
wire n_558;
wire n_269;
wire n_529;
wire n_128;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_135;
wire n_126;
wire n_644;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_262;
wire n_238;
wire n_639;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_79),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_36),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_0),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_121),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_41),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_60),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_12),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_34),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_15),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_37),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_30),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_56),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_111),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_75),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_48),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_8),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_22),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_20),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_90),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_46),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_15),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_14),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_35),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_6),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_29),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_69),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_58),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_122),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_84),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_40),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_77),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_66),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_113),
.Y(n_166)
);

NOR2xp67_ASAP7_75t_L g167 ( 
.A(n_14),
.B(n_100),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_44),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_67),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_70),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_83),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_42),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_54),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_112),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_57),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

AND2x4_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_129),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

OA21x2_ASAP7_75t_L g187 ( 
.A1(n_136),
.A2(n_0),
.B(n_1),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_134),
.A2(n_152),
.B1(n_143),
.B2(n_156),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_167),
.B(n_1),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_125),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_130),
.B(n_2),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g196 ( 
.A1(n_150),
.A2(n_2),
.B(n_3),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

AOI22x1_ASAP7_75t_SL g198 ( 
.A1(n_132),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

NOR2x1_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_17),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_139),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_127),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_131),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_175),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

NAND2xp33_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_168),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_192),
.B(n_142),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_189),
.A2(n_165),
.B1(n_169),
.B2(n_166),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_207),
.Y(n_226)
);

NAND2xp33_ASAP7_75t_SL g227 ( 
.A(n_195),
.B(n_138),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_140),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

INVxp67_ASAP7_75t_SL g233 ( 
.A(n_176),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_172),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_182),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_141),
.Y(n_237)
);

INVxp33_ASAP7_75t_SL g238 ( 
.A(n_194),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_145),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_185),
.B(n_146),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_185),
.B(n_149),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_182),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_197),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_209),
.B(n_153),
.Y(n_248)
);

NAND2xp33_ASAP7_75t_L g249 ( 
.A(n_176),
.B(n_157),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_185),
.B(n_159),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_185),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_197),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_176),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_176),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_203),
.Y(n_256)
);

NOR2x1p5_ASAP7_75t_L g257 ( 
.A(n_186),
.B(n_161),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_179),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_258),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_258),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_177),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_177),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_224),
.A2(n_206),
.B1(n_183),
.B2(n_207),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_217),
.B(n_183),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_218),
.B(n_183),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_215),
.B(n_177),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_216),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_177),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_186),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_204),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_204),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_219),
.Y(n_276)
);

A2O1A1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_227),
.A2(n_212),
.B(n_213),
.C(n_180),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_227),
.A2(n_196),
.B1(n_187),
.B2(n_203),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_236),
.B(n_200),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_235),
.B(n_203),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_225),
.B(n_162),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_248),
.B(n_181),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_257),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_236),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_180),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_251),
.B(n_181),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_255),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_241),
.B(n_242),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_244),
.B(n_179),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_241),
.B(n_242),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_221),
.B(n_191),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_221),
.B(n_191),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_224),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_220),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_231),
.B(n_191),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_231),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_232),
.Y(n_300)
);

O2A1O1Ixp33_ASAP7_75t_L g301 ( 
.A1(n_222),
.A2(n_212),
.B(n_196),
.C(n_187),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_232),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_238),
.B(n_191),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_223),
.B(n_184),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_229),
.B(n_184),
.Y(n_305)
);

OAI22x1_ASAP7_75t_SL g306 ( 
.A1(n_238),
.A2(n_198),
.B1(n_5),
.B2(n_6),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_245),
.B(n_188),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_246),
.B(n_188),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_234),
.Y(n_309)
);

NAND2xp33_ASAP7_75t_L g310 ( 
.A(n_234),
.B(n_199),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g311 ( 
.A(n_240),
.B(n_199),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_243),
.B(n_201),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_230),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_281),
.A2(n_264),
.B(n_283),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_259),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_296),
.A2(n_249),
.B1(n_187),
.B2(n_196),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_271),
.B(n_303),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_285),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_301),
.A2(n_214),
.B(n_208),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_266),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_288),
.A2(n_230),
.B(n_73),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_274),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_272),
.B(n_230),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_260),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_266),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_262),
.A2(n_230),
.B(n_74),
.Y(n_330)
);

AO21x1_ASAP7_75t_L g331 ( 
.A1(n_282),
.A2(n_198),
.B(n_7),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_265),
.B(n_4),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_294),
.A2(n_298),
.B(n_295),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_291),
.A2(n_71),
.B(n_124),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_280),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_293),
.A2(n_279),
.B1(n_284),
.B2(n_292),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_289),
.B(n_18),
.Y(n_337)
);

CKINVDCx8_ASAP7_75t_R g338 ( 
.A(n_306),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_279),
.B(n_7),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_268),
.A2(n_76),
.B(n_123),
.Y(n_340)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_274),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_19),
.Y(n_342)
);

BUFx4f_ASAP7_75t_L g343 ( 
.A(n_284),
.Y(n_343)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_267),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_292),
.B(n_21),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_267),
.B(n_8),
.Y(n_346)
);

NAND2x1_ASAP7_75t_L g347 ( 
.A(n_260),
.B(n_23),
.Y(n_347)
);

AOI21x1_ASAP7_75t_L g348 ( 
.A1(n_304),
.A2(n_78),
.B(n_119),
.Y(n_348)
);

NOR2x1_ASAP7_75t_L g349 ( 
.A(n_270),
.B(n_24),
.Y(n_349)
);

AOI21xp33_ASAP7_75t_L g350 ( 
.A1(n_278),
.A2(n_9),
.B(n_10),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_312),
.A2(n_80),
.B(n_118),
.Y(n_351)
);

NOR2x1_ASAP7_75t_L g352 ( 
.A(n_277),
.B(n_25),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_273),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_297),
.A2(n_82),
.B1(n_117),
.B2(n_116),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_290),
.B(n_26),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_309),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_275),
.A2(n_81),
.B1(n_115),
.B2(n_110),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_305),
.A2(n_68),
.B(n_109),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_290),
.B(n_11),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_263),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_269),
.B(n_65),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_307),
.A2(n_308),
.B(n_310),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_261),
.A2(n_64),
.B(n_107),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_276),
.A2(n_63),
.B(n_106),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_L g365 ( 
.A(n_276),
.B(n_62),
.Y(n_365)
);

AO31x2_ASAP7_75t_L g366 ( 
.A1(n_359),
.A2(n_302),
.A3(n_300),
.B(n_299),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_324),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_318),
.B(n_286),
.Y(n_368)
);

OAI21x1_ASAP7_75t_L g369 ( 
.A1(n_333),
.A2(n_286),
.B(n_313),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_321),
.A2(n_61),
.B(n_105),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_314),
.A2(n_59),
.B(n_104),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_323),
.B(n_13),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_319),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_335),
.Y(n_374)
);

AO31x2_ASAP7_75t_L g375 ( 
.A1(n_339),
.A2(n_13),
.A3(n_16),
.B(n_27),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_319),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_315),
.Y(n_377)
);

NAND2x1p5_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_28),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_338),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_316),
.A2(n_38),
.B(n_39),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_329),
.B(n_43),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_362),
.A2(n_45),
.B(n_47),
.Y(n_382)
);

A2O1A1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_350),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_326),
.B(n_52),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_344),
.B(n_53),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_327),
.A2(n_345),
.B(n_322),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_322),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_328),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_341),
.B(n_86),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_320),
.B(n_87),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_343),
.Y(n_391)
);

AOI21xp33_ASAP7_75t_L g392 ( 
.A1(n_332),
.A2(n_91),
.B(n_92),
.Y(n_392)
);

NAND2x1p5_ASAP7_75t_L g393 ( 
.A(n_341),
.B(n_93),
.Y(n_393)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_356),
.A2(n_95),
.B(n_96),
.Y(n_394)
);

OAI21x1_ASAP7_75t_L g395 ( 
.A1(n_360),
.A2(n_97),
.B(n_98),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_317),
.A2(n_99),
.B(n_101),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_360),
.A2(n_102),
.B(n_103),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_346),
.B(n_353),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_363),
.A2(n_342),
.B(n_337),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_343),
.B(n_331),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_354),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_352),
.B(n_358),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_365),
.A2(n_361),
.B(n_325),
.Y(n_403)
);

OAI21x1_ASAP7_75t_L g404 ( 
.A1(n_330),
.A2(n_348),
.B(n_334),
.Y(n_404)
);

OAI21x1_ASAP7_75t_L g405 ( 
.A1(n_347),
.A2(n_364),
.B(n_351),
.Y(n_405)
);

AOI21x1_ASAP7_75t_L g406 ( 
.A1(n_349),
.A2(n_340),
.B(n_357),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_344),
.B(n_318),
.Y(n_407)
);

OAI21x1_ASAP7_75t_L g408 ( 
.A1(n_369),
.A2(n_404),
.B(n_405),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_367),
.Y(n_409)
);

OAI21x1_ASAP7_75t_L g410 ( 
.A1(n_403),
.A2(n_386),
.B(n_406),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_368),
.B(n_374),
.Y(n_411)
);

OAI21x1_ASAP7_75t_L g412 ( 
.A1(n_394),
.A2(n_395),
.B(n_397),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_388),
.Y(n_413)
);

AO21x2_ASAP7_75t_L g414 ( 
.A1(n_380),
.A2(n_399),
.B(n_370),
.Y(n_414)
);

AO21x2_ASAP7_75t_L g415 ( 
.A1(n_380),
.A2(n_371),
.B(n_382),
.Y(n_415)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_373),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_384),
.Y(n_417)
);

OAI21x1_ASAP7_75t_L g418 ( 
.A1(n_402),
.A2(n_396),
.B(n_385),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_377),
.B(n_398),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_400),
.A2(n_407),
.B1(n_384),
.B2(n_389),
.Y(n_420)
);

AOI21x1_ASAP7_75t_L g421 ( 
.A1(n_388),
.A2(n_401),
.B(n_381),
.Y(n_421)
);

INVx5_ASAP7_75t_L g422 ( 
.A(n_373),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g423 ( 
.A1(n_387),
.A2(n_393),
.B(n_378),
.Y(n_423)
);

AO31x2_ASAP7_75t_L g424 ( 
.A1(n_383),
.A2(n_366),
.A3(n_375),
.B(n_392),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_387),
.B(n_376),
.Y(n_425)
);

OAI21x1_ASAP7_75t_L g426 ( 
.A1(n_390),
.A2(n_372),
.B(n_366),
.Y(n_426)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_366),
.A2(n_373),
.B(n_376),
.Y(n_427)
);

NAND2x1p5_ASAP7_75t_L g428 ( 
.A(n_376),
.B(n_377),
.Y(n_428)
);

AO21x1_ASAP7_75t_L g429 ( 
.A1(n_375),
.A2(n_379),
.B(n_391),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_375),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_379),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_377),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_L g433 ( 
.A1(n_380),
.A2(n_350),
.B1(n_339),
.B2(n_370),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_384),
.Y(n_434)
);

OAI21xp33_ASAP7_75t_L g435 ( 
.A1(n_377),
.A2(n_282),
.B(n_224),
.Y(n_435)
);

AO21x2_ASAP7_75t_L g436 ( 
.A1(n_380),
.A2(n_399),
.B(n_370),
.Y(n_436)
);

OAI21x1_ASAP7_75t_L g437 ( 
.A1(n_369),
.A2(n_405),
.B(n_404),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_377),
.Y(n_438)
);

CKINVDCx11_ASAP7_75t_R g439 ( 
.A(n_377),
.Y(n_439)
);

OAI21x1_ASAP7_75t_L g440 ( 
.A1(n_369),
.A2(n_405),
.B(n_404),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_377),
.B(n_259),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_369),
.A2(n_404),
.B(n_405),
.Y(n_442)
);

NAND2x1p5_ASAP7_75t_L g443 ( 
.A(n_373),
.B(n_376),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_413),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_439),
.Y(n_445)
);

OAI22xp33_ASAP7_75t_L g446 ( 
.A1(n_431),
.A2(n_420),
.B1(n_438),
.B2(n_434),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_427),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_432),
.Y(n_448)
);

AO21x2_ASAP7_75t_L g449 ( 
.A1(n_415),
.A2(n_436),
.B(n_414),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_441),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_428),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_417),
.B(n_434),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_416),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_419),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_409),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_411),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_411),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_430),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_419),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_428),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_430),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_417),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_425),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_421),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_416),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_439),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_425),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_416),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_410),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_431),
.A2(n_433),
.B1(n_415),
.B2(n_429),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_416),
.B(n_422),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_433),
.B(n_426),
.Y(n_472)
);

CKINVDCx10_ASAP7_75t_R g473 ( 
.A(n_422),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_443),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_408),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_422),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_442),
.Y(n_477)
);

BUFx4f_ASAP7_75t_SL g478 ( 
.A(n_422),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_456),
.B(n_424),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_424),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_457),
.B(n_424),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_457),
.B(n_467),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_459),
.B(n_443),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_458),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_418),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_467),
.B(n_424),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_450),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_471),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_458),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_461),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_444),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_461),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_473),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_463),
.B(n_414),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_448),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_451),
.Y(n_496)
);

BUFx2_ASAP7_75t_SL g497 ( 
.A(n_471),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_451),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_455),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_470),
.B(n_423),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_460),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_460),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_473),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_464),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_446),
.B(n_436),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_472),
.B(n_412),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_447),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_452),
.B(n_437),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_449),
.B(n_440),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_462),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_452),
.B(n_474),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_487),
.B(n_452),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_504),
.Y(n_513)
);

AND2x4_ASAP7_75t_SL g514 ( 
.A(n_501),
.B(n_452),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_484),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_482),
.B(n_466),
.Y(n_516)
);

OAI22xp33_ASAP7_75t_L g517 ( 
.A1(n_505),
.A2(n_466),
.B1(n_445),
.B2(n_478),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_496),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_484),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_488),
.Y(n_520)
);

OR2x6_ASAP7_75t_L g521 ( 
.A(n_497),
.B(n_469),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_485),
.B(n_468),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_495),
.B(n_449),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_486),
.B(n_449),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_496),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_489),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_486),
.B(n_481),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_493),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_498),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_489),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_492),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_483),
.B(n_445),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_504),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_488),
.B(n_476),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_494),
.B(n_477),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_492),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_490),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_479),
.B(n_477),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_500),
.A2(n_465),
.B1(n_453),
.B2(n_468),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_498),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_480),
.B(n_475),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_511),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_499),
.B(n_476),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_480),
.B(n_475),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_515),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_527),
.B(n_506),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_513),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_513),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_519),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_533),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_523),
.B(n_509),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_527),
.B(n_506),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_526),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_524),
.B(n_509),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_518),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_521),
.B(n_508),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_530),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_521),
.B(n_508),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_531),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_542),
.B(n_540),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_521),
.B(n_536),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_537),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_541),
.B(n_544),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_532),
.B(n_510),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_535),
.B(n_507),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_560),
.B(n_522),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_547),
.Y(n_567)
);

NOR2x1p5_ASAP7_75t_L g568 ( 
.A(n_554),
.B(n_516),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_555),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_546),
.B(n_544),
.Y(n_570)
);

INVxp33_ASAP7_75t_L g571 ( 
.A(n_564),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_546),
.B(n_541),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_547),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_548),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_561),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_552),
.B(n_538),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_561),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_552),
.B(n_517),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_548),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_573),
.B(n_551),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_577),
.B(n_575),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_577),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_567),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_567),
.Y(n_584)
);

AND3x2_ASAP7_75t_L g585 ( 
.A(n_578),
.B(n_529),
.C(n_502),
.Y(n_585)
);

OAI22xp33_ASAP7_75t_L g586 ( 
.A1(n_571),
.A2(n_520),
.B1(n_522),
.B2(n_521),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_573),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_574),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_569),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_586),
.A2(n_568),
.B1(n_566),
.B2(n_575),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_585),
.A2(n_577),
.B1(n_556),
.B2(n_558),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_587),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_589),
.A2(n_554),
.B1(n_569),
.B2(n_551),
.Y(n_593)
);

A2O1A1Ixp33_ASAP7_75t_L g594 ( 
.A1(n_589),
.A2(n_503),
.B(n_493),
.C(n_528),
.Y(n_594)
);

AOI221xp5_ASAP7_75t_L g595 ( 
.A1(n_593),
.A2(n_580),
.B1(n_588),
.B2(n_562),
.C(n_583),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_591),
.B(n_581),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_594),
.B(n_528),
.Y(n_597)
);

O2A1O1Ixp33_ASAP7_75t_L g598 ( 
.A1(n_592),
.A2(n_580),
.B(n_503),
.C(n_512),
.Y(n_598)
);

AOI221x1_ASAP7_75t_L g599 ( 
.A1(n_590),
.A2(n_581),
.B1(n_579),
.B2(n_574),
.C(n_584),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_591),
.B(n_582),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_600),
.A2(n_556),
.B(n_558),
.Y(n_601)
);

AOI221xp5_ASAP7_75t_L g602 ( 
.A1(n_595),
.A2(n_579),
.B1(n_549),
.B2(n_557),
.C(n_553),
.Y(n_602)
);

NOR3xp33_ASAP7_75t_L g603 ( 
.A(n_596),
.B(n_597),
.C(n_598),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_599),
.A2(n_556),
.B1(n_558),
.B2(n_561),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_603),
.B(n_572),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_602),
.B(n_572),
.Y(n_606)
);

AOI211xp5_ASAP7_75t_L g607 ( 
.A1(n_601),
.A2(n_525),
.B(n_520),
.C(n_559),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_605),
.Y(n_608)
);

NOR2x1_ASAP7_75t_SL g609 ( 
.A(n_606),
.B(n_607),
.Y(n_609)
);

XOR2x1_ASAP7_75t_L g610 ( 
.A(n_605),
.B(n_471),
.Y(n_610)
);

NOR2x1_ASAP7_75t_L g611 ( 
.A(n_605),
.B(n_465),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_608),
.Y(n_612)
);

NOR2x1_ASAP7_75t_L g613 ( 
.A(n_611),
.B(n_465),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_609),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_610),
.Y(n_615)
);

NOR2x1_ASAP7_75t_L g616 ( 
.A(n_611),
.B(n_471),
.Y(n_616)
);

NAND4xp75_ASAP7_75t_L g617 ( 
.A(n_611),
.B(n_604),
.C(n_545),
.D(n_500),
.Y(n_617)
);

AOI211x1_ASAP7_75t_L g618 ( 
.A1(n_609),
.A2(n_570),
.B(n_576),
.C(n_563),
.Y(n_618)
);

NOR2xp67_ASAP7_75t_L g619 ( 
.A(n_614),
.B(n_525),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_615),
.A2(n_612),
.B1(n_617),
.B2(n_613),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_618),
.Y(n_621)
);

AND2x2_ASAP7_75t_SL g622 ( 
.A(n_616),
.B(n_453),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_612),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_612),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_614),
.A2(n_520),
.B1(n_534),
.B2(n_514),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_614),
.Y(n_626)
);

OAI22x1_ASAP7_75t_L g627 ( 
.A1(n_626),
.A2(n_624),
.B1(n_620),
.B2(n_623),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_622),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_621),
.A2(n_534),
.B1(n_520),
.B2(n_514),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_619),
.A2(n_539),
.B1(n_565),
.B2(n_570),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_625),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_626),
.B(n_576),
.Y(n_632)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_626),
.B(n_534),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_626),
.B(n_488),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_632),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_627),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_633),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_634),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_628),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_631),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_629),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_636),
.A2(n_630),
.B1(n_565),
.B2(n_550),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_640),
.A2(n_453),
.B1(n_468),
.B2(n_497),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_639),
.A2(n_641),
.B1(n_637),
.B2(n_638),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_638),
.A2(n_635),
.B(n_543),
.Y(n_645)
);

AO21x2_ASAP7_75t_L g646 ( 
.A1(n_645),
.A2(n_499),
.B(n_491),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_644),
.A2(n_453),
.B1(n_468),
.B2(n_476),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_642),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_646),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_648),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_650),
.B(n_647),
.Y(n_651)
);

OR2x6_ASAP7_75t_L g652 ( 
.A(n_651),
.B(n_649),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_652),
.A2(n_643),
.B1(n_453),
.B2(n_468),
.Y(n_653)
);


endmodule