module real_jpeg_27216_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_334, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_334;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_0),
.A2(n_27),
.B1(n_35),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_0),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_0),
.A2(n_31),
.B1(n_33),
.B2(n_121),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_0),
.A2(n_46),
.B1(n_47),
.B2(n_121),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_0),
.A2(n_62),
.B1(n_64),
.B2(n_121),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_1),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_1),
.B(n_30),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_1),
.B(n_33),
.Y(n_221)
);

AOI21xp33_ASAP7_75t_L g225 ( 
.A1(n_1),
.A2(n_33),
.B(n_221),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_180),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_1),
.A2(n_59),
.B(n_62),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_1),
.B(n_87),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_1),
.A2(n_109),
.B1(n_127),
.B2(n_269),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_2),
.Y(n_104)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_2),
.Y(n_109)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_2),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_3),
.A2(n_27),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_3),
.A2(n_31),
.B1(n_33),
.B2(n_38),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_3),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_3),
.A2(n_38),
.B1(n_62),
.B2(n_64),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_7),
.A2(n_27),
.B1(n_35),
.B2(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_7),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_7),
.A2(n_31),
.B1(n_33),
.B2(n_182),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_182),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_7),
.A2(n_62),
.B1(n_64),
.B2(n_182),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_8),
.A2(n_27),
.B1(n_35),
.B2(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_8),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_8),
.A2(n_31),
.B1(n_33),
.B2(n_148),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_148),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_8),
.A2(n_62),
.B1(n_64),
.B2(n_148),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_9),
.A2(n_31),
.B1(n_33),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_9),
.A2(n_27),
.B1(n_35),
.B2(n_53),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_9),
.A2(n_53),
.B1(n_62),
.B2(n_64),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_10),
.A2(n_31),
.B1(n_33),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_10),
.A2(n_50),
.B1(n_62),
.B2(n_64),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_10),
.A2(n_27),
.B1(n_35),
.B2(n_50),
.Y(n_123)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_13),
.A2(n_31),
.B1(n_33),
.B2(n_48),
.Y(n_55)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_13),
.Y(n_220)
);

INVx11_ASAP7_75t_SL g63 ( 
.A(n_14),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_15),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_15),
.A2(n_36),
.B1(n_46),
.B2(n_47),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_15),
.A2(n_31),
.B1(n_33),
.B2(n_36),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_15),
.A2(n_36),
.B1(n_62),
.B2(n_64),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_94),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_79),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_19),
.B(n_79),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_69),
.C(n_73),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_20),
.A2(n_21),
.B1(n_69),
.B2(n_320),
.Y(n_324)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_40),
.B1(n_41),
.B2(n_68),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_22),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_23),
.A2(n_120),
.B(n_122),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_23),
.A2(n_39),
.B1(n_120),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_23),
.A2(n_39),
.B1(n_147),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_24),
.B(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_24),
.A2(n_83),
.B(n_84),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_24),
.A2(n_84),
.B(n_123),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_24),
.A2(n_30),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_25),
.B(n_33),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g179 ( 
.A(n_27),
.B(n_180),
.CON(n_179),
.SN(n_179)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_29),
.A2(n_31),
.B1(n_179),
.B2(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_30),
.B(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

AOI32xp33_ASAP7_75t_L g217 ( 
.A1(n_31),
.A2(n_46),
.A3(n_218),
.B1(n_221),
.B2(n_222),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_34),
.A2(n_39),
.B(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_37),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_39),
.B(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_56),
.B2(n_67),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_56),
.C(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_51),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_44),
.A2(n_75),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_45),
.A2(n_54),
.B1(n_77),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_45),
.A2(n_54),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_45),
.A2(n_54),
.B1(n_176),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_45),
.A2(n_54),
.B1(n_204),
.B2(n_225),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_47),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g222 ( 
.A(n_47),
.B(n_219),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_47),
.A2(n_60),
.B(n_180),
.C(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_51),
.A2(n_87),
.B(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_56),
.A2(n_67),
.B1(n_74),
.B2(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_61),
.B(n_65),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_57),
.A2(n_61),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_57),
.A2(n_113),
.B(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_57),
.A2(n_65),
.B(n_131),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_57),
.A2(n_61),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_57),
.A2(n_154),
.B(n_229),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_57),
.A2(n_61),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_57),
.A2(n_61),
.B1(n_228),
.B2(n_246),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_64),
.Y(n_61)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_61),
.A2(n_112),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_61),
.B(n_180),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_62),
.Y(n_64)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_64),
.B(n_273),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_66),
.B(n_133),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_69),
.C(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_69),
.A2(n_317),
.B1(n_319),
.B2(n_320),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_69),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_73),
.B(n_324),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_74),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B(n_78),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_75),
.A2(n_78),
.B(n_88),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_85),
.B2(n_86),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI321xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_313),
.A3(n_325),
.B1(n_331),
.B2(n_332),
.C(n_334),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_165),
.B(n_312),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_149),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_97),
.B(n_149),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_124),
.C(n_135),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_98),
.A2(n_99),
.B1(n_124),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_114),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_100),
.B(n_116),
.C(n_118),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_111),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_101),
.B(n_111),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_102),
.A2(n_195),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_103),
.A2(n_110),
.B(n_140),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_103),
.A2(n_108),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_128),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_107),
.A2(n_127),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

INVx11_ASAP7_75t_L g208 ( 
.A(n_108),
.Y(n_208)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_109),
.A2(n_127),
.B1(n_138),
.B2(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_110),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_117),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_124),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_134),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_125),
.A2(n_126),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_130),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_126),
.A2(n_159),
.B(n_162),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B(n_129),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_138),
.B(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_127),
.A2(n_208),
.B1(n_261),
.B2(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_130),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_132),
.B(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_135),
.B(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_144),
.C(n_145),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_136),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_141),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_144),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_163),
.B2(n_164),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_158),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_152),
.B(n_158),
.C(n_164),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_155),
.B(n_157),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_155),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_157),
.B(n_315),
.C(n_321),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_157),
.A2(n_315),
.B1(n_316),
.B2(n_330),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_157),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_163),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_306),
.B(n_311),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_209),
.B(n_292),
.C(n_305),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_196),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_168),
.B(n_196),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_183),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_170),
.B(n_171),
.C(n_183),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.C(n_178),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_178),
.B(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_180),
.B(n_208),
.Y(n_273)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_191),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_185),
.B(n_189),
.C(n_191),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_194),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.C(n_202),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_197),
.A2(n_198),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_202),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.C(n_207),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_207),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_291),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_284),
.B(n_290),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_239),
.B(n_283),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_230),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_213),
.B(n_230),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_223),
.C(n_226),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_214),
.A2(n_215),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_217),
.Y(n_237)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_235),
.B2(n_236),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_231),
.B(n_237),
.C(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_277),
.B(n_282),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_257),
.B(n_276),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_249),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_242),
.B(n_249),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_243),
.A2(n_244),
.B1(n_247),
.B2(n_264),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_247),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_255),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_254),
.C(n_255),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_256),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_265),
.B(n_275),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_263),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_259),
.B(n_263),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_270),
.B(n_274),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_267),
.B(n_268),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_285),
.B(n_286),
.Y(n_290)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_293),
.B(n_294),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_303),
.B2(n_304),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_300),
.C(n_304),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_303),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_323),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_323),
.Y(n_332)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_321),
.A2(n_322),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_326),
.B(n_327),
.Y(n_331)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);


endmodule