module fake_jpeg_15309_n_189 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_189);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_37),
.Y(n_70)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_40),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_19),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_32),
.B1(n_31),
.B2(n_45),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_65),
.B(n_72),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_57),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_63),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_17),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_16),
.B(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_46),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_35),
.A2(n_31),
.B1(n_33),
.B2(n_28),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_23),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_24),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_3),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_39),
.A2(n_31),
.B1(n_33),
.B2(n_28),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_78),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_86),
.Y(n_104)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_17),
.A3(n_43),
.B1(n_22),
.B2(n_21),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_81),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_25),
.Y(n_78)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_26),
.B1(n_24),
.B2(n_27),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_30),
.B(n_6),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_59),
.A2(n_26),
.B1(n_21),
.B2(n_18),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_5),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_25),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_93),
.Y(n_101)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_2),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_3),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_30),
.B1(n_4),
.B2(n_5),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_5),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_15),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

AND2x4_ASAP7_75t_SL g105 ( 
.A(n_73),
.B(n_89),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_119),
.B(n_30),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_113),
.B1(n_91),
.B2(n_83),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_79),
.C(n_85),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_118),
.C(n_51),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_114),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_117),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_71),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_57),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_74),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_49),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_51),
.C(n_50),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_87),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_123),
.B(n_126),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_134),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_97),
.B1(n_82),
.B2(n_94),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_128),
.B1(n_137),
.B2(n_106),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_103),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_91),
.B(n_50),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_136),
.C(n_115),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_97),
.B1(n_82),
.B2(n_83),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_76),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_133),
.B(n_135),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_74),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_99),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_50),
.Y(n_135)
);

XNOR2x1_ASAP7_75t_SL g136 ( 
.A(n_101),
.B(n_81),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_152),
.B1(n_128),
.B2(n_126),
.Y(n_157)
);

NOR2x1_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_104),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_139),
.A2(n_140),
.B(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_102),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_146),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_119),
.B1(n_107),
.B2(n_102),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_104),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_100),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_116),
.B1(n_113),
.B2(n_119),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_160),
.B1(n_138),
.B2(n_150),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_135),
.C(n_130),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_151),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_156),
.A2(n_139),
.B(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_157),
.B(n_150),
.Y(n_168)
);

BUFx24_ASAP7_75t_SL g159 ( 
.A(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_141),
.Y(n_171)
);

OAI321xp33_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_132),
.A3(n_111),
.B1(n_116),
.B2(n_109),
.C(n_98),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_146),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_144),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_167),
.C(n_169),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_165),
.A2(n_166),
.B(n_170),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_158),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_147),
.B(n_145),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_171),
.B(n_109),
.Y(n_176)
);

AOI321xp33_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_153),
.A3(n_158),
.B1(n_161),
.B2(n_162),
.C(n_154),
.Y(n_174)
);

AOI211xp5_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_175),
.B(n_14),
.C(n_8),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_176),
.B(n_7),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_55),
.C(n_52),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_170),
.C(n_165),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_179),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_52),
.C(n_98),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_182),
.B(n_7),
.Y(n_184)
);

AOI322xp5_ASAP7_75t_L g185 ( 
.A1(n_181),
.A2(n_7),
.A3(n_8),
.B1(n_10),
.B2(n_11),
.C1(n_75),
.C2(n_179),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_173),
.A2(n_75),
.B1(n_14),
.B2(n_9),
.Y(n_182)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_11),
.B(n_8),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_10),
.B1(n_183),
.B2(n_187),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_10),
.Y(n_189)
);


endmodule