module fake_jpeg_32084_n_122 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_122);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_0),
.B(n_37),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_59),
.Y(n_61)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_47),
.Y(n_69)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_48),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_73),
.B(n_52),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_58),
.A2(n_48),
.B1(n_51),
.B2(n_50),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_51),
.B1(n_41),
.B2(n_43),
.Y(n_74)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_49),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_71),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_74),
.A2(n_86),
.B(n_9),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_84),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_47),
.B(n_21),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_78),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_10),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_20),
.C(n_39),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_82),
.C(n_18),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_19),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_85),
.Y(n_100)
);

AO22x1_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_24),
.B1(n_36),
.B2(n_35),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_4),
.C(n_5),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_12),
.B1(n_14),
.B2(n_17),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_76),
.A2(n_64),
.B1(n_70),
.B2(n_7),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_94),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_9),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_64),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_96),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_104),
.B(n_28),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_99),
.B(n_101),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_80),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_103),
.C(n_27),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_22),
.C(n_25),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_112),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_78),
.C(n_29),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_100),
.C(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_109),
.A2(n_100),
.B1(n_90),
.B2(n_99),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_107),
.B(n_111),
.Y(n_116)
);

OAI211xp5_ASAP7_75t_L g118 ( 
.A1(n_116),
.A2(n_107),
.B(n_108),
.C(n_113),
.Y(n_118)
);

OAI21x1_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_114),
.B(n_117),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_106),
.C(n_32),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_30),
.C(n_33),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_34),
.Y(n_122)
);


endmodule