module fake_jpeg_190_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_52),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_36),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_41),
.B1(n_36),
.B2(n_39),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_56),
.B1(n_53),
.B2(n_50),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_50),
.A2(n_41),
.B1(n_45),
.B2(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_63),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_45),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_69),
.Y(n_77)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_49),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_51),
.B(n_50),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_58),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_75),
.B1(n_58),
.B2(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_34),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_34),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_46),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_38),
.Y(n_76)
);

A2O1A1O1Ixp25_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_0),
.B(n_2),
.C(n_3),
.D(n_4),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_79),
.B1(n_71),
.B2(n_66),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_56),
.B1(n_52),
.B2(n_48),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_88),
.B(n_81),
.C(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_82),
.B(n_85),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_63),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_5),
.C(n_7),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_46),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_59),
.B(n_43),
.C(n_52),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_59),
.B(n_68),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_48),
.B1(n_36),
.B2(n_42),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_94),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_84),
.A2(n_81),
.B1(n_77),
.B2(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_65),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_28),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_43),
.C(n_42),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_95),
.C(n_96),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_72),
.B(n_2),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_98),
.Y(n_103)
);

OAI32xp33_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_99)
);

AOI322xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_16),
.C2(n_18),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_8),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_100),
.Y(n_111)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

NAND2xp67_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_24),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_104),
.B(n_111),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_112),
.B1(n_114),
.B2(n_108),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_25),
.C(n_31),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_103),
.C(n_107),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_27),
.A3(n_30),
.B1(n_29),
.B2(n_20),
.C1(n_26),
.C2(n_32),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_113),
.Y(n_118)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_119),
.C(n_110),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_109),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_94),
.C(n_93),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_120),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_119),
.C(n_116),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_124),
.B(n_125),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_118),
.C(n_122),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_106),
.C(n_104),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_94),
.C(n_14),
.Y(n_130)
);

BUFx24_ASAP7_75t_SL g131 ( 
.A(n_130),
.Y(n_131)
);


endmodule