module fake_netlist_6_1682_n_39 (n_7, n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_8, n_39);

input n_7;
input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;
input n_8;

output n_39;

wire n_16;
wire n_34;
wire n_9;
wire n_18;
wire n_21;
wire n_24;
wire n_10;
wire n_37;
wire n_15;
wire n_33;
wire n_27;
wire n_14;
wire n_38;
wire n_32;
wire n_36;
wire n_22;
wire n_26;
wire n_13;
wire n_35;
wire n_11;
wire n_28;
wire n_17;
wire n_23;
wire n_12;
wire n_20;
wire n_30;
wire n_19;
wire n_29;
wire n_31;
wire n_25;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

AND2x2_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_2),
.Y(n_10)
);

CKINVDCx5p33_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

OR2x4_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

AND2x6_ASAP7_75t_SL g21 ( 
.A(n_12),
.B(n_1),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_17),
.A2(n_11),
.B1(n_10),
.B2(n_14),
.Y(n_22)
);

CKINVDCx11_ASAP7_75t_R g23 ( 
.A(n_21),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_17),
.B1(n_11),
.B2(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

AOI221xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_18),
.B1(n_20),
.B2(n_19),
.C(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_16),
.B1(n_20),
.B2(n_17),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_3),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_28),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

AOI221xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_31),
.B1(n_5),
.B2(n_4),
.C(n_8),
.Y(n_35)
);

AO22x2_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_31),
.B1(n_5),
.B2(n_4),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_37),
.B1(n_36),
.B2(n_7),
.Y(n_39)
);


endmodule