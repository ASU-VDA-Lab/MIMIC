module real_jpeg_25726_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_0),
.A2(n_12),
.B1(n_13),
.B2(n_19),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_12),
.B1(n_13),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_4),
.B(n_10),
.Y(n_9)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_4),
.A2(n_12),
.B1(n_13),
.B2(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_4),
.B(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

XOR2xp5_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_24),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_15),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_9),
.B(n_12),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_10),
.B(n_18),
.Y(n_17)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_12),
.A2(n_13),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

INVx6_ASAP7_75t_SL g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_20),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_23),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_26),
.B(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);


endmodule