module fake_jpeg_17546_n_58 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_58);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_58;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_19),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_36),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_25),
.Y(n_35)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

AO21x1_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_38),
.B(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_30),
.C(n_26),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_38),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_28),
.B1(n_25),
.B2(n_10),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_45),
.B1(n_36),
.B2(n_1),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_7),
.B1(n_21),
.B2(n_20),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.C(n_50),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

INVxp33_ASAP7_75t_SL g52 ( 
.A(n_49),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_0),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_41),
.B1(n_47),
.B2(n_46),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_51),
.B1(n_46),
.B2(n_43),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_43),
.C(n_1),
.Y(n_55)
);

AOI322xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_0),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_56)
);

AO21x1_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_11),
.B(n_15),
.Y(n_57)
);

A2O1A1O1Ixp25_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_16),
.B(n_22),
.C(n_2),
.D(n_3),
.Y(n_58)
);


endmodule