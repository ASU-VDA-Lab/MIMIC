module fake_jpeg_3520_n_543 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_543);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_543;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_455;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_11),
.B(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_12),
.B(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx8_ASAP7_75t_SL g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_44),
.B(n_51),
.Y(n_129)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_48),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_50),
.Y(n_131)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_52),
.B(n_59),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVxp67_ASAP7_75t_SL g109 ( 
.A(n_53),
.Y(n_109)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_57),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_64),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_62),
.B(n_70),
.Y(n_155)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g114 ( 
.A(n_63),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_21),
.B(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_21),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_17),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_71),
.B(n_72),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_22),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_25),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_73),
.Y(n_123)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_76),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_77),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_35),
.B(n_7),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_35),
.B(n_7),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_37),
.B(n_1),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_1),
.Y(n_119)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_87),
.Y(n_151)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_89),
.B(n_99),
.Y(n_163)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_26),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_16),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_105),
.B(n_133),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_61),
.B(n_36),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_110),
.A2(n_111),
.B(n_39),
.Y(n_177)
);

HAxp5_ASAP7_75t_SL g111 ( 
.A(n_64),
.B(n_73),
.CON(n_111),
.SN(n_111)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_119),
.B(n_15),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

INVx11_ASAP7_75t_L g197 ( 
.A(n_121),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_54),
.A2(n_42),
.B1(n_38),
.B2(n_39),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_127),
.A2(n_20),
.B1(n_29),
.B2(n_16),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_90),
.A2(n_38),
.B1(n_36),
.B2(n_16),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_47),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_78),
.Y(n_133)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

INVx11_ASAP7_75t_L g142 ( 
.A(n_49),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_46),
.A2(n_15),
.B1(n_29),
.B2(n_20),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_93),
.B1(n_76),
.B2(n_18),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_57),
.Y(n_150)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_65),
.Y(n_160)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_53),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_66),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_100),
.B(n_45),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_164),
.B(n_167),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_166),
.B(n_177),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_55),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_170),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_56),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g227 ( 
.A1(n_171),
.A2(n_142),
.B1(n_140),
.B2(n_113),
.Y(n_227)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_104),
.Y(n_175)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_114),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_176),
.B(n_181),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_111),
.A2(n_69),
.B1(n_67),
.B2(n_36),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_178),
.A2(n_198),
.B1(n_200),
.B2(n_206),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_155),
.Y(n_181)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_182),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_106),
.B(n_50),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_183),
.B(n_187),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_184),
.A2(n_77),
.B1(n_140),
.B2(n_158),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_108),
.B(n_87),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_204),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_91),
.Y(n_187)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_189),
.Y(n_211)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_135),
.Y(n_191)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_191),
.Y(n_238)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

CKINVDCx12_ASAP7_75t_R g193 ( 
.A(n_123),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_132),
.B(n_88),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_195),
.B(n_196),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_92),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_109),
.A2(n_18),
.B1(n_98),
.B2(n_96),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_109),
.A2(n_18),
.B1(n_95),
.B2(n_82),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_203),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_116),
.B(n_80),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_149),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_208),
.Y(n_232)
);

HAxp5_ASAP7_75t_SL g206 ( 
.A(n_128),
.B(n_25),
.CON(n_206),
.SN(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_117),
.Y(n_207)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_128),
.B(n_147),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_141),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_103),
.Y(n_240)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_107),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_210),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_166),
.A2(n_58),
.B1(n_68),
.B2(n_60),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_212),
.A2(n_214),
.B1(n_221),
.B2(n_227),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_208),
.A2(n_148),
.B1(n_102),
.B2(n_158),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_164),
.A2(n_102),
.B1(n_148),
.B2(n_156),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_234),
.A2(n_239),
.B1(n_241),
.B2(n_103),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_172),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_243),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_184),
.A2(n_154),
.B1(n_107),
.B2(n_125),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_240),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_206),
.A2(n_156),
.B1(n_138),
.B2(n_130),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_176),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_187),
.B(n_175),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_246),
.A2(n_268),
.B(n_275),
.Y(n_282)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_249),
.A2(n_256),
.B1(n_259),
.B2(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_215),
.Y(n_250)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_215),
.Y(n_251)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_251),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_220),
.B(n_167),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_252),
.B(n_253),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_222),
.B(n_167),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_245),
.Y(n_254)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_254),
.Y(n_293)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_255),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_186),
.C(n_168),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_218),
.C(n_240),
.Y(n_283)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_260),
.B(n_261),
.Y(n_276)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_232),
.A2(n_170),
.B1(n_204),
.B2(n_138),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_262),
.A2(n_256),
.B1(n_251),
.B2(n_250),
.Y(n_300)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

AND2x6_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_233),
.Y(n_264)
);

AND2x6_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_243),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_216),
.B(n_191),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_265),
.B(n_266),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_209),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_220),
.B(n_192),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_267),
.B(n_269),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_226),
.A2(n_190),
.B(n_205),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_268),
.A2(n_242),
.B(n_224),
.Y(n_294)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_271),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_199),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_233),
.B(n_203),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_274),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_236),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_273),
.A2(n_232),
.B1(n_226),
.B2(n_241),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_277),
.A2(n_279),
.B1(n_287),
.B2(n_252),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_216),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_283),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_273),
.A2(n_214),
.B1(n_218),
.B2(n_221),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_282),
.A2(n_294),
.B(n_276),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_275),
.A2(n_246),
.B1(n_265),
.B2(n_253),
.Y(n_287)
);

AND2x6_ASAP7_75t_L g329 ( 
.A(n_288),
.B(n_248),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_258),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_291),
.Y(n_324)
);

OAI32xp33_ASAP7_75t_L g292 ( 
.A1(n_264),
.A2(n_228),
.A3(n_229),
.B1(n_212),
.B2(n_224),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_297),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_234),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_120),
.C(n_112),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_298),
.B(n_304),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_260),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_242),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_301),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_266),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_267),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_264),
.B(n_246),
.C(n_262),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_316),
.Y(n_341)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_276),
.Y(n_307)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_307),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_282),
.A2(n_249),
.B(n_272),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_308),
.Y(n_343)
);

NOR3xp33_ASAP7_75t_L g347 ( 
.A(n_309),
.B(n_325),
.C(n_327),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_299),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_310),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_311),
.B(n_313),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_261),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_290),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_314),
.B(n_317),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_315),
.A2(n_329),
.B1(n_330),
.B2(n_295),
.Y(n_351)
);

FAx1_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_270),
.CI(n_269),
.CON(n_316),
.SN(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_247),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_254),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_318),
.B(n_321),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_286),
.B(n_255),
.Y(n_319)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_254),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_320),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_254),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_259),
.Y(n_322)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_322),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_303),
.Y(n_325)
);

NAND2x1_ASAP7_75t_SL g327 ( 
.A(n_287),
.B(n_249),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_263),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_328),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_279),
.A2(n_231),
.B1(n_217),
.B2(n_237),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_284),
.Y(n_331)
);

NOR3xp33_ASAP7_75t_L g362 ( 
.A(n_331),
.B(n_335),
.C(n_336),
.Y(n_362)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_284),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_300),
.A2(n_231),
.B1(n_237),
.B2(n_217),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_333),
.A2(n_280),
.B1(n_277),
.B2(n_297),
.Y(n_339)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_285),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_293),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_285),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_294),
.A2(n_213),
.B(n_202),
.Y(n_336)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_337),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_339),
.A2(n_351),
.B1(n_356),
.B2(n_310),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_283),
.C(n_278),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_340),
.B(n_346),
.C(n_358),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_312),
.B(n_301),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_353),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_298),
.C(n_292),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_324),
.B(n_281),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_349),
.B(n_350),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_325),
.B(n_281),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_323),
.B(n_288),
.Y(n_353)
);

AO22x1_ASAP7_75t_SL g355 ( 
.A1(n_316),
.A2(n_288),
.B1(n_280),
.B2(n_289),
.Y(n_355)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_355),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_306),
.A2(n_289),
.B1(n_274),
.B2(n_217),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_317),
.Y(n_357)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_357),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_213),
.C(n_236),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_307),
.Y(n_359)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_359),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_211),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_365),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_326),
.B(n_236),
.C(n_146),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_364),
.B(n_336),
.C(n_320),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_326),
.B(n_211),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_348),
.B(n_363),
.Y(n_368)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_368),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_348),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_369),
.B(n_375),
.Y(n_402)
);

A2O1A1Ixp33_ASAP7_75t_SL g372 ( 
.A1(n_341),
.A2(n_305),
.B(n_329),
.C(n_327),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_372),
.A2(n_355),
.B(n_343),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_340),
.B(n_309),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_380),
.Y(n_399)
);

INVxp33_ASAP7_75t_SL g375 ( 
.A(n_344),
.Y(n_375)
);

XNOR2x2_ASAP7_75t_SL g376 ( 
.A(n_341),
.B(n_305),
.Y(n_376)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_376),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_339),
.A2(n_315),
.B1(n_314),
.B2(n_330),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_378),
.A2(n_383),
.B1(n_396),
.B2(n_352),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_366),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_379),
.B(n_388),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_345),
.B(n_315),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_360),
.Y(n_382)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_382),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_338),
.A2(n_329),
.B1(n_321),
.B2(n_318),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_360),
.Y(n_385)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_385),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_346),
.B(n_327),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_387),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_353),
.B(n_327),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_363),
.Y(n_388)
);

AOI21xp33_ASAP7_75t_L g389 ( 
.A1(n_342),
.A2(n_308),
.B(n_311),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_SL g424 ( 
.A(n_389),
.B(n_230),
.C(n_165),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_364),
.C(n_352),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_361),
.B(n_316),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_358),
.Y(n_405)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_359),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_394),
.B(n_395),
.Y(n_412)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_367),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_354),
.A2(n_322),
.B1(n_331),
.B2(n_335),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_397),
.B(n_219),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_398),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_400),
.A2(n_372),
.B(n_392),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_374),
.B(n_365),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_403),
.B(n_405),
.Y(n_432)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_390),
.Y(n_404)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_404),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_408),
.B(n_423),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_381),
.A2(n_343),
.B1(n_355),
.B2(n_316),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_409),
.A2(n_411),
.B1(n_417),
.B2(n_419),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_377),
.B(n_313),
.C(n_328),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_410),
.B(n_413),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_381),
.A2(n_319),
.B1(n_347),
.B2(n_356),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_368),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_377),
.B(n_320),
.C(n_334),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_415),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_380),
.B(n_320),
.C(n_332),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_382),
.A2(n_362),
.B1(n_333),
.B2(n_274),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_376),
.A2(n_237),
.B1(n_248),
.B2(n_207),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_370),
.B(n_386),
.C(n_387),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_421),
.B(n_173),
.Y(n_446)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_422),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_378),
.A2(n_122),
.B1(n_173),
.B2(n_201),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_424),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_383),
.A2(n_194),
.B1(n_219),
.B2(n_130),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_425),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_420),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_426),
.B(n_442),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_370),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_434),
.B(n_437),
.Y(n_463)
);

AOI322xp5_ASAP7_75t_L g435 ( 
.A1(n_418),
.A2(n_391),
.A3(n_371),
.B1(n_384),
.B2(n_372),
.C1(n_393),
.C2(n_390),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_435),
.B(n_447),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_421),
.B(n_373),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_402),
.Y(n_438)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_438),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_439),
.B(n_444),
.Y(n_453)
);

CKINVDCx14_ASAP7_75t_R g440 ( 
.A(n_412),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_440),
.A2(n_448),
.B1(n_409),
.B2(n_419),
.Y(n_460)
);

AOI322xp5_ASAP7_75t_SL g442 ( 
.A1(n_407),
.A2(n_372),
.A3(n_373),
.B1(n_230),
.B2(n_188),
.C1(n_197),
.C2(n_159),
.Y(n_442)
);

A2O1A1O1Ixp25_ASAP7_75t_L g443 ( 
.A1(n_406),
.A2(n_165),
.B(n_210),
.C(n_197),
.D(n_189),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_443),
.A2(n_423),
.B(n_400),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_410),
.B(n_159),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_404),
.Y(n_445)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_445),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_446),
.B(n_450),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_417),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_411),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_416),
.Y(n_449)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_449),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_408),
.B(n_188),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_401),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_452),
.B(n_454),
.Y(n_481)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_430),
.Y(n_455)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_451),
.B(n_415),
.C(n_399),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_457),
.B(n_464),
.Y(n_477)
);

AO21x1_ASAP7_75t_L g489 ( 
.A1(n_458),
.A2(n_157),
.B(n_131),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_460),
.A2(n_471),
.B(n_169),
.Y(n_490)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_445),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_434),
.B(n_399),
.C(n_405),
.Y(n_465)
);

NOR2xp67_ASAP7_75t_SL g486 ( 
.A(n_465),
.B(n_467),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_450),
.B(n_401),
.C(n_398),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_433),
.A2(n_431),
.B1(n_428),
.B2(n_436),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_468),
.A2(n_469),
.B1(n_470),
.B2(n_153),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_431),
.A2(n_425),
.B1(n_403),
.B2(n_117),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_428),
.A2(n_185),
.B1(n_188),
.B2(n_180),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_427),
.B(n_182),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_444),
.B(n_185),
.C(n_180),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_472),
.B(n_125),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_437),
.C(n_432),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_474),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_432),
.C(n_441),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_467),
.B(n_439),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_481),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_441),
.C(n_429),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_476),
.B(n_479),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_455),
.B(n_443),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_452),
.B(n_162),
.C(n_157),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_480),
.B(n_454),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_459),
.A2(n_152),
.B(n_162),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_482),
.A2(n_169),
.B(n_462),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_152),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_483),
.B(n_461),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_453),
.B(n_174),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_489),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_485),
.A2(n_490),
.B1(n_471),
.B2(n_472),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_487),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_456),
.B(n_131),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_488),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_493),
.B(n_498),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_497),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_473),
.B(n_474),
.Y(n_498)
);

OA21x2_ASAP7_75t_SL g499 ( 
.A1(n_477),
.A2(n_478),
.B(n_486),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_499),
.B(n_10),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_501),
.B(n_103),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_476),
.B(n_453),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_503),
.A2(n_489),
.B(n_484),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_475),
.B(n_97),
.C(n_113),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_504),
.B(n_505),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_481),
.A2(n_48),
.B1(n_94),
.B2(n_126),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_508),
.B(n_509),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_492),
.B(n_480),
.C(n_137),
.Y(n_509)
);

NAND3xp33_ASAP7_75t_L g510 ( 
.A(n_495),
.B(n_12),
.C(n_8),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_510),
.A2(n_517),
.B(n_518),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_SL g511 ( 
.A1(n_491),
.A2(n_136),
.B1(n_126),
.B2(n_115),
.Y(n_511)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_511),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_500),
.A2(n_124),
.B(n_150),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_512),
.A2(n_513),
.B(n_515),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_495),
.A2(n_124),
.B(n_150),
.Y(n_513)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_516),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_503),
.B(n_9),
.Y(n_517)
);

OAI221xp5_ASAP7_75t_L g518 ( 
.A1(n_494),
.A2(n_115),
.B1(n_25),
.B2(n_32),
.C(n_31),
.Y(n_518)
);

OAI21xp33_ASAP7_75t_SL g519 ( 
.A1(n_507),
.A2(n_502),
.B(n_496),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_519),
.A2(n_2),
.B(n_3),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_506),
.A2(n_502),
.B1(n_25),
.B2(n_31),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_521),
.B(n_523),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_31),
.C(n_32),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_514),
.A2(n_7),
.B(n_14),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_526),
.A2(n_528),
.B(n_2),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_506),
.A2(n_32),
.B(n_28),
.Y(n_528)
);

AOI322xp5_ASAP7_75t_L g529 ( 
.A1(n_520),
.A2(n_32),
.A3(n_28),
.B1(n_8),
.B2(n_9),
.C1(n_14),
.C2(n_11),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_529),
.B(n_530),
.Y(n_538)
);

AOI322xp5_ASAP7_75t_L g530 ( 
.A1(n_524),
.A2(n_28),
.A3(n_14),
.B1(n_11),
.B2(n_9),
.C1(n_8),
.C2(n_1),
.Y(n_530)
);

AOI322xp5_ASAP7_75t_L g532 ( 
.A1(n_519),
.A2(n_28),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_2),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_532),
.B(n_525),
.C(n_531),
.Y(n_536)
);

AOI21x1_ASAP7_75t_L g535 ( 
.A1(n_533),
.A2(n_534),
.B(n_522),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_535),
.A2(n_536),
.B(n_537),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_534),
.B(n_527),
.C(n_28),
.Y(n_537)
);

BUFx24_ASAP7_75t_SL g540 ( 
.A(n_538),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_540),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_541)
);

AOI211xp5_ASAP7_75t_L g542 ( 
.A1(n_541),
.A2(n_539),
.B(n_4),
.C(n_6),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_542),
.B(n_3),
.Y(n_543)
);


endmodule