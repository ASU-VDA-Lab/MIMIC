module fake_jpeg_20461_n_100 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_100);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_31),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_48),
.B(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_0),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_53),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_39),
.B1(n_35),
.B2(n_38),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_55),
.A2(n_44),
.B1(n_36),
.B2(n_2),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_37),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_59),
.B1(n_0),
.B2(n_1),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx12_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_67),
.B1(n_70),
.B2(n_5),
.Y(n_78)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_58),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_66),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_13),
.C(n_29),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_57),
.B1(n_59),
.B2(n_2),
.Y(n_70)
);

AO21x1_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_3),
.B(n_4),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_3),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_80),
.B(n_10),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_78),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_82)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_82),
.Y(n_89)
);

AOI221xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_86),
.B1(n_30),
.B2(n_12),
.C(n_14),
.Y(n_87)
);

AO22x2_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_75),
.B1(n_79),
.B2(n_72),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_87),
.A2(n_85),
.B1(n_86),
.B2(n_17),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_89),
.Y(n_92)
);

AO21x1_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_90),
.B(n_15),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_11),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_19),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_20),
.B(n_22),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_96),
.A2(n_23),
.B(n_25),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_27),
.Y(n_100)
);


endmodule