module fake_jpeg_20067_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVxp67_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_6),
.B(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g15 ( 
.A(n_9),
.B(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_15),
.B(n_17),
.Y(n_22)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_18),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_1),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_19),
.B(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_19),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_10),
.B(n_12),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_10),
.B(n_8),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_21),
.A2(n_25),
.B(n_20),
.C(n_14),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_22),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_31),
.B(n_32),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_13),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

XNOR2x1_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_28),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_40),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_35),
.B(n_37),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_26),
.C(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_3),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_44),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_49),
.B(n_48),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);


endmodule