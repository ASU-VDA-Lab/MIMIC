module fake_jpeg_17106_n_168 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_23),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_9),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_8),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_0),
.Y(n_67)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_19),
.B1(n_42),
.B2(n_40),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_52),
.B1(n_63),
.B2(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_73),
.Y(n_75)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_59),
.B1(n_62),
.B2(n_50),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_92),
.B1(n_56),
.B2(n_45),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_65),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_78),
.B(n_85),
.Y(n_111)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_80),
.Y(n_118)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_51),
.B1(n_1),
.B2(n_2),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_44),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_49),
.B1(n_66),
.B2(n_58),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_114)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_69),
.A2(n_55),
.B1(n_64),
.B2(n_46),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_85),
.A2(n_66),
.B1(n_53),
.B2(n_58),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_101),
.B1(n_104),
.B2(n_105),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_98),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_102),
.B(n_113),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_61),
.B1(n_48),
.B2(n_51),
.Y(n_104)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_75),
.A2(n_60),
.B1(n_57),
.B2(n_3),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_110),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_116),
.B1(n_5),
.B2(n_7),
.Y(n_124)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_130),
.Y(n_137)
);

OR2x2_ASAP7_75t_SL g130 ( 
.A(n_111),
.B(n_7),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_125),
.A2(n_118),
.B(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_125),
.Y(n_142)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_134),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_103),
.C(n_94),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_135),
.B(n_136),
.Y(n_138)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_133),
.A2(n_105),
.B1(n_126),
.B2(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_95),
.Y(n_147)
);

AOI32xp33_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_137),
.A3(n_123),
.B1(n_124),
.B2(n_135),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_SL g151 ( 
.A1(n_143),
.A2(n_147),
.B(n_112),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_134),
.Y(n_145)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_146),
.B(n_147),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_144),
.A2(n_138),
.B(n_114),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_149),
.B(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_121),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_153),
.C(n_150),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_155),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_148),
.C(n_139),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_30),
.B1(n_38),
.B2(n_37),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_120),
.B1(n_109),
.B2(n_96),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_107),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_100),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_24),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_26),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_22),
.B(n_43),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_121),
.C(n_17),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_165),
.A2(n_16),
.B(n_35),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_15),
.C(n_34),
.Y(n_167)
);

FAx1_ASAP7_75t_SL g168 ( 
.A(n_167),
.B(n_13),
.CI(n_31),
.CON(n_168),
.SN(n_168)
);


endmodule