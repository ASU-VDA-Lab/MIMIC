module fake_jpeg_21676_n_124 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_124);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_24),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_64),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_0),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_0),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_1),
.Y(n_67)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_77),
.Y(n_86)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_42),
.B1(n_56),
.B2(n_55),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_57),
.B1(n_43),
.B2(n_48),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_88),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_38),
.B1(n_55),
.B2(n_39),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_87),
.B1(n_51),
.B2(n_47),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_38),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_83),
.B1(n_85),
.B2(n_2),
.Y(n_103)
);

OR2x2_ASAP7_75t_SL g83 ( 
.A(n_73),
.B(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_39),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_70),
.B(n_50),
.Y(n_88)
);

BUFx12f_ASAP7_75t_SL g89 ( 
.A(n_73),
.Y(n_89)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

BUFx24_ASAP7_75t_SL g92 ( 
.A(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_101),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_41),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_7),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_46),
.B1(n_40),
.B2(n_54),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_103),
.B(n_8),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_84),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_6),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_109),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_93),
.C(n_96),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_107),
.Y(n_115)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_113),
.B(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_111),
.B(n_115),
.Y(n_117)
);

OAI31xp33_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_108),
.A3(n_102),
.B(n_14),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_11),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_12),
.C(n_15),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_120),
.A2(n_17),
.B(n_18),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_94),
.B(n_23),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);


endmodule