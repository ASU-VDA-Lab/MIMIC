module real_jpeg_4271_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_1),
.B(n_73),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_1),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_1),
.B(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_1),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_1),
.B(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_1),
.B(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_2),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_2),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_2),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_2),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_2),
.B(n_133),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_2),
.B(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_2),
.B(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_3),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_3),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_3),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_3),
.B(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_3),
.B(n_418),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_4),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_4),
.Y(n_174)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_4),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g136 ( 
.A(n_5),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_5),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_5),
.B(n_224),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_5),
.B(n_241),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_5),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_5),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_5),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_5),
.B(n_409),
.Y(n_408)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_6),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_6),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_6),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_6),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_6),
.B(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_6),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_6),
.B(n_185),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_6),
.B(n_197),
.Y(n_196)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_8),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_8),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_9),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_9),
.B(n_41),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_9),
.B(n_81),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_9),
.B(n_170),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_9),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_9),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_9),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_9),
.B(n_342),
.Y(n_341)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_10),
.Y(n_144)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_10),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_11),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_11),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_11),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_11),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_11),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_11),
.B(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_11),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_11),
.B(n_266),
.Y(n_265)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_13),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_13),
.Y(n_137)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_13),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_13),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_14),
.Y(n_135)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_14),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_14),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_15),
.Y(n_25)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_15),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_15),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_15),
.B(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_15),
.B(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_156),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_155),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_92),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_20),
.B(n_92),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_75),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_42),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.C(n_39),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_23),
.B(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_31),
.C(n_33),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_46),
.C(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_24),
.A2(n_46),
.B1(n_47),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_24),
.A2(n_91),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_24),
.A2(n_91),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_24),
.B(n_166),
.C(n_169),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

OR2x2_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_35),
.Y(n_34)
);

OR2x2_ASAP7_75t_SL g47 ( 
.A(n_25),
.B(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_25),
.B(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_29),
.Y(n_109)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_29),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_29),
.Y(n_386)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_30),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_30),
.Y(n_287)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_30),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_31),
.A2(n_33),
.B1(n_34),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_31),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_33),
.A2(n_34),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_33),
.A2(n_34),
.B1(n_179),
.B2(n_298),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_34),
.B(n_99),
.C(n_102),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_34),
.B(n_176),
.C(n_179),
.Y(n_175)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_36),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_37),
.A2(n_39),
.B1(n_40),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_37),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_64),
.B1(n_65),
.B2(n_74),
.Y(n_42)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_59),
.B2(n_63),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_52),
.B2(n_58),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_46),
.A2(n_47),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_47),
.B(n_195),
.C(n_199),
.Y(n_288)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_48),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_50),
.Y(n_311)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_51),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_52),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_52),
.B(n_264),
.Y(n_263)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_56),
.Y(n_167)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_57),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_57),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_58),
.B(n_265),
.C(n_268),
.Y(n_325)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_59),
.A2(n_63),
.B1(n_111),
.B2(n_120),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_59),
.B(n_112),
.C(n_119),
.Y(n_151)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_71),
.B2(n_72),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_69),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_99),
.C(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_68),
.A2(n_69),
.B1(n_107),
.B2(n_108),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.C(n_88),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_76),
.B(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_79),
.B(n_88),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.C(n_87),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_80),
.A2(n_83),
.B1(n_84),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_83),
.A2(n_84),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_84),
.B(n_127),
.C(n_184),
.Y(n_346)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_85),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_86),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_145),
.C(n_153),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_93),
.B(n_485),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_121),
.C(n_124),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_94),
.B(n_479),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_106),
.C(n_110),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_95),
.B(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_105),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_98),
.A2(n_99),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_99),
.B(n_196),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_99),
.B(n_196),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx8_ASAP7_75t_L g376 ( 
.A(n_101),
.Y(n_376)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_106),
.B(n_110),
.Y(n_355)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_115),
.B1(n_118),
.B2(n_119),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_115),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_115),
.B(n_248),
.C(n_255),
.Y(n_262)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_121),
.B(n_124),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_138),
.C(n_140),
.Y(n_124)
);

AO22x1_ASAP7_75t_SL g362 ( 
.A1(n_125),
.A2(n_126),
.B1(n_363),
.B2(n_364),
.Y(n_362)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.C(n_136),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_127),
.A2(n_184),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_127),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_127),
.A2(n_136),
.B1(n_273),
.B2(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_127),
.B(n_373),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_127),
.A2(n_273),
.B1(n_373),
.B2(n_374),
.Y(n_411)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_129),
.Y(n_238)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_129),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_129),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_130),
.A2(n_223),
.B1(n_227),
.B2(n_228),
.Y(n_222)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_130),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_130),
.B(n_219),
.C(n_223),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_130),
.A2(n_227),
.B1(n_330),
.B2(n_332),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_135),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_135),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_136),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_140),
.A2(n_141),
.B1(n_340),
.B2(n_341),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_141),
.B(n_341),
.C(n_346),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_142),
.Y(n_216)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_143),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_145),
.B(n_153),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_151),
.C(n_152),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_146),
.A2(n_147),
.B1(n_481),
.B2(n_482),
.Y(n_480)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_151),
.B(n_152),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_475),
.B(n_489),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_365),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_319),
.B(n_348),
.C(n_349),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_289),
.B(n_318),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_160),
.B(n_473),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_257),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_161),
.B(n_257),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_217),
.C(n_244),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_162),
.B(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_191),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_163),
.B(n_192),
.C(n_200),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_175),
.C(n_182),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_164),
.B(n_314),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_173),
.B(n_220),
.Y(n_433)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_175),
.A2(n_182),
.B1(n_183),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_175),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_176),
.B(n_297),
.Y(n_296)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_179),
.Y(n_298)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_184),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_184),
.A2(n_187),
.B1(n_188),
.B2(n_274),
.Y(n_312)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_200),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_197),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_208),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_202),
.B(n_204),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_201),
.B(n_209),
.C(n_214),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_214),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_215),
.B(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_217),
.B(n_244),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_229),
.C(n_231),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_218),
.A2(n_229),
.B1(n_230),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_218),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_220),
.B(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_223),
.Y(n_228)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_231),
.B(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.C(n_239),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_232),
.A2(n_233),
.B1(n_462),
.B2(n_463),
.Y(n_461)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_234),
.A2(n_235),
.B1(n_239),
.B2(n_240),
.Y(n_463)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_256),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_247),
.C(n_256),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_254),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_253),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_253),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_258),
.B(n_260),
.C(n_275),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_275),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_270),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_262),
.B(n_263),
.C(n_270),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_276),
.B(n_278),
.C(n_279),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_288),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_281),
.B(n_283),
.C(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_288),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_316),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_290),
.B(n_316),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_295),
.C(n_313),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_291),
.A2(n_292),
.B1(n_467),
.B2(n_468),
.Y(n_466)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_295),
.B(n_313),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_299),
.C(n_312),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_296),
.B(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_299),
.B(n_312),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_305),
.C(n_308),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_300),
.A2(n_301),
.B1(n_308),
.B2(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_305),
.B(n_393),
.Y(n_392)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_307),
.Y(n_418)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_308),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_309),
.B(n_385),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_309),
.B(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_320),
.B(n_350),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_321),
.B(n_322),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_322),
.B(n_351),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_322),
.B(n_351),
.Y(n_474)
);

FAx1_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_333),
.CI(n_347),
.CON(n_322),
.SN(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_329),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_326),
.C(n_329),
.Y(n_358)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_330),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_336),
.C(n_338),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_338),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_346),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx8_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_352),
.B(n_354),
.C(n_356),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_356),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_359),
.B2(n_360),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_357),
.B(n_361),
.C(n_362),
.Y(n_483)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

OAI31xp33_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_471),
.A3(n_472),
.B(n_474),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_465),
.B(n_470),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_452),
.B(n_464),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_412),
.B(n_451),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_370),
.B(n_395),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_370),
.B(n_395),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_382),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_371),
.B(n_383),
.C(n_392),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_377),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_372),
.B(n_378),
.C(n_381),
.Y(n_460)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.Y(n_377)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_392),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_387),
.C(n_390),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_384),
.B(n_397),
.Y(n_396)
);

INVx11_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_387),
.A2(n_388),
.B1(n_390),
.B2(n_391),
.Y(n_397)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_398),
.C(n_411),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_396),
.B(n_448),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_398),
.A2(n_399),
.B1(n_411),
.B2(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_407),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_400),
.A2(n_401),
.B1(n_407),
.B2(n_408),
.Y(n_421)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_411),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_445),
.B(n_450),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_431),
.B(n_444),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_422),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_422),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_421),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_419),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_417),
.B(n_419),
.C(n_421),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_428),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_423),
.A2(n_424),
.B1(n_428),
.B2(n_429),
.Y(n_442)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_429),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_438),
.B(n_443),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx8_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_442),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_439),
.B(n_442),
.Y(n_443)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_446),
.B(n_447),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_453),
.B(n_454),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_455),
.A2(n_456),
.B1(n_458),
.B2(n_459),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_460),
.C(n_461),
.Y(n_469)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_461),
.Y(n_459)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_466),
.B(n_469),
.Y(n_470)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_467),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_486),
.Y(n_475)
);

OAI21xp33_ASAP7_75t_L g489 ( 
.A1(n_476),
.A2(n_490),
.B(n_491),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_484),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_484),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_480),
.C(n_483),
.Y(n_477)
);

FAx1_ASAP7_75t_SL g488 ( 
.A(n_478),
.B(n_480),
.CI(n_483),
.CON(n_488),
.SN(n_488)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_487),
.B(n_488),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g493 ( 
.A(n_488),
.Y(n_493)
);


endmodule