module fake_jpeg_10287_n_284 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_284);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_18),
.Y(n_51)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NAND2xp33_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_26),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_41),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_26),
.B1(n_23),
.B2(n_19),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_39),
.A2(n_33),
.B1(n_37),
.B2(n_20),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_36),
.B1(n_37),
.B2(n_33),
.Y(n_69)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_51),
.A2(n_35),
.B(n_36),
.C(n_23),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_35),
.B(n_29),
.Y(n_81)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_26),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_62),
.Y(n_84)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_23),
.B1(n_24),
.B2(n_15),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_37),
.B1(n_49),
.B2(n_36),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_23),
.B1(n_37),
.B2(n_33),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_28),
.B1(n_31),
.B2(n_53),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_34),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_70),
.Y(n_85)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx4f_ASAP7_75t_SL g96 ( 
.A(n_68),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_18),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_34),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_53),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_47),
.B1(n_24),
.B2(n_54),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_81),
.B1(n_91),
.B2(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_83),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_87),
.B(n_71),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_55),
.B1(n_50),
.B2(n_47),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_98),
.B1(n_57),
.B2(n_68),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_61),
.Y(n_89)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_58),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_53),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_83),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_27),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_63),
.A2(n_31),
.B1(n_28),
.B2(n_54),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_60),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_104),
.C(n_112),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_56),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_109),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_101),
.A2(n_110),
.B1(n_95),
.B2(n_59),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_56),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_105),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

FAx1_ASAP7_75t_SL g108 ( 
.A(n_85),
.B(n_73),
.CI(n_57),
.CON(n_108),
.SN(n_108)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_117),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_71),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_65),
.B1(n_66),
.B2(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_67),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_109),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_24),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_82),
.C(n_97),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_115),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_74),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_88),
.B(n_74),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_80),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_80),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_120),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_114),
.A2(n_68),
.B1(n_89),
.B2(n_82),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_121),
.A2(n_32),
.B(n_15),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_133),
.Y(n_147)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_128),
.B(n_129),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_108),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_17),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_96),
.B1(n_21),
.B2(n_22),
.Y(n_160)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_88),
.Y(n_134)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_138),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_88),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_137),
.A2(n_139),
.B1(n_43),
.B2(n_31),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_95),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_59),
.B1(n_93),
.B2(n_58),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_27),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_99),
.B(n_83),
.Y(n_142)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_102),
.Y(n_143)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_138),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_146),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_108),
.B1(n_116),
.B2(n_112),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_145),
.A2(n_148),
.B1(n_150),
.B2(n_156),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_116),
.B1(n_114),
.B2(n_119),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_166),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_93),
.B1(n_58),
.B2(n_43),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_153),
.Y(n_187)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_96),
.B1(n_28),
.B2(n_90),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_158),
.B(n_132),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_159),
.A2(n_167),
.B(n_168),
.Y(n_190)
);

XNOR2x1_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_167),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_136),
.A2(n_96),
.B1(n_20),
.B2(n_22),
.Y(n_162)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_134),
.A2(n_20),
.B1(n_15),
.B2(n_22),
.Y(n_164)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_122),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_133),
.A2(n_16),
.B1(n_27),
.B2(n_13),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_169),
.A2(n_168),
.B1(n_140),
.B2(n_16),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_147),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_176),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_126),
.C(n_143),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_184),
.C(n_191),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_162),
.B1(n_164),
.B2(n_154),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_147),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_152),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_177),
.B(n_150),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_151),
.Y(n_183)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_126),
.C(n_123),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_131),
.Y(n_185)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_142),
.Y(n_186)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_189),
.B(n_144),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_152),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_145),
.B(n_123),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_163),
.C(n_161),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_195),
.C(n_204),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_161),
.C(n_157),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_157),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_171),
.B(n_190),
.Y(n_221)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_201),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_203),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_186),
.B(n_127),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_148),
.C(n_156),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_141),
.C(n_128),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_170),
.C(n_176),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_208),
.B(n_209),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_185),
.B(n_32),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_8),
.C(n_12),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_9),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_182),
.B1(n_189),
.B2(n_171),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_212),
.A2(n_222),
.B1(n_179),
.B2(n_190),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_173),
.B(n_183),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_193),
.B(n_180),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_205),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_219),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_178),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_209),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_225),
.C(n_227),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_181),
.C(n_182),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_188),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_214),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_180),
.C(n_178),
.Y(n_227)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_211),
.A2(n_204),
.B1(n_179),
.B2(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_236),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_241),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_195),
.B1(n_27),
.B2(n_13),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_232),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_13),
.B1(n_7),
.B2(n_12),
.Y(n_233)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_212),
.A2(n_215),
.B1(n_225),
.B2(n_224),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_237),
.B1(n_9),
.B2(n_8),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_32),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_227),
.A2(n_13),
.B1(n_7),
.B2(n_12),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_5),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_5),
.C(n_11),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_214),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_21),
.Y(n_247)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_248),
.C(n_253),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_252),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_0),
.C(n_1),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_0),
.C(n_1),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_231),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_254),
.A2(n_235),
.B(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_239),
.Y(n_255)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_259),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_244),
.A2(n_240),
.B(n_236),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_262),
.C(n_246),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_230),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_263),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_249),
.A2(n_6),
.B(n_8),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_6),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_264),
.B(n_245),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_265),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_269),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_259),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_254),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_257),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_261),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_267),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_276),
.A2(n_273),
.B(n_268),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_272),
.B(n_270),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_279),
.A2(n_277),
.B(n_250),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_280),
.A2(n_250),
.B(n_6),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_0),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_3),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_3),
.B(n_4),
.Y(n_284)
);


endmodule