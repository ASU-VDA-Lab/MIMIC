module fake_jpeg_10087_n_147 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_147);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx5p33_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx24_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_22),
.A2(n_25),
.B1(n_18),
.B2(n_20),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_5),
.Y(n_26)
);

OR2x2_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx2_ASAP7_75t_R g29 ( 
.A(n_27),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_26),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_18),
.B1(n_17),
.B2(n_10),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_14),
.B1(n_28),
.B2(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_38),
.B(n_45),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_25),
.B1(n_31),
.B2(n_23),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_13),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_32),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_27),
.B(n_24),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_35),
.B1(n_37),
.B2(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_9),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_32),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_54),
.B1(n_56),
.B2(n_59),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_25),
.B1(n_31),
.B2(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_49),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_31),
.B1(n_21),
.B2(n_12),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_11),
.B1(n_12),
.B2(n_2),
.Y(n_62)
);

OR2x4_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_45),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_65),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_66),
.B(n_70),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_9),
.B(n_1),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_43),
.C(n_39),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_73),
.C(n_79),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_74),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_43),
.Y(n_79)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_52),
.B(n_63),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_85),
.B(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_79),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_62),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_82),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_32),
.C(n_50),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_67),
.C(n_72),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_46),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_32),
.B(n_34),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_95),
.A2(n_96),
.B1(n_33),
.B2(n_23),
.Y(n_106)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_98),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_89),
.C(n_81),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_72),
.B1(n_66),
.B2(n_32),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_108),
.B1(n_84),
.B2(n_91),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_90),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_104),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_106),
.B1(n_95),
.B2(n_88),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_21),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_97),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_33),
.B1(n_0),
.B2(n_3),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_118),
.C(n_98),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_114),
.B(n_116),
.Y(n_119)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_113),
.B(n_117),
.Y(n_121)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_33),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_104),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_33),
.Y(n_130)
);

BUFx24_ASAP7_75t_SL g123 ( 
.A(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_92),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_107),
.C(n_105),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_85),
.C(n_33),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_87),
.B1(n_102),
.B2(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

BUFx24_ASAP7_75t_SL g133 ( 
.A(n_127),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_129),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_131),
.B(n_132),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_2),
.Y(n_131)
);

AOI21x1_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_3),
.B(n_5),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_130),
.A2(n_121),
.B(n_6),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_8),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_128),
.C(n_6),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_141),
.B(n_8),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_139),
.B(n_140),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_133),
.B(n_6),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_135),
.C(n_8),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_143),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_144),
.Y(n_147)
);


endmodule