module fake_jpeg_29596_n_44 (n_3, n_2, n_1, n_0, n_4, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_2),
.B(n_3),
.Y(n_6)
);

BUFx2_ASAP7_75t_R g7 ( 
.A(n_5),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_4),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_19),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_15),
.B(n_20),
.Y(n_26)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_12),
.Y(n_21)
);

MAJx2_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_7),
.C(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_19),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_20),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_32),
.B1(n_9),
.B2(n_11),
.Y(n_34)
);

OAI32xp33_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_27),
.A3(n_15),
.B1(n_21),
.B2(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_22),
.B1(n_12),
.B2(n_23),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_17),
.B(n_12),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_16),
.C(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_9),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_23),
.C(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_36),
.C(n_33),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_40),
.B(n_39),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_38),
.B(n_31),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_3),
.Y(n_44)
);


endmodule