module fake_jpeg_7964_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_14),
.A2(n_0),
.B(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_11),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_13),
.C(n_8),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_14),
.B1(n_12),
.B2(n_7),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_14),
.B1(n_7),
.B2(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_24),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_34),
.A2(n_9),
.B1(n_8),
.B2(n_7),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_26),
.B1(n_24),
.B2(n_21),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_32),
.C(n_40),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_39),
.B1(n_36),
.B2(n_15),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_26),
.B1(n_21),
.B2(n_9),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_43),
.B1(n_44),
.B2(n_6),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_4),
.Y(n_43)
);

XOR2x2_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_23),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_41),
.Y(n_47)
);

OAI31xp33_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_48),
.A3(n_6),
.B(n_0),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_45),
.C(n_17),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_50),
.Y(n_51)
);


endmodule