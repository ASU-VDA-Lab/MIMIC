module fake_jpeg_847_n_292 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_292);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_292;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_40),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_20),
.B(n_39),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_50),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_23),
.B1(n_34),
.B2(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_46),
.Y(n_99)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_0),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_30),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_16),
.B(n_15),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_22),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_16),
.B(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_57),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_14),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_58),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_6),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_65),
.A2(n_81),
.B1(n_82),
.B2(n_101),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_30),
.B1(n_26),
.B2(n_25),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_70),
.A2(n_59),
.B1(n_38),
.B2(n_8),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_72),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_23),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_34),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_74),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_29),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_75),
.B(n_80),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_28),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_88),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_17),
.B1(n_37),
.B2(n_45),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_41),
.A2(n_37),
.B1(n_39),
.B2(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_20),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_28),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_19),
.B(n_27),
.C(n_21),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_89),
.B(n_95),
.Y(n_111)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_27),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_94),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_30),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_26),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_37),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_6),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_100),
.B(n_93),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_52),
.A2(n_36),
.B1(n_38),
.B2(n_8),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_55),
.A2(n_36),
.B1(n_38),
.B2(n_8),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_38),
.B1(n_7),
.B2(n_9),
.Y(n_119)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_109),
.A2(n_84),
.B1(n_99),
.B2(n_96),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_80),
.A2(n_67),
.B(n_66),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_114),
.A2(n_131),
.B(n_116),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_89),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_137),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_134),
.B1(n_138),
.B2(n_140),
.Y(n_156)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_6),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_135),
.Y(n_143)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_124),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_103),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_128),
.Y(n_147)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_131),
.Y(n_144)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_128),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_82),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_14),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_64),
.B(n_68),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_84),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_93),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_79),
.A2(n_106),
.B1(n_76),
.B2(n_105),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_137),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_79),
.A2(n_106),
.B1(n_76),
.B2(n_105),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_68),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_142),
.B(n_163),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_SL g192 ( 
.A(n_149),
.B(n_143),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_113),
.A2(n_83),
.B1(n_96),
.B2(n_90),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_152),
.B1(n_166),
.B2(n_156),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_90),
.B(n_86),
.C(n_83),
.Y(n_155)
);

OA21x2_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_168),
.B(n_166),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_86),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_160),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_109),
.A2(n_119),
.B1(n_129),
.B2(n_122),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_162),
.B1(n_161),
.B2(n_152),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_159),
.B(n_146),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_129),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_141),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_114),
.B(n_126),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_117),
.B(n_118),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_133),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_175),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_130),
.A2(n_120),
.B1(n_116),
.B2(n_132),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_107),
.B(n_110),
.C(n_132),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_172),
.C(n_170),
.Y(n_178)
);

NOR2x1p5_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_110),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_170),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_128),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_171),
.B(n_154),
.Y(n_196)
);

AOI22x1_ASAP7_75t_SL g174 ( 
.A1(n_108),
.A2(n_115),
.B1(n_111),
.B2(n_113),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_174),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_123),
.B(n_137),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_181),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_204),
.Y(n_214)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_144),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_185),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_144),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_144),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_186),
.Y(n_227)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_157),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_193),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_142),
.A2(n_172),
.B(n_149),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_190),
.A2(n_179),
.B(n_184),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_173),
.C(n_189),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_158),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_194),
.A2(n_202),
.B1(n_164),
.B2(n_168),
.Y(n_206)
);

O2A1O1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_174),
.A2(n_155),
.B(n_168),
.C(n_148),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_178),
.B(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_170),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_197),
.B(n_199),
.Y(n_211)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_145),
.Y(n_198)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_167),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_200),
.B(n_205),
.Y(n_210)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_148),
.A2(n_164),
.B1(n_151),
.B2(n_147),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_173),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_213),
.B1(n_217),
.B2(n_197),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_190),
.A2(n_147),
.B(n_171),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_208),
.A2(n_191),
.B(n_185),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_204),
.Y(n_242)
);

NAND3xp33_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_191),
.C(n_176),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_199),
.B1(n_193),
.B2(n_181),
.Y(n_213)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_195),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_179),
.A2(n_204),
.B1(n_195),
.B2(n_177),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_180),
.B(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_224),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_221),
.A2(n_223),
.B(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_186),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_192),
.C(n_188),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_233),
.C(n_241),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_239),
.B1(n_224),
.B2(n_216),
.Y(n_248)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_209),
.C(n_221),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

FAx1_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_216),
.CI(n_217),
.CON(n_237),
.SN(n_237)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_204),
.B1(n_182),
.B2(n_187),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_243),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_198),
.C(n_203),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_244),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_213),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_220),
.B(n_210),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_247),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_227),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

AOI321xp33_ASAP7_75t_L g252 ( 
.A1(n_237),
.A2(n_208),
.A3(n_222),
.B1(n_207),
.B2(n_212),
.C(n_225),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_240),
.B(n_238),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_206),
.B1(n_212),
.B2(n_225),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_257),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_235),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_259),
.B(n_233),
.C(n_230),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_254),
.C(n_248),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_259),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_265),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_270),
.B(n_254),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_245),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_244),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_234),
.Y(n_270)
);

OAI21xp33_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_252),
.B(n_255),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_263),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_274),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g274 ( 
.A(n_261),
.B(n_253),
.CI(n_258),
.CON(n_274),
.SN(n_274)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_275),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_262),
.B(n_226),
.CI(n_228),
.CON(n_278),
.SN(n_278)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_278),
.A2(n_269),
.B1(n_250),
.B2(n_228),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_280),
.B(n_282),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_266),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_283),
.B(n_271),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_280),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_279),
.B(n_277),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_285),
.A2(n_282),
.B(n_281),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_288),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_289),
.Y(n_290)
);

OA21x2_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_286),
.B(n_271),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_283),
.Y(n_292)
);


endmodule