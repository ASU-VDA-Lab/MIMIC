module real_aes_6185_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
OAI22xp5_ASAP7_75t_SL g519 ( .A1(n_0), .A2(n_14), .B1(n_520), .B2(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_0), .Y(n_520) );
INVx1_ASAP7_75t_L g320 ( .A(n_1), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_2), .A2(n_47), .B1(n_170), .B2(n_173), .Y(n_169) );
AOI21xp33_ASAP7_75t_L g227 ( .A1(n_3), .A2(n_228), .B(n_229), .Y(n_227) );
INVx1_ASAP7_75t_L g185 ( .A(n_4), .Y(n_185) );
AND2x6_ASAP7_75t_L g202 ( .A(n_4), .B(n_183), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_4), .B(n_535), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_5), .A2(n_296), .B(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g236 ( .A(n_6), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_7), .B(n_288), .Y(n_287) );
AO22x2_ASAP7_75t_L g90 ( .A1(n_8), .A2(n_25), .B1(n_91), .B2(n_92), .Y(n_90) );
INVx1_ASAP7_75t_L g199 ( .A(n_9), .Y(n_199) );
INVx1_ASAP7_75t_L g302 ( .A(n_10), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_11), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_12), .B(n_247), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_12), .A2(n_518), .B1(n_519), .B2(n_522), .Y(n_517) );
INVx1_ASAP7_75t_L g522 ( .A(n_12), .Y(n_522) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_13), .A2(n_26), .B1(n_91), .B2(n_96), .Y(n_95) );
INVx1_ASAP7_75t_L g521 ( .A(n_14), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_15), .B(n_228), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_16), .B(n_224), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g299 ( .A1(n_17), .A2(n_300), .B(n_301), .C(n_303), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g107 ( .A1(n_18), .A2(n_33), .B1(n_108), .B2(n_115), .Y(n_107) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_19), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_20), .B(n_234), .Y(n_321) );
INVx1_ASAP7_75t_L g212 ( .A(n_21), .Y(n_212) );
AOI22xp33_ASAP7_75t_SL g148 ( .A1(n_22), .A2(n_45), .B1(n_149), .B2(n_156), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g83 ( .A1(n_23), .A2(n_63), .B1(n_84), .B2(n_101), .Y(n_83) );
INVx2_ASAP7_75t_L g206 ( .A(n_24), .Y(n_206) );
OAI221xp5_ASAP7_75t_L g527 ( .A1(n_26), .A2(n_41), .B1(n_51), .B2(n_528), .C(n_529), .Y(n_527) );
INVxp67_ASAP7_75t_L g530 ( .A(n_26), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_27), .A2(n_202), .B(n_213), .C(n_258), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_28), .Y(n_120) );
INVx1_ASAP7_75t_L g210 ( .A(n_29), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_29), .A2(n_509), .B1(n_524), .B2(n_532), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_30), .B(n_234), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_31), .B(n_165), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_32), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_34), .B(n_162), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_35), .Y(n_129) );
CKINVDCx16_ASAP7_75t_R g216 ( .A(n_36), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_37), .B(n_228), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_38), .A2(n_204), .B1(n_207), .B2(n_213), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_39), .Y(n_267) );
CKINVDCx16_ASAP7_75t_R g317 ( .A(n_40), .Y(n_317) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_41), .A2(n_59), .B1(n_91), .B2(n_96), .Y(n_100) );
INVxp67_ASAP7_75t_L g531 ( .A(n_41), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_42), .A2(n_233), .B(n_235), .C(n_238), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g277 ( .A(n_43), .Y(n_277) );
INVx1_ASAP7_75t_L g230 ( .A(n_44), .Y(n_230) );
INVx1_ASAP7_75t_L g183 ( .A(n_46), .Y(n_183) );
INVx1_ASAP7_75t_L g198 ( .A(n_48), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_49), .Y(n_528) );
AOI22xp5_ASAP7_75t_SL g79 ( .A1(n_50), .A2(n_80), .B1(n_176), .B2(n_177), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_50), .Y(n_177) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_51), .A2(n_66), .B1(n_91), .B2(n_92), .Y(n_98) );
A2O1A1Ixp33_ASAP7_75t_SL g246 ( .A1(n_52), .A2(n_238), .B(n_247), .C(n_248), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_53), .Y(n_138) );
INVxp67_ASAP7_75t_L g249 ( .A(n_54), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_55), .Y(n_221) );
INVx1_ASAP7_75t_L g270 ( .A(n_56), .Y(n_270) );
INVx1_ASAP7_75t_L g516 ( .A(n_57), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_58), .A2(n_202), .B(n_213), .C(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_60), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g196 ( .A(n_61), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_62), .B(n_247), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g318 ( .A1(n_64), .A2(n_202), .B(n_213), .C(n_319), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_65), .A2(n_513), .B1(n_514), .B2(n_515), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_65), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_67), .B(n_241), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_68), .Y(n_324) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_69), .A2(n_202), .B(n_213), .C(n_285), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_70), .Y(n_292) );
INVx1_ASAP7_75t_L g245 ( .A(n_71), .Y(n_245) );
CKINVDCx16_ASAP7_75t_R g298 ( .A(n_72), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_73), .B(n_260), .Y(n_286) );
INVx1_ASAP7_75t_L g91 ( .A(n_74), .Y(n_91) );
INVx1_ASAP7_75t_L g93 ( .A(n_74), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_75), .B(n_226), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_76), .A2(n_228), .B(n_244), .Y(n_243) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_178), .B1(n_186), .B2(n_498), .C(n_506), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
INVx1_ASAP7_75t_L g176 ( .A(n_80), .Y(n_176) );
OAI322xp33_ASAP7_75t_L g506 ( .A1(n_80), .A2(n_212), .A3(n_507), .B1(n_508), .B2(n_536), .C1(n_537), .C2(n_542), .Y(n_506) );
AND2x2_ASAP7_75t_SL g80 ( .A(n_81), .B(n_142), .Y(n_80) );
INVxp67_ASAP7_75t_L g507 ( .A(n_81), .Y(n_507) );
NOR3xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_119), .C(n_133), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g82 ( .A(n_83), .B(n_107), .Y(n_82) );
INVx4_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx4_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x4_ASAP7_75t_L g87 ( .A(n_88), .B(n_97), .Y(n_87) );
AND2x4_ASAP7_75t_L g104 ( .A(n_88), .B(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g137 ( .A(n_88), .B(n_127), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_88), .B(n_112), .Y(n_141) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_94), .Y(n_88) );
AND2x2_ASAP7_75t_L g114 ( .A(n_89), .B(n_95), .Y(n_114) );
OR2x2_ASAP7_75t_L g126 ( .A(n_89), .B(n_95), .Y(n_126) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
AND2x2_ASAP7_75t_L g146 ( .A(n_90), .B(n_95), .Y(n_146) );
AND2x2_ASAP7_75t_L g155 ( .A(n_90), .B(n_100), .Y(n_155) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g96 ( .A(n_93), .Y(n_96) );
AND2x2_ASAP7_75t_L g153 ( .A(n_94), .B(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g118 ( .A(n_95), .Y(n_118) );
AND2x6_ASAP7_75t_L g163 ( .A(n_97), .B(n_114), .Y(n_163) );
AND2x4_ASAP7_75t_L g168 ( .A(n_97), .B(n_125), .Y(n_168) );
AND2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_99), .Y(n_97) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_98), .B(n_100), .Y(n_106) );
INVx1_ASAP7_75t_L g113 ( .A(n_98), .Y(n_113) );
INVx1_ASAP7_75t_L g128 ( .A(n_98), .Y(n_128) );
INVx1_ASAP7_75t_L g154 ( .A(n_98), .Y(n_154) );
AND2x2_ASAP7_75t_L g127 ( .A(n_99), .B(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g112 ( .A(n_100), .B(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
BUFx3_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OR2x6_ASAP7_75t_L g117 ( .A(n_106), .B(n_118), .Y(n_117) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx4_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx8_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
INVx1_ASAP7_75t_L g175 ( .A(n_113), .Y(n_175) );
AND2x4_ASAP7_75t_L g132 ( .A(n_114), .B(n_127), .Y(n_132) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx6_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g172 ( .A(n_118), .Y(n_172) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_121), .B1(n_129), .B2(n_130), .Y(n_119) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx5_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
INVx11_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x6_ASAP7_75t_L g145 ( .A(n_127), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OAI22xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_135), .B1(n_138), .B2(n_139), .Y(n_133) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx2_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVxp67_ASAP7_75t_L g536 ( .A(n_142), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_143), .B(n_160), .Y(n_142) );
OAI21xp5_ASAP7_75t_SL g143 ( .A1(n_144), .A2(n_147), .B(n_148), .Y(n_143) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g174 ( .A(n_146), .B(n_175), .Y(n_174) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
INVx1_ASAP7_75t_L g159 ( .A(n_154), .Y(n_159) );
AND2x4_ASAP7_75t_L g158 ( .A(n_155), .B(n_159), .Y(n_158) );
AND2x4_ASAP7_75t_L g171 ( .A(n_155), .B(n_172), .Y(n_171) );
BUFx4f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NAND3xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_164), .C(n_169), .Y(n_160) );
BUFx4f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx5_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_179), .Y(n_178) );
OR2x2_ASAP7_75t_SL g179 ( .A(n_180), .B(n_184), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND3x1_ASAP7_75t_SL g526 ( .A(n_181), .B(n_184), .C(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g532 ( .A(n_181), .B(n_533), .Y(n_532) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_181), .A2(n_539), .B(n_541), .Y(n_538) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_182), .B(n_185), .Y(n_541) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND3x1_ASAP7_75t_L g187 ( .A(n_188), .B(n_423), .C(n_472), .Y(n_187) );
NOR3xp33_ASAP7_75t_SL g188 ( .A(n_189), .B(n_330), .C(n_368), .Y(n_188) );
OAI222xp33_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_251), .B1(n_305), .B2(n_311), .C1(n_325), .C2(n_328), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_222), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_191), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_191), .B(n_373), .Y(n_464) );
BUFx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
OR2x2_ASAP7_75t_L g341 ( .A(n_192), .B(n_242), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_192), .B(n_223), .Y(n_349) );
AND2x2_ASAP7_75t_L g384 ( .A(n_192), .B(n_361), .Y(n_384) );
OR2x2_ASAP7_75t_L g408 ( .A(n_192), .B(n_223), .Y(n_408) );
OR2x2_ASAP7_75t_L g416 ( .A(n_192), .B(n_315), .Y(n_416) );
AND2x2_ASAP7_75t_L g419 ( .A(n_192), .B(n_242), .Y(n_419) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
OR2x2_ASAP7_75t_L g313 ( .A(n_193), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g327 ( .A(n_193), .B(n_242), .Y(n_327) );
AND2x2_ASAP7_75t_L g377 ( .A(n_193), .B(n_315), .Y(n_377) );
AND2x2_ASAP7_75t_L g390 ( .A(n_193), .B(n_223), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_193), .B(n_476), .Y(n_497) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_200), .B(n_220), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_194), .B(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g265 ( .A(n_194), .Y(n_265) );
AO21x2_ASAP7_75t_L g315 ( .A1(n_194), .A2(n_316), .B(n_323), .Y(n_315) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_195), .Y(n_226) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
AND2x2_ASAP7_75t_SL g241 ( .A(n_196), .B(n_197), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
OAI22xp33_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_203), .B1(n_216), .B2(n_217), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_201), .A2(n_230), .B(n_231), .C(n_232), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_201), .A2(n_231), .B(n_245), .C(n_246), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g297 ( .A1(n_201), .A2(n_231), .B(n_298), .C(n_299), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_201), .B(n_504), .Y(n_503) );
INVx4_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
NAND2x1p5_ASAP7_75t_L g217 ( .A(n_202), .B(n_218), .Y(n_217) );
AND2x4_ASAP7_75t_L g228 ( .A(n_202), .B(n_218), .Y(n_228) );
INVx2_ASAP7_75t_L g322 ( .A(n_204), .Y(n_322) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g214 ( .A(n_206), .Y(n_214) );
INVx1_ASAP7_75t_L g219 ( .A(n_206), .Y(n_219) );
OAI22xp5_ASAP7_75t_SL g207 ( .A1(n_208), .A2(n_210), .B1(n_211), .B2(n_212), .Y(n_207) );
INVx2_ASAP7_75t_L g211 ( .A(n_208), .Y(n_211) );
INVx4_ASAP7_75t_L g300 ( .A(n_208), .Y(n_300) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g215 ( .A(n_209), .Y(n_215) );
AND2x2_ASAP7_75t_L g218 ( .A(n_209), .B(n_219), .Y(n_218) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_209), .Y(n_234) );
INVx3_ASAP7_75t_L g237 ( .A(n_209), .Y(n_237) );
INVx1_ASAP7_75t_L g247 ( .A(n_209), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_210), .A2(n_510), .B1(n_524), .B2(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g502 ( .A(n_211), .Y(n_502) );
INVx5_ASAP7_75t_L g231 ( .A(n_213), .Y(n_231) );
AND2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_214), .Y(n_239) );
BUFx3_ASAP7_75t_L g264 ( .A(n_214), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g269 ( .A1(n_217), .A2(n_270), .B(n_271), .Y(n_269) );
OAI21xp5_ASAP7_75t_L g316 ( .A1(n_217), .A2(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g505 ( .A(n_219), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_L g415 ( .A1(n_222), .A2(n_416), .B(n_417), .C(n_420), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_222), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_222), .B(n_360), .Y(n_482) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_242), .Y(n_222) );
AND2x2_ASAP7_75t_SL g326 ( .A(n_223), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g340 ( .A(n_223), .Y(n_340) );
AND2x2_ASAP7_75t_L g367 ( .A(n_223), .B(n_361), .Y(n_367) );
INVx1_ASAP7_75t_SL g375 ( .A(n_223), .Y(n_375) );
AND2x2_ASAP7_75t_L g398 ( .A(n_223), .B(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_L g476 ( .A(n_223), .Y(n_476) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_227), .B(n_240), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_SL g266 ( .A(n_225), .B(n_267), .Y(n_266) );
INVx4_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_226), .A2(n_243), .B(n_250), .Y(n_242) );
BUFx2_ASAP7_75t_L g296 ( .A(n_228), .Y(n_296) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx4_ASAP7_75t_L g288 ( .A(n_234), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_237), .B(n_249), .Y(n_248) );
INVx5_ASAP7_75t_L g260 ( .A(n_237), .Y(n_260) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_239), .Y(n_289) );
INVx1_ASAP7_75t_L g278 ( .A(n_241), .Y(n_278) );
INVx2_ASAP7_75t_L g282 ( .A(n_241), .Y(n_282) );
OA21x2_ASAP7_75t_L g294 ( .A1(n_241), .A2(n_295), .B(n_304), .Y(n_294) );
BUFx2_ASAP7_75t_L g312 ( .A(n_242), .Y(n_312) );
INVx1_ASAP7_75t_L g374 ( .A(n_242), .Y(n_374) );
INVx3_ASAP7_75t_L g399 ( .A(n_242), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_251), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_279), .Y(n_251) );
INVx1_ASAP7_75t_L g395 ( .A(n_252), .Y(n_395) );
OAI32xp33_ASAP7_75t_L g401 ( .A1(n_252), .A2(n_340), .A3(n_402), .B1(n_403), .B2(n_404), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_252), .A2(n_406), .B1(n_409), .B2(n_414), .Y(n_405) );
INVx4_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g343 ( .A(n_253), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g421 ( .A(n_253), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g491 ( .A(n_253), .B(n_437), .Y(n_491) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_268), .Y(n_253) );
AND2x2_ASAP7_75t_L g306 ( .A(n_254), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g336 ( .A(n_254), .Y(n_336) );
INVx1_ASAP7_75t_L g355 ( .A(n_254), .Y(n_355) );
OR2x2_ASAP7_75t_L g363 ( .A(n_254), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g370 ( .A(n_254), .B(n_344), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_254), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g391 ( .A(n_254), .B(n_309), .Y(n_391) );
INVx3_ASAP7_75t_L g413 ( .A(n_254), .Y(n_413) );
AND2x2_ASAP7_75t_L g438 ( .A(n_254), .B(n_310), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_254), .B(n_403), .Y(n_486) );
OR2x6_ASAP7_75t_L g254 ( .A(n_255), .B(n_266), .Y(n_254) );
AOI21xp5_ASAP7_75t_SL g255 ( .A1(n_256), .A2(n_257), .B(n_265), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_261), .B(n_262), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g319 ( .A1(n_260), .A2(n_320), .B(n_321), .C(n_322), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_262), .A2(n_273), .B(n_274), .Y(n_272) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g303 ( .A(n_264), .Y(n_303) );
INVx1_ASAP7_75t_L g275 ( .A(n_265), .Y(n_275) );
INVx2_ASAP7_75t_L g310 ( .A(n_268), .Y(n_310) );
AND2x2_ASAP7_75t_L g442 ( .A(n_268), .B(n_280), .Y(n_442) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_275), .B(n_276), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_278), .B(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_278), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g484 ( .A(n_279), .Y(n_484) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_293), .Y(n_279) );
INVx1_ASAP7_75t_L g329 ( .A(n_280), .Y(n_329) );
AND2x2_ASAP7_75t_L g356 ( .A(n_280), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_280), .B(n_310), .Y(n_364) );
AND2x2_ASAP7_75t_L g422 ( .A(n_280), .B(n_345), .Y(n_422) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g308 ( .A(n_281), .Y(n_308) );
AND2x2_ASAP7_75t_L g335 ( .A(n_281), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g344 ( .A(n_281), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_281), .B(n_310), .Y(n_410) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B(n_291), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_290), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_289), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_293), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g357 ( .A(n_293), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_293), .B(n_310), .Y(n_403) );
AND2x2_ASAP7_75t_L g412 ( .A(n_293), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g437 ( .A(n_293), .Y(n_437) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g309 ( .A(n_294), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g345 ( .A(n_294), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_300), .B(n_302), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_305), .A2(n_315), .B1(n_474), .B2(n_477), .Y(n_473) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
OAI21xp5_ASAP7_75t_SL g496 ( .A1(n_307), .A2(n_418), .B(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_308), .B(n_413), .Y(n_430) );
INVx1_ASAP7_75t_L g455 ( .A(n_308), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_309), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g382 ( .A(n_309), .B(n_335), .Y(n_382) );
INVx2_ASAP7_75t_L g338 ( .A(n_310), .Y(n_338) );
INVx1_ASAP7_75t_L g388 ( .A(n_310), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g479 ( .A1(n_311), .A2(n_463), .B1(n_480), .B2(n_483), .C(n_485), .Y(n_479) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g350 ( .A(n_312), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_312), .B(n_361), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_313), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g404 ( .A(n_313), .B(n_350), .Y(n_404) );
INVx3_ASAP7_75t_SL g445 ( .A(n_313), .Y(n_445) );
AND2x2_ASAP7_75t_L g389 ( .A(n_314), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g418 ( .A(n_314), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_314), .B(n_327), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_314), .B(n_373), .Y(n_459) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx3_ASAP7_75t_L g361 ( .A(n_315), .Y(n_361) );
OAI322xp33_ASAP7_75t_L g456 ( .A1(n_315), .A2(n_387), .A3(n_409), .B1(n_457), .B2(n_459), .C1(n_460), .C2(n_461), .Y(n_456) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI21xp33_ASAP7_75t_L g480 ( .A1(n_326), .A2(n_329), .B(n_481), .Y(n_480) );
NOR2xp33_ASAP7_75t_SL g406 ( .A(n_327), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g428 ( .A(n_327), .B(n_340), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_327), .B(n_367), .Y(n_443) );
INVxp67_ASAP7_75t_L g394 ( .A(n_329), .Y(n_394) );
AOI211xp5_ASAP7_75t_L g400 ( .A1(n_329), .A2(n_401), .B(n_405), .C(n_415), .Y(n_400) );
OAI221xp5_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_339), .B1(n_342), .B2(n_346), .C(n_351), .Y(n_330) );
INVxp67_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_337), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g354 ( .A(n_338), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g471 ( .A(n_338), .Y(n_471) );
OAI221xp5_ASAP7_75t_L g487 ( .A1(n_339), .A2(n_488), .B1(n_493), .B2(n_494), .C(n_496), .Y(n_487) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_340), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g387 ( .A(n_340), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_340), .B(n_418), .Y(n_425) );
AND2x2_ASAP7_75t_L g467 ( .A(n_340), .B(n_445), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_341), .B(n_366), .Y(n_365) );
OAI22xp33_ASAP7_75t_L g462 ( .A1(n_341), .A2(n_353), .B1(n_463), .B2(n_464), .Y(n_462) );
OR2x2_ASAP7_75t_L g493 ( .A(n_341), .B(n_361), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g470 ( .A(n_344), .Y(n_470) );
AND2x2_ASAP7_75t_L g495 ( .A(n_344), .B(n_438), .Y(n_495) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR2xp33_ASAP7_75t_SL g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g359 ( .A(n_349), .B(n_360), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_358), .B1(n_362), .B2(n_365), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g426 ( .A(n_354), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_354), .B(n_394), .Y(n_461) );
AOI322xp5_ASAP7_75t_L g385 ( .A1(n_356), .A2(n_386), .A3(n_388), .B1(n_389), .B2(n_391), .C1(n_392), .C2(n_396), .Y(n_385) );
INVxp67_ASAP7_75t_L g379 ( .A(n_357), .Y(n_379) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_359), .A2(n_364), .B1(n_381), .B2(n_383), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_360), .B(n_373), .Y(n_460) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_361), .B(n_399), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_361), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g457 ( .A(n_363), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
NAND3xp33_ASAP7_75t_SL g368 ( .A(n_369), .B(n_385), .C(n_400), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B1(n_376), .B2(n_378), .C(n_380), .Y(n_369) );
AND2x2_ASAP7_75t_L g376 ( .A(n_372), .B(n_377), .Y(n_376) );
INVx3_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
AND2x2_ASAP7_75t_L g386 ( .A(n_377), .B(n_387), .Y(n_386) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_379), .Y(n_458) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_384), .B(n_398), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_387), .B(n_445), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_388), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g463 ( .A(n_391), .Y(n_463) );
AND2x2_ASAP7_75t_L g478 ( .A(n_391), .B(n_455), .Y(n_478) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AOI211xp5_ASAP7_75t_L g472 ( .A1(n_402), .A2(n_473), .B(n_479), .C(n_487), .Y(n_472) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g441 ( .A(n_412), .B(n_442), .Y(n_441) );
NAND2x1_ASAP7_75t_SL g483 ( .A(n_413), .B(n_484), .Y(n_483) );
CKINVDCx16_ASAP7_75t_R g453 ( .A(n_416), .Y(n_453) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g448 ( .A(n_422), .Y(n_448) );
AND2x2_ASAP7_75t_L g452 ( .A(n_422), .B(n_438), .Y(n_452) );
NOR5xp2_ASAP7_75t_L g423 ( .A(n_424), .B(n_439), .C(n_456), .D(n_462), .E(n_465), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_427), .B2(n_429), .C(n_431), .Y(n_424) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_428), .B(n_486), .Y(n_485) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g454 ( .A(n_438), .B(n_455), .Y(n_454) );
OAI221xp5_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_443), .B1(n_444), .B2(n_446), .C(n_449), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_452), .B1(n_453), .B2(n_454), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g492 ( .A(n_452), .Y(n_492) );
AOI211xp5_ASAP7_75t_SL g465 ( .A1(n_466), .A2(n_468), .B(n_470), .C(n_471), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVxp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_492), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
CKINVDCx14_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .Y(n_500) );
INVx1_ASAP7_75t_L g540 ( .A(n_501), .Y(n_540) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_504), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_510), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_517), .B2(n_523), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_517), .Y(n_523) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
INVxp67_ASAP7_75t_L g535 ( .A(n_527), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_532), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_534), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g537 ( .A(n_538), .Y(n_537) );
CKINVDCx16_ASAP7_75t_R g543 ( .A(n_544), .Y(n_543) );
endmodule