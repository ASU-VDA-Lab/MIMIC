module fake_jpeg_19229_n_254 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_254);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx6_ASAP7_75t_SL g11 ( 
.A(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_SL g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_25),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_32),
.B(n_33),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_12),
.B1(n_11),
.B2(n_23),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_12),
.B1(n_24),
.B2(n_11),
.Y(n_46)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_42),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_47),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_12),
.B1(n_30),
.B2(n_15),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_12),
.B1(n_36),
.B2(n_39),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_50),
.Y(n_61)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_53),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_25),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_34),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_56),
.B(n_34),
.Y(n_74)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_72),
.Y(n_85)
);

INVxp67_ASAP7_75t_SL g62 ( 
.A(n_54),
.Y(n_62)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_36),
.B(n_39),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_81),
.B(n_73),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_84),
.Y(n_97)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_86),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_56),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_51),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_69),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_53),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_20),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_84),
.A2(n_73),
.B1(n_70),
.B2(n_46),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_98),
.B1(n_37),
.B2(n_15),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_103),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_32),
.B(n_25),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_102),
.B(n_40),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_79),
.B(n_29),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_40),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_89),
.B1(n_77),
.B2(n_92),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_35),
.B1(n_49),
.B2(n_43),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_99),
.A2(n_109),
.B1(n_63),
.B2(n_64),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_67),
.C(n_35),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_104),
.C(n_108),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_80),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_44),
.B(n_28),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_35),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_33),
.C(n_31),
.Y(n_104)
);

OAI22x1_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_40),
.B1(n_28),
.B2(n_27),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_37),
.B1(n_64),
.B2(n_58),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_33),
.C(n_31),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_43),
.B1(n_49),
.B2(n_57),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_23),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_120),
.Y(n_154)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_138),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_116),
.A2(n_134),
.B(n_27),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_94),
.C(n_96),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_18),
.C(n_13),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_119),
.Y(n_144)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_78),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_40),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_78),
.Y(n_126)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_64),
.B1(n_63),
.B2(n_86),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_129),
.B1(n_133),
.B2(n_68),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_100),
.B(n_20),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_132),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_88),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_37),
.B1(n_71),
.B2(n_11),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_102),
.A2(n_88),
.B(n_60),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_71),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_68),
.B(n_26),
.Y(n_155)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_136),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_78),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_137),
.B(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_149),
.Y(n_176)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_143),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_71),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_152),
.B(n_119),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_18),
.C(n_13),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_157),
.C(n_158),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_155),
.A2(n_135),
.B1(n_147),
.B2(n_134),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_131),
.A2(n_33),
.B1(n_31),
.B2(n_54),
.Y(n_156)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_18),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_14),
.B1(n_21),
.B2(n_19),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_150),
.B1(n_156),
.B2(n_153),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_179),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_113),
.C(n_136),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_170),
.C(n_174),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_147),
.A2(n_140),
.B1(n_144),
.B2(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_138),
.C(n_122),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_120),
.Y(n_172)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_9),
.B1(n_10),
.B2(n_8),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_118),
.C(n_125),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_118),
.C(n_27),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_26),
.C(n_21),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_141),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_195),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_181),
.A2(n_159),
.B1(n_155),
.B2(n_162),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g199 ( 
.A1(n_185),
.A2(n_196),
.A3(n_168),
.B1(n_189),
.B2(n_197),
.C1(n_187),
.C2(n_191),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_186),
.A2(n_180),
.B1(n_164),
.B2(n_175),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_9),
.Y(n_188)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_9),
.B1(n_10),
.B2(n_8),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_190),
.A2(n_5),
.B1(n_1),
.B2(n_2),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_179),
.A2(n_8),
.B(n_7),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_3),
.B(n_4),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_26),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_18),
.Y(n_195)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_192),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_201),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_203),
.B1(n_205),
.B2(n_193),
.Y(n_218)
);

FAx1_ASAP7_75t_SL g201 ( 
.A(n_182),
.B(n_184),
.CI(n_165),
.CON(n_201),
.SN(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_170),
.C(n_174),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_209),
.C(n_207),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_7),
.B(n_5),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_204),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_211),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_21),
.C(n_19),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_190),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_217),
.Y(n_229)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_195),
.Y(n_217)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_201),
.C(n_200),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_219),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_194),
.B(n_14),
.Y(n_220)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_206),
.B(n_14),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_211),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_224),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_210),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_227),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_219),
.B(n_205),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_213),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_234),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_217),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_212),
.C(n_221),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_235),
.B(n_237),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_14),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_13),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_238),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_230),
.A2(n_21),
.B1(n_13),
.B2(n_4),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_239),
.A2(n_3),
.B(n_4),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_236),
.A2(n_231),
.B1(n_224),
.B2(n_13),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_241),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_233),
.B(n_232),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_245),
.A2(n_244),
.B1(n_4),
.B2(n_3),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_242),
.A2(n_237),
.B(n_13),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

NOR3xp33_ASAP7_75t_SL g251 ( 
.A(n_250),
.B(n_249),
.C(n_247),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_251),
.B(n_3),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_SL g253 ( 
.A1(n_252),
.A2(n_22),
.B(n_233),
.C(n_248),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_22),
.Y(n_254)
);


endmodule