module real_jpeg_2262_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_361, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_361;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_0),
.B(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_0),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_0),
.B(n_69),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_0),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_0),
.B(n_43),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_0),
.B(n_34),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_2),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_2),
.B(n_43),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_2),
.B(n_72),
.Y(n_256)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_4),
.B(n_43),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_4),
.B(n_54),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_4),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_4),
.B(n_61),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_4),
.B(n_72),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_6),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_6),
.B(n_43),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_6),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_6),
.B(n_39),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_6),
.B(n_31),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_6),
.B(n_69),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_6),
.B(n_61),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_10),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_10),
.B(n_54),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_10),
.B(n_39),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_10),
.B(n_61),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_10),
.B(n_69),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_11),
.B(n_43),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_11),
.B(n_72),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_11),
.B(n_34),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_11),
.B(n_54),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_11),
.B(n_61),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_11),
.B(n_69),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_12),
.B(n_69),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_12),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_12),
.B(n_61),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_12),
.B(n_72),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_12),
.B(n_34),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_12),
.B(n_54),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_12),
.B(n_39),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_13),
.B(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_13),
.B(n_34),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_13),
.B(n_39),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_13),
.B(n_54),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_13),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_13),
.B(n_43),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_13),
.B(n_72),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

XNOR2x2_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_158),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_157),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_135),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_20),
.B(n_135),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_83),
.C(n_102),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_21),
.B(n_83),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_64),
.B2(n_82),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_22),
.B(n_65),
.C(n_74),
.Y(n_156)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.C(n_48),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_24),
.B(n_342),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_36),
.B2(n_37),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_35),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_28),
.B(n_33),
.C(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_29),
.B(n_38),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_30),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_30),
.B(n_40),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_30),
.B(n_173),
.Y(n_291)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_67),
.C(n_68),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_33),
.A2(n_35),
.B1(n_67),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_33),
.A2(n_35),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_33),
.B(n_190),
.Y(n_230)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_34),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_36),
.A2(n_37),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_36),
.B(n_290),
.C(n_291),
.Y(n_320)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_38),
.B(n_173),
.Y(n_196)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_40),
.B(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_41),
.A2(n_48),
.B1(n_49),
.B2(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_41),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.C(n_47),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_42),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_42),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_45),
.A2(n_46),
.B1(n_47),
.B2(n_120),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_47),
.Y(n_120)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_56),
.B2(n_63),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_51),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_50),
.A2(n_51),
.B1(n_126),
.B2(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_50),
.B(n_229),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_57),
.C(n_60),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_51),
.B(n_86),
.C(n_89),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_53),
.B(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_53),
.B(n_173),
.Y(n_200)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_61),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_74),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.C(n_71),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_66),
.B(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_67),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_67),
.A2(n_109),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_67),
.B(n_246),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_68),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_68),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_68),
.A2(n_110),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx3_ASAP7_75t_SL g183 ( 
.A(n_69),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_70),
.A2(n_71),
.B1(n_81),
.B2(n_134),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_70),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_71),
.A2(n_77),
.B1(n_78),
.B2(n_81),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_71),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_71),
.B(n_75),
.C(n_78),
.Y(n_149)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_72),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_80),
.B(n_124),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_91),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_84),
.B(n_92),
.C(n_93),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_85),
.A2(n_86),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_85),
.A2(n_86),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_86),
.B(n_240),
.C(n_241),
.Y(n_276)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_89),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_100),
.B2(n_101),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_96),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_97),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_112),
.C(n_114),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_99),
.C(n_101),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_97),
.A2(n_98),
.B1(n_114),
.B2(n_115),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_102),
.A2(n_103),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_121),
.C(n_132),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_104),
.A2(n_105),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_111),
.C(n_116),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_106),
.B(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_111),
.B(n_116),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_112),
.B(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_121),
.B(n_132),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_128),
.C(n_130),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_122),
.B(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.C(n_126),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_123),
.A2(n_126),
.B1(n_229),
.B2(n_303),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_123),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_124),
.B(n_127),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_124),
.B(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_125),
.A2(n_301),
.B1(n_302),
.B2(n_304),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_125),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_126),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_330)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx24_ASAP7_75t_SL g360 ( 
.A(n_135),
.Y(n_360)
);

FAx1_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_147),
.CI(n_156),
.CON(n_135),
.SN(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_144),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_139),
.A2(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_139),
.B(n_282),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_155),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_153),
.Y(n_154)
);

AOI321xp33_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_336),
.A3(n_348),
.B1(n_353),
.B2(n_358),
.C(n_361),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_293),
.C(n_332),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_260),
.B(n_292),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_232),
.B(n_259),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_212),
.B(n_231),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_193),
.B(n_211),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_175),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_165),
.B(n_175),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.C(n_174),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_166),
.A2(n_167),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_167),
.A2(n_168),
.B(n_169),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_170),
.A2(n_171),
.B1(n_174),
.B2(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_172),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_183),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_174),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_184),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_185),
.C(n_189),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_182),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_178),
.B(n_181),
.C(n_182),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_183),
.B(n_223),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_188),
.B1(n_189),
.B2(n_192),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_192),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_202),
.B(n_210),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_198),
.B(n_201),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_196),
.B(n_197),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_203),
.B(n_206),
.Y(n_210)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_213),
.B(n_214),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_225),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_224),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_224),
.C(n_225),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_221),
.C(n_222),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_219),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_228),
.C(n_230),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_233),
.B(n_234),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_248),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_249),
.C(n_250),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_242),
.B2(n_243),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_244),
.C(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_245),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_258),
.Y(n_250)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_251),
.Y(n_258)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_257),
.C(n_258),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_256),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_261),
.B(n_262),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_279),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_277),
.B2(n_278),
.Y(n_263)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_265),
.B(n_278),
.C(n_279),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_274),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_275),
.C(n_276),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_267),
.B(n_271),
.C(n_273),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_270),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_287),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_280)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_281),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_283),
.B(n_308),
.C(n_311),
.Y(n_328)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_284),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_285),
.C(n_287),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_291),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI21xp33_ASAP7_75t_L g354 ( 
.A1(n_294),
.A2(n_355),
.B(n_356),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_321),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_295),
.B(n_321),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_312),
.C(n_313),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_296),
.B(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_299),
.C(n_306),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_305),
.B2(n_306),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_302),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_310),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_313),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_320),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_318),
.C(n_320),
.Y(n_326)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_331),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_325),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_325),
.C(n_331),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_328),
.C(n_329),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_333),
.B(n_334),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_345),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_337),
.B(n_345),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_341),
.C(n_344),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_338),
.B(n_341),
.Y(n_352)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_344),
.B(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_346),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_349),
.A2(n_354),
.B(n_357),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_350),
.B(n_351),
.Y(n_357)
);


endmodule