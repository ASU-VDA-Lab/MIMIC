module fake_jpeg_679_n_551 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_551);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_551;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_11),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_60),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_62),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_63),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_64),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_65),
.Y(n_205)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_66),
.Y(n_208)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_67),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_68),
.Y(n_178)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_70),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_73),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_74),
.Y(n_173)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

INVx11_ASAP7_75t_SL g76 ( 
.A(n_25),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_27),
.B(n_18),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_77),
.B(n_80),
.Y(n_147)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_78),
.Y(n_168)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_79),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_0),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_81),
.Y(n_175)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_82),
.Y(n_172)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g181 ( 
.A(n_83),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_85),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_87),
.Y(n_166)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_30),
.Y(n_88)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_89),
.Y(n_176)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_19),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_99),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_91),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_94),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_96),
.Y(n_187)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_27),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_37),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_102),
.Y(n_150)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_19),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_25),
.Y(n_104)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

CKINVDCx10_ASAP7_75t_R g105 ( 
.A(n_25),
.Y(n_105)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_105),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_54),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_112),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_24),
.B(n_0),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_113),
.Y(n_158)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_19),
.Y(n_110)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_29),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_21),
.B(n_17),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_21),
.B(n_17),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_1),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_118),
.Y(n_139)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_116),
.B(n_122),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_34),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_117),
.B(n_123),
.Y(n_182)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

HAxp5_ASAP7_75t_SL g119 ( 
.A(n_29),
.B(n_1),
.CON(n_119),
.SN(n_119)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_119),
.A2(n_10),
.B(n_12),
.Y(n_201)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_120),
.B(n_121),
.Y(n_174)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_44),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_44),
.Y(n_123)
);

INVx6_ASAP7_75t_SL g124 ( 
.A(n_51),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_124),
.B(n_6),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_90),
.A2(n_47),
.B1(n_42),
.B2(n_36),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_126),
.A2(n_128),
.B1(n_130),
.B2(n_133),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_102),
.A2(n_104),
.B1(n_76),
.B2(n_60),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_61),
.A2(n_42),
.B1(n_34),
.B2(n_36),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_62),
.A2(n_47),
.B1(n_55),
.B2(n_39),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_63),
.A2(n_33),
.B1(n_53),
.B2(n_52),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_135),
.A2(n_149),
.B1(n_155),
.B2(n_156),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_98),
.A2(n_33),
.B1(n_53),
.B2(n_52),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_140),
.A2(n_16),
.B1(n_200),
.B2(n_157),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_55),
.B(n_48),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g216 ( 
.A1(n_144),
.A2(n_161),
.B(n_15),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_74),
.A2(n_48),
.B1(n_35),
.B2(n_39),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_64),
.A2(n_43),
.B1(n_41),
.B2(n_40),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_70),
.A2(n_43),
.B1(n_41),
.B2(n_40),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_91),
.A2(n_35),
.B1(n_38),
.B2(n_46),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_160),
.A2(n_167),
.B1(n_184),
.B2(n_132),
.Y(n_227)
);

AOI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_67),
.A2(n_46),
.B(n_38),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_165),
.B(n_193),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_123),
.A2(n_46),
.B1(n_44),
.B2(n_4),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_117),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_170),
.B(n_197),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_88),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_171),
.A2(n_167),
.B(n_195),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_123),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_65),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_186),
.A2(n_195),
.B1(n_16),
.B2(n_184),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_110),
.B(n_3),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_194),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_84),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_58),
.B(n_7),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_58),
.B(n_16),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_203),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_118),
.B(n_8),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_199),
.B(n_202),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_12),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_122),
.B(n_115),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_89),
.B(n_10),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_121),
.B(n_12),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_206),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_86),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_136),
.Y(n_209)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_209),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_210),
.B(n_216),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_158),
.B(n_95),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_211),
.B(n_218),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_L g214 ( 
.A1(n_160),
.A2(n_94),
.B1(n_106),
.B2(n_87),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_214),
.A2(n_235),
.B1(n_205),
.B2(n_257),
.Y(n_296)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_164),
.Y(n_215)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_215),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_133),
.A2(n_92),
.B1(n_96),
.B2(n_103),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_217),
.A2(n_228),
.B1(n_240),
.B2(n_247),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_163),
.B(n_107),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_137),
.Y(n_219)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_219),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_142),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_220),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_168),
.B(n_15),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_221),
.B(n_223),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_169),
.B(n_175),
.Y(n_223)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_137),
.Y(n_224)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_224),
.Y(n_284)
);

BUFx12f_ASAP7_75t_L g225 ( 
.A(n_137),
.Y(n_225)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_225),
.Y(n_287)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_151),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_226),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_227),
.Y(n_301)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_151),
.Y(n_229)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_229),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_142),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_230),
.Y(n_330)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_233),
.Y(n_303)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_164),
.Y(n_234)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_234),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_SL g236 ( 
.A(n_147),
.B(n_150),
.C(n_134),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_236),
.Y(n_305)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_145),
.Y(n_237)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_237),
.Y(n_297)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_176),
.Y(n_238)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_238),
.Y(n_298)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_239),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_208),
.A2(n_196),
.B1(n_178),
.B2(n_143),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_152),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_241),
.B(n_242),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_174),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_127),
.B(n_182),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_243),
.B(n_246),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_125),
.B(n_174),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_244),
.B(n_253),
.C(n_263),
.Y(n_326)
);

AO22x1_ASAP7_75t_SL g245 ( 
.A1(n_139),
.A2(n_154),
.B1(n_131),
.B2(n_207),
.Y(n_245)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_245),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_196),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_208),
.A2(n_178),
.B1(n_143),
.B2(n_189),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_159),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_248),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_129),
.B(n_138),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_250),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_138),
.B(n_181),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_189),
.A2(n_132),
.B1(n_207),
.B2(n_191),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_252),
.A2(n_278),
.B1(n_258),
.B2(n_246),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_172),
.B(n_181),
.Y(n_253)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_179),
.Y(n_254)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_254),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_136),
.Y(n_255)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_255),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_128),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_265),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_148),
.Y(n_258)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_258),
.Y(n_321)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_139),
.Y(n_259)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_148),
.Y(n_260)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_260),
.Y(n_328)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_173),
.Y(n_262)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_262),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_172),
.B(n_183),
.C(n_188),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_201),
.B(n_126),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_264),
.B(n_270),
.Y(n_322)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_159),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_187),
.B(n_141),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_267),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_192),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_268),
.B(n_269),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_192),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_187),
.B(n_156),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_141),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_271),
.B(n_272),
.Y(n_320)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_146),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_173),
.B(n_179),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_273),
.B(n_274),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_146),
.B(n_177),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_149),
.B(n_153),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_275),
.Y(n_308)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_153),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_276),
.A2(n_258),
.B1(n_272),
.B2(n_260),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_166),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_277),
.A2(n_180),
.B(n_185),
.Y(n_281)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_180),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_270),
.A2(n_186),
.B1(n_166),
.B2(n_177),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_280),
.A2(n_296),
.B1(n_304),
.B2(n_309),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_281),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_264),
.A2(n_162),
.B(n_185),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_292),
.A2(n_294),
.B(n_301),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_210),
.A2(n_162),
.B(n_205),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_294),
.A2(n_253),
.B(n_224),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_211),
.A2(n_228),
.B1(n_218),
.B2(n_256),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_306),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_259),
.A2(n_235),
.B1(n_232),
.B2(n_221),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g361 ( 
.A(n_310),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_213),
.A2(n_267),
.B1(n_231),
.B2(n_223),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_314),
.A2(n_324),
.B1(n_329),
.B2(n_278),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_251),
.B(n_261),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_219),
.C(n_209),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_222),
.A2(n_212),
.B1(n_214),
.B2(n_268),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_263),
.B1(n_238),
.B2(n_254),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_245),
.A2(n_210),
.B1(n_244),
.B2(n_276),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_245),
.A2(n_244),
.B1(n_237),
.B2(n_239),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_283),
.B(n_241),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_332),
.B(n_339),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_302),
.A2(n_271),
.B1(n_233),
.B2(n_234),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_334),
.A2(n_363),
.B1(n_367),
.B2(n_279),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_335),
.A2(n_352),
.B1(n_354),
.B2(n_298),
.Y(n_381)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_321),
.Y(n_336)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_336),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_320),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_337),
.B(n_345),
.Y(n_377)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_321),
.Y(n_338)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_338),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_295),
.B(n_215),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_299),
.Y(n_340)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_340),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_295),
.B(n_253),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_341),
.B(n_344),
.Y(n_389)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_299),
.Y(n_342)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_342),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_312),
.B(n_229),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_283),
.B(n_226),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_346),
.A2(n_358),
.B(n_371),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_316),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_348),
.Y(n_387)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_303),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_262),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_349),
.A2(n_355),
.B(n_287),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_351),
.B(n_353),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_302),
.A2(n_220),
.B1(n_230),
.B2(n_248),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_312),
.B(n_255),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_322),
.B(n_225),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_265),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_356),
.B(n_365),
.C(n_327),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_304),
.B(n_225),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_357),
.B(n_359),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_286),
.A2(n_225),
.B(n_308),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_328),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_360),
.Y(n_374)
);

OA21x2_ASAP7_75t_L g362 ( 
.A1(n_314),
.A2(n_292),
.B(n_329),
.Y(n_362)
);

AO22x2_ASAP7_75t_L g392 ( 
.A1(n_362),
.A2(n_311),
.B1(n_297),
.B2(n_293),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_309),
.A2(n_280),
.B1(n_324),
.B2(n_296),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_282),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_364),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_326),
.B(n_325),
.C(n_290),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_282),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_366),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_308),
.A2(n_301),
.B1(n_325),
.B2(n_288),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_291),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_368),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_307),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_369),
.Y(n_395)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_303),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_370),
.Y(n_399)
);

O2A1O1Ixp33_ASAP7_75t_L g372 ( 
.A1(n_281),
.A2(n_285),
.B(n_291),
.C(n_298),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_372),
.A2(n_319),
.B(n_284),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_375),
.C(n_378),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_315),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_376),
.A2(n_357),
.B1(n_335),
.B2(n_350),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_365),
.B(n_290),
.C(n_289),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_381),
.A2(n_393),
.B1(n_398),
.B2(n_352),
.Y(n_423)
);

AND2x2_ASAP7_75t_SL g382 ( 
.A(n_354),
.B(n_290),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_382),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_333),
.A2(n_305),
.B1(n_311),
.B2(n_331),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_384),
.A2(n_402),
.B1(n_338),
.B2(n_368),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_341),
.B(n_331),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_386),
.B(n_388),
.C(n_336),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_353),
.B(n_297),
.Y(n_388)
);

OAI21x1_ASAP7_75t_SL g430 ( 
.A1(n_392),
.A2(n_401),
.B(n_403),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_333),
.A2(n_305),
.B1(n_300),
.B2(n_330),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_363),
.A2(n_350),
.B1(n_367),
.B2(n_343),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_332),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_400),
.B(n_364),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_362),
.A2(n_300),
.B1(n_330),
.B2(n_318),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_387),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_407),
.B(n_408),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_339),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_385),
.Y(n_409)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_409),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_369),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_410),
.B(n_413),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_377),
.B(n_344),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_411),
.B(n_418),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_412),
.A2(n_429),
.B1(n_432),
.B2(n_403),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_395),
.B(n_337),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_375),
.B(n_351),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_414),
.B(n_415),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_362),
.Y(n_415)
);

OAI32xp33_ASAP7_75t_L g416 ( 
.A1(n_389),
.A2(n_362),
.A3(n_349),
.B1(n_372),
.B2(n_359),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_416),
.A2(n_419),
.B(n_396),
.Y(n_447)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_385),
.Y(n_417)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_417),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_377),
.B(n_349),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_396),
.A2(n_358),
.B(n_371),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_379),
.B(n_347),
.Y(n_420)
);

NAND3xp33_ASAP7_75t_L g451 ( 
.A(n_420),
.B(n_421),
.C(n_422),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_380),
.B(n_348),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_423),
.A2(n_434),
.B1(n_390),
.B2(n_380),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_379),
.B(n_355),
.Y(n_424)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_424),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_389),
.B(n_355),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_425),
.B(n_428),
.Y(n_459)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_383),
.Y(n_427)
);

NAND2x1_ASAP7_75t_SL g455 ( 
.A(n_427),
.B(n_431),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_388),
.B(n_372),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_398),
.A2(n_361),
.B1(n_346),
.B2(n_366),
.Y(n_429)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_383),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_376),
.A2(n_393),
.B1(n_381),
.B2(n_402),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_433),
.B(n_378),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_437),
.A2(n_439),
.B1(n_441),
.B2(n_444),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_421),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_438),
.B(n_340),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_440),
.B(n_445),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_432),
.A2(n_401),
.B1(n_404),
.B2(n_384),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_406),
.B(n_394),
.C(n_386),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_442),
.B(n_449),
.C(n_452),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_434),
.A2(n_430),
.B1(n_426),
.B2(n_423),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_406),
.B(n_414),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_429),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_446),
.Y(n_471)
);

OA21x2_ASAP7_75t_L g467 ( 
.A1(n_447),
.A2(n_425),
.B(n_418),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_415),
.B(n_394),
.C(n_382),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_433),
.B(n_382),
.C(n_404),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_419),
.B(n_382),
.C(n_397),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_453),
.B(n_454),
.C(n_458),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_397),
.C(n_387),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_428),
.B(n_392),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_411),
.B(n_412),
.C(n_408),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_460),
.B(n_392),
.Y(n_469)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_455),
.Y(n_462)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_462),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_407),
.Y(n_463)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_463),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_457),
.B(n_424),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_464),
.B(n_469),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_455),
.B(n_422),
.Y(n_465)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_465),
.Y(n_493)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_435),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_466),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_467),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_459),
.Y(n_483)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_436),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_475),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_439),
.A2(n_446),
.B1(n_437),
.B2(n_441),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_474),
.A2(n_478),
.B1(n_458),
.B2(n_447),
.Y(n_491)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_451),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_445),
.B(n_392),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_477),
.B(n_479),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_444),
.A2(n_430),
.B1(n_416),
.B2(n_392),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_460),
.B(n_405),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_443),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_480),
.B(n_481),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_456),
.B(n_391),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_454),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_482),
.B(n_452),
.Y(n_498)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_483),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_457),
.C(n_442),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_497),
.C(n_472),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_491),
.A2(n_464),
.B1(n_472),
.B2(n_417),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_465),
.B(n_453),
.Y(n_495)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_495),
.Y(n_509)
);

AO221x1_ASAP7_75t_L g496 ( 
.A1(n_474),
.A2(n_374),
.B1(n_448),
.B2(n_390),
.C(n_391),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_496),
.B(n_498),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_461),
.B(n_440),
.C(n_449),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_463),
.B(n_370),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_499),
.A2(n_448),
.B1(n_374),
.B2(n_405),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_501),
.B(n_511),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_494),
.A2(n_473),
.B(n_478),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_502),
.A2(n_505),
.B(n_484),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_476),
.Y(n_504)
);

NOR2xp67_ASAP7_75t_SL g513 ( 
.A(n_504),
.B(n_507),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_494),
.A2(n_467),
.B(n_473),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_488),
.A2(n_471),
.B1(n_467),
.B2(n_469),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_506),
.A2(n_508),
.B1(n_484),
.B2(n_493),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_492),
.B(n_476),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_488),
.A2(n_477),
.B1(n_431),
.B2(n_427),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_510),
.A2(n_495),
.B1(n_493),
.B2(n_489),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_491),
.B(n_409),
.Y(n_511)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_512),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_501),
.B(n_487),
.C(n_497),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_514),
.B(n_516),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_515),
.A2(n_519),
.B(n_505),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_495),
.C(n_486),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_489),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_517),
.B(n_522),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_511),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_509),
.B(n_485),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_502),
.A2(n_489),
.B1(n_483),
.B2(n_496),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_523),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_490),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_524),
.B(n_525),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_515),
.A2(n_509),
.B(n_510),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_526),
.A2(n_529),
.B(n_500),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_514),
.B(n_506),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_528),
.B(n_531),
.Y(n_537)
);

AOI21xp33_ASAP7_75t_L g529 ( 
.A1(n_518),
.A2(n_500),
.B(n_508),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_516),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_533),
.B(n_539),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_527),
.B(n_523),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_534),
.A2(n_536),
.B(n_538),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_530),
.B(n_521),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_525),
.B(n_519),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_537),
.B(n_531),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_542),
.B(n_507),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_535),
.A2(n_534),
.B1(n_518),
.B2(n_512),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_543),
.A2(n_399),
.B(n_360),
.Y(n_546)
);

OAI21xp33_ASAP7_75t_L g547 ( 
.A1(n_544),
.A2(n_545),
.B(n_546),
.Y(n_547)
);

NAND4xp25_ASAP7_75t_L g545 ( 
.A(n_540),
.B(n_513),
.C(n_399),
.D(n_342),
.Y(n_545)
);

AOI322xp5_ASAP7_75t_SL g548 ( 
.A1(n_544),
.A2(n_541),
.A3(n_318),
.B1(n_330),
.B2(n_287),
.C1(n_313),
.C2(n_284),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_548),
.A2(n_313),
.B(n_319),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_547),
.B(n_293),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_550),
.A2(n_323),
.B(n_318),
.Y(n_551)
);


endmodule