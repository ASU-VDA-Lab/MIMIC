module fake_jpeg_22489_n_192 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_192);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_39),
.Y(n_65)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_40),
.A2(n_23),
.B1(n_17),
.B2(n_24),
.Y(n_71)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_15),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_16),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_15),
.B(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_19),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_16),
.C(n_28),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_22),
.C(n_24),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_51),
.B(n_55),
.Y(n_99)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_59),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_33),
.A2(n_30),
.B1(n_27),
.B2(n_18),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_57),
.A2(n_37),
.B1(n_35),
.B2(n_29),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_34),
.B(n_17),
.Y(n_68)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_64),
.B1(n_67),
.B2(n_66),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_37),
.B1(n_25),
.B2(n_2),
.Y(n_95)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_34),
.B(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_61),
.B1(n_57),
.B2(n_55),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_77),
.A2(n_80),
.B1(n_83),
.B2(n_89),
.Y(n_109)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_22),
.B1(n_41),
.B2(n_20),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_87),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_12),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_41),
.B1(n_29),
.B2(n_35),
.Y(n_83)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_95),
.B1(n_100),
.B2(n_75),
.Y(n_105)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_97),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_8),
.C(n_14),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_42),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_102),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_100),
.A2(n_75),
.B1(n_69),
.B2(n_54),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_0),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_98),
.A2(n_76),
.B(n_50),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_101),
.B(n_93),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_139)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_112),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_76),
.B1(n_50),
.B2(n_69),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_65),
.B1(n_49),
.B2(n_4),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_65),
.B1(n_12),
.B2(n_13),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_87),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_65),
.B(n_3),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_121),
.B(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_123),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_1),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_121),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_1),
.B1(n_3),
.B2(n_6),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_122),
.C(n_124),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_6),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_6),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_78),
.B1(n_85),
.B2(n_96),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_125),
.A2(n_134),
.B(n_126),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_118),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_130),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

INVxp33_ASAP7_75t_SL g132 ( 
.A(n_118),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_116),
.A2(n_93),
.B1(n_86),
.B2(n_90),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_117),
.Y(n_135)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_99),
.Y(n_137)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_111),
.B(n_79),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_138),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_119),
.B(n_85),
.Y(n_140)
);

OAI21x1_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_142),
.B(n_113),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_108),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_122),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_109),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_114),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_144),
.A2(n_155),
.B(n_127),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_157),
.Y(n_160)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_150),
.B(n_131),
.CI(n_134),
.CON(n_161),
.SN(n_161)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_151),
.B(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_109),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_152),
.B(n_145),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_110),
.C(n_103),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_143),
.C(n_139),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_136),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_144),
.C(n_146),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_152),
.A2(n_133),
.B1(n_156),
.B2(n_130),
.Y(n_159)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_165),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_148),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_166),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_127),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_164),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_154),
.B(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_168),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_147),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_160),
.Y(n_172)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_163),
.C(n_164),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_161),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_165),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_161),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_179),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_171),
.C(n_180),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_158),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_182),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_160),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_169),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_176),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_172),
.B(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_187),
.B(n_189),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_186),
.C(n_183),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_185),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_191),
.Y(n_192)
);


endmodule