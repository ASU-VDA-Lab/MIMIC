module fake_jpeg_23542_n_322 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_0),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_39),
.A2(n_45),
.B(n_1),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_40),
.Y(n_85)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx12_ASAP7_75t_R g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_23),
.B(n_36),
.C(n_28),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_35),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_25),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_31),
.B1(n_30),
.B2(n_37),
.Y(n_68)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_51),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_47),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_56),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_48),
.A2(n_36),
.B(n_25),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_46),
.C(n_44),
.Y(n_92)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_36),
.B1(n_24),
.B2(n_34),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_57),
.A2(n_68),
.B1(n_80),
.B2(n_82),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_58),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_28),
.B1(n_24),
.B2(n_34),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_63),
.B1(n_33),
.B2(n_38),
.Y(n_96)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_69),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_28),
.B1(n_24),
.B2(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_35),
.B1(n_25),
.B2(n_31),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_70),
.B1(n_74),
.B2(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_35),
.B1(n_37),
.B2(n_30),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_78),
.Y(n_91)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_75),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_27),
.B1(n_29),
.B2(n_22),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_82),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_29),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_79),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_21),
.B1(n_22),
.B2(n_26),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_21),
.B1(n_26),
.B2(n_19),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_98),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_20),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_52),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_106),
.C(n_53),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_56),
.A2(n_38),
.B1(n_18),
.B2(n_26),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_93),
.A2(n_102),
.B1(n_109),
.B2(n_110),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_96),
.A2(n_114),
.B1(n_117),
.B2(n_54),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_11),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_97),
.B(n_14),
.Y(n_134)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_38),
.B1(n_18),
.B2(n_11),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_66),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_104),
.B(n_113),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_19),
.C(n_18),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_107),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_75),
.A2(n_9),
.B1(n_17),
.B2(n_16),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_20),
.B1(n_8),
.B2(n_11),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_111),
.A2(n_120),
.B1(n_121),
.B2(n_51),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_80),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_71),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_77),
.A2(n_12),
.B1(n_4),
.B2(n_5),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_57),
.Y(n_123)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_138),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_127),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_142),
.B(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_139),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_95),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_131),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_119),
.B(n_111),
.C(n_114),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_132),
.A2(n_104),
.B(n_108),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_106),
.C(n_112),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_134),
.B(n_116),
.Y(n_172)
);

AO21x2_ASAP7_75t_L g135 ( 
.A1(n_87),
.A2(n_81),
.B(n_72),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_135),
.A2(n_148),
.B1(n_153),
.B2(n_147),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_95),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_136),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_118),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_137),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_53),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_90),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_141),
.Y(n_180)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_3),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_72),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_144),
.B(n_7),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_50),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_152),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_147),
.B(n_153),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_96),
.A2(n_76),
.B1(n_73),
.B2(n_60),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_120),
.A2(n_76),
.B1(n_51),
.B2(n_66),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_105),
.B1(n_107),
.B2(n_101),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_150),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_103),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_4),
.B(n_5),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_90),
.B(n_103),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_125),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_160),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_122),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_161),
.A2(n_182),
.B1(n_185),
.B2(n_135),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_94),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_165),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_145),
.A2(n_105),
.B1(n_101),
.B2(n_98),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_164),
.A2(n_176),
.B1(n_183),
.B2(n_166),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_94),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_179),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_167),
.A2(n_168),
.B(n_16),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_123),
.B(n_121),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_173),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_172),
.B(n_175),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_121),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_177),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_140),
.B(n_139),
.Y(n_175)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_132),
.A2(n_108),
.B1(n_116),
.B2(n_115),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_148),
.A2(n_115),
.B1(n_108),
.B2(n_14),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_6),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_188),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_135),
.A2(n_7),
.B1(n_14),
.B2(n_15),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_138),
.B(n_126),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_189),
.A2(n_201),
.B(n_208),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_177),
.A2(n_135),
.B1(n_186),
.B2(n_156),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_190),
.A2(n_197),
.B(n_211),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_152),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_196),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_193),
.B(n_183),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_167),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_204),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_143),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_142),
.B(n_124),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_157),
.A2(n_137),
.B1(n_154),
.B2(n_142),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_198),
.A2(n_203),
.B1(n_212),
.B2(n_185),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_159),
.A2(n_130),
.B(n_127),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_179),
.B(n_136),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_209),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_159),
.A2(n_144),
.B(n_146),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_175),
.B(n_15),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_184),
.B(n_15),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_210),
.B(n_214),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_187),
.A2(n_17),
.B1(n_173),
.B2(n_170),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_162),
.A2(n_17),
.B(n_165),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_213),
.A2(n_163),
.B(n_172),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_169),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_215),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_184),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_158),
.B(n_187),
.C(n_182),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_164),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_176),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_218),
.B(n_163),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_221),
.A2(n_223),
.B1(n_212),
.B2(n_194),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_203),
.A2(n_186),
.B1(n_161),
.B2(n_178),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_242),
.C(n_222),
.Y(n_260)
);

INVx13_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_230),
.Y(n_255)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_232),
.B(n_233),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_171),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_180),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_237),
.A2(n_240),
.B1(n_241),
.B2(n_191),
.Y(n_247)
);

NAND2xp33_ASAP7_75t_SL g238 ( 
.A(n_207),
.B(n_160),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_238),
.B(n_208),
.Y(n_258)
);

OA22x2_ASAP7_75t_L g239 ( 
.A1(n_193),
.A2(n_169),
.B1(n_181),
.B2(n_156),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_239),
.A2(n_207),
.B1(n_211),
.B2(n_202),
.Y(n_246)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_192),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_204),
.C(n_214),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_226),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_244),
.A2(n_252),
.B1(n_257),
.B2(n_233),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_246),
.A2(n_223),
.B1(n_219),
.B2(n_240),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_237),
.A2(n_217),
.B1(n_200),
.B2(n_198),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_254),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_196),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_213),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_258),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_221),
.A2(n_202),
.B1(n_197),
.B2(n_189),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_241),
.B(n_195),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_259),
.B(n_261),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_229),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_226),
.B(n_195),
.Y(n_261)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_262),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_265),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_277),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_228),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_236),
.B(n_234),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_268),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_257),
.A2(n_236),
.B1(n_219),
.B2(n_234),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_269),
.A2(n_271),
.B1(n_246),
.B2(n_252),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_274),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_239),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_222),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_288),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_228),
.C(n_231),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_289),
.C(n_290),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_273),
.A2(n_239),
.B1(n_244),
.B2(n_224),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_270),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_269),
.A2(n_239),
.B1(n_230),
.B2(n_224),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_286),
.B(n_287),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_254),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_258),
.C(n_201),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_253),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_268),
.B(n_239),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_297),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_256),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_296),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_291),
.B(n_275),
.Y(n_296)
);

FAx1_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_277),
.CI(n_272),
.CON(n_297),
.SN(n_297)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_285),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_263),
.C(n_278),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_290),
.Y(n_309)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_181),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_304),
.B(n_305),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_282),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_299),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_301),
.B(n_283),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_308),
.B(n_309),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_311),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_292),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_312),
.A2(n_302),
.A3(n_300),
.B1(n_294),
.B2(n_305),
.C1(n_306),
.C2(n_297),
.Y(n_316)
);

OAI21x1_ASAP7_75t_L g318 ( 
.A1(n_316),
.A2(n_317),
.B(n_238),
.Y(n_318)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_314),
.A2(n_297),
.A3(n_295),
.B1(n_299),
.B2(n_191),
.C1(n_209),
.C2(n_210),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_318),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_313),
.B(n_174),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_320),
.B(n_313),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_319),
.Y(n_322)
);


endmodule