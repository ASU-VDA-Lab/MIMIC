module fake_jpeg_11149_n_631 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_631);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_631;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_60),
.B(n_70),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_61),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_62),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_63),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_65),
.Y(n_164)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_67),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_68),
.Y(n_194)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_24),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_72),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_75),
.Y(n_198)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_77),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_20),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_78),
.B(n_80),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_79),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_24),
.B(n_18),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_81),
.Y(n_179)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_84),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g169 ( 
.A(n_87),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_88),
.Y(n_186)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_92),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_50),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_93),
.B(n_104),
.Y(n_180)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_96),
.Y(n_192)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_97),
.Y(n_175)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_102),
.Y(n_191)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_103),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_38),
.B(n_0),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_26),
.Y(n_107)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_107),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_108),
.Y(n_207)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

BUFx10_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_110),
.Y(n_213)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_26),
.Y(n_111)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

CKINVDCx6p67_ASAP7_75t_R g170 ( 
.A(n_112),
.Y(n_170)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_40),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_114),
.B(n_120),
.Y(n_185)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_38),
.Y(n_116)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_33),
.Y(n_118)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_118),
.Y(n_204)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_35),
.Y(n_119)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_119),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_46),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_121),
.B(n_56),
.Y(n_193)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_35),
.Y(n_122)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_43),
.Y(n_124)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_45),
.Y(n_125)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_125),
.Y(n_203)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_38),
.Y(n_126)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_126),
.Y(n_205)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_127),
.Y(n_212)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_48),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_128),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_40),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_129),
.B(n_167),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_78),
.B(n_46),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_130),
.B(n_142),
.Y(n_247)
);

BUFx2_ASAP7_75t_R g133 ( 
.A(n_60),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_133),
.B(n_187),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_71),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_L g281 ( 
.A(n_135),
.B(n_30),
.C(n_18),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_136),
.B(n_145),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_87),
.A2(n_27),
.B1(n_55),
.B2(n_58),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_141),
.A2(n_149),
.B1(n_162),
.B2(n_214),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_92),
.B(n_46),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_81),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_67),
.B(n_57),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_147),
.B(n_166),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_62),
.A2(n_27),
.B1(n_55),
.B2(n_56),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_84),
.A2(n_56),
.B1(n_41),
.B2(n_55),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_103),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_25),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_105),
.B(n_57),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_171),
.B(n_208),
.Y(n_231)
);

INVx4_ASAP7_75t_SL g187 ( 
.A(n_64),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_84),
.B(n_45),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_190),
.B(n_216),
.C(n_34),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

OA22x2_ASAP7_75t_L g197 ( 
.A1(n_127),
.A2(n_55),
.B1(n_27),
.B2(n_56),
.Y(n_197)
);

OA22x2_ASAP7_75t_SL g278 ( 
.A1(n_197),
.A2(n_199),
.B1(n_149),
.B2(n_141),
.Y(n_278)
);

OA22x2_ASAP7_75t_L g199 ( 
.A1(n_65),
.A2(n_27),
.B1(n_41),
.B2(n_52),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_61),
.B(n_22),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_201),
.B(n_47),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_118),
.B(n_54),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_68),
.B(n_22),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_211),
.B(n_44),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_72),
.A2(n_41),
.B1(n_53),
.B2(n_52),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_61),
.B(n_23),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_217),
.Y(n_296)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_218),
.Y(n_300)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_219),
.Y(n_292)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_138),
.Y(n_220)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_220),
.Y(n_302)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_221),
.Y(n_323)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_154),
.Y(n_222)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_222),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_79),
.B1(n_108),
.B2(n_96),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_223),
.A2(n_227),
.B1(n_230),
.B2(n_276),
.Y(n_307)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_152),
.Y(n_224)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_224),
.Y(n_348)
);

INVx11_ASAP7_75t_L g225 ( 
.A(n_137),
.Y(n_225)
);

BUFx8_ASAP7_75t_L g330 ( 
.A(n_225),
.Y(n_330)
);

INVx11_ASAP7_75t_L g226 ( 
.A(n_137),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_226),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_88),
.B1(n_77),
.B2(n_75),
.Y(n_227)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_165),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_229),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_143),
.A2(n_42),
.B1(n_25),
.B2(n_53),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_SL g232 ( 
.A1(n_190),
.A2(n_63),
.B(n_48),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_232),
.B(n_162),
.Y(n_312)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_173),
.Y(n_234)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_234),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_151),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_235),
.Y(n_329)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_236),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_180),
.A2(n_121),
.B1(n_23),
.B2(n_47),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_237),
.A2(n_266),
.B1(n_244),
.B2(n_258),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_151),
.Y(n_238)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_238),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_216),
.A2(n_63),
.B1(n_44),
.B2(n_54),
.Y(n_239)
);

AO21x1_ASAP7_75t_L g344 ( 
.A1(n_239),
.A2(n_266),
.B(n_277),
.Y(n_344)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_146),
.Y(n_240)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_240),
.Y(n_306)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_174),
.Y(n_241)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_241),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_185),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_242),
.B(n_252),
.Y(n_313)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_181),
.Y(n_243)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_243),
.Y(n_317)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_182),
.Y(n_245)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_245),
.Y(n_321)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_187),
.Y(n_246)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_246),
.Y(n_322)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_161),
.Y(n_248)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_248),
.Y(n_327)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_183),
.Y(n_249)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_249),
.Y(n_331)
);

INVx8_ASAP7_75t_L g250 ( 
.A(n_188),
.Y(n_250)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_250),
.Y(n_335)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_176),
.Y(n_251)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_251),
.Y(n_341)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_185),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_253),
.B(n_254),
.Y(n_314)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_150),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_159),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_255),
.A2(n_259),
.B1(n_272),
.B2(n_280),
.Y(n_347)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_256),
.B(n_261),
.Y(n_319)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_157),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_257),
.B(n_260),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_159),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_132),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_158),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_139),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_262),
.B(n_264),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_208),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_263),
.Y(n_345)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_140),
.Y(n_264)
);

CKINVDCx12_ASAP7_75t_R g265 ( 
.A(n_179),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_265),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_180),
.B(n_121),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_201),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_267),
.B(n_268),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_196),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_269),
.B(n_273),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_270),
.B(n_283),
.Y(n_295)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_184),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_271),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_164),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_156),
.B(n_42),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_275),
.B(n_281),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_202),
.A2(n_34),
.B1(n_54),
.B2(n_30),
.Y(n_276)
);

FAx1_ASAP7_75t_L g277 ( 
.A(n_130),
.B(n_48),
.CI(n_18),
.CON(n_277),
.SN(n_277)
);

OA22x2_ASAP7_75t_L g315 ( 
.A1(n_278),
.A2(n_197),
.B1(n_210),
.B2(n_200),
.Y(n_315)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_191),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_279),
.B(n_284),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_164),
.Y(n_280)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_148),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_282),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_156),
.B(n_17),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_203),
.Y(n_284)
);

INVx11_ASAP7_75t_L g285 ( 
.A(n_137),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_290),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_172),
.B(n_17),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_286),
.B(n_172),
.Y(n_311)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_209),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_287),
.B(n_289),
.Y(n_309)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_205),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_177),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_206),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_213),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_263),
.A2(n_147),
.B1(n_215),
.B2(n_178),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_294),
.A2(n_0),
.B(n_1),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_298),
.A2(n_318),
.B1(n_287),
.B2(n_271),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_233),
.B(n_142),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_301),
.B(n_339),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_223),
.A2(n_227),
.B1(n_278),
.B2(n_231),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_308),
.A2(n_324),
.B1(n_328),
.B2(n_337),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_311),
.B(n_304),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_312),
.B(n_315),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_288),
.A2(n_197),
.B1(n_169),
.B2(n_192),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_233),
.A2(n_171),
.B1(n_193),
.B2(n_169),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_247),
.A2(n_163),
.B1(n_198),
.B2(n_195),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_336),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_277),
.A2(n_207),
.B1(n_198),
.B2(n_195),
.Y(n_337)
);

OA22x2_ASAP7_75t_L g338 ( 
.A1(n_246),
.A2(n_144),
.B1(n_131),
.B2(n_194),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_338),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_228),
.B(n_30),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_244),
.B(n_189),
.C(n_170),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_170),
.C(n_272),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_274),
.B(n_155),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_346),
.B(n_281),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_319),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_350),
.B(n_371),
.Y(n_395)
);

NOR3xp33_ASAP7_75t_L g397 ( 
.A(n_351),
.B(n_370),
.C(n_394),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_352),
.A2(n_357),
.B1(n_355),
.B2(n_335),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_304),
.B(n_256),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_353),
.B(n_356),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_324),
.A2(n_250),
.B1(n_218),
.B2(n_268),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_354),
.A2(n_380),
.B1(n_347),
.B2(n_303),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_318),
.A2(n_194),
.B1(n_252),
.B2(n_249),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_292),
.Y(n_358)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_358),
.Y(n_408)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_292),
.Y(n_361)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_361),
.Y(n_403)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_362),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_325),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_363),
.B(n_377),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_301),
.B(n_241),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_364),
.B(n_382),
.Y(n_406)
);

INVx13_ASAP7_75t_L g365 ( 
.A(n_300),
.Y(n_365)
);

INVxp33_ASAP7_75t_L g421 ( 
.A(n_365),
.Y(n_421)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_296),
.Y(n_366)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_366),
.Y(n_420)
);

INVx13_ASAP7_75t_L g367 ( 
.A(n_300),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_367),
.Y(n_413)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_296),
.Y(n_368)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_368),
.Y(n_411)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_302),
.Y(n_369)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_369),
.Y(n_414)
);

AOI32xp33_ASAP7_75t_L g370 ( 
.A1(n_312),
.A2(n_226),
.A3(n_225),
.B1(n_285),
.B2(n_221),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_319),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_372),
.B(n_393),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_326),
.A2(n_170),
.B(n_221),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_373),
.A2(n_379),
.B(n_390),
.Y(n_422)
);

INVx8_ASAP7_75t_L g375 ( 
.A(n_329),
.Y(n_375)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_375),
.Y(n_400)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_302),
.Y(n_376)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_320),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_348),
.Y(n_378)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_378),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_344),
.A2(n_153),
.B(n_160),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_335),
.A2(n_160),
.B1(n_153),
.B2(n_255),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_329),
.Y(n_381)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_381),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_313),
.B(n_280),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_305),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_383),
.B(n_384),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_305),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_385),
.B(n_387),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_333),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_386),
.B(n_388),
.Y(n_412)
);

INVx5_ASAP7_75t_SL g387 ( 
.A(n_330),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_314),
.B(n_259),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_349),
.B(n_238),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_389),
.B(n_340),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_344),
.A2(n_2),
.B(n_3),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_345),
.A2(n_235),
.B1(n_17),
.B2(n_16),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_391),
.A2(n_339),
.B(n_334),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_298),
.B(n_16),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_295),
.B(n_14),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_359),
.A2(n_307),
.B1(n_328),
.B2(n_315),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_396),
.A2(n_423),
.B(n_429),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_360),
.B(n_342),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_398),
.B(n_418),
.C(n_431),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_402),
.A2(n_391),
.B(n_389),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_364),
.B(n_338),
.Y(n_404)
);

AO21x1_ASAP7_75t_L g461 ( 
.A1(n_404),
.A2(n_425),
.B(n_322),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_374),
.A2(n_315),
.B1(n_326),
.B2(n_346),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_409),
.B(n_426),
.Y(n_453)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_410),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_360),
.B(n_294),
.Y(n_418)
);

AO22x1_ASAP7_75t_L g423 ( 
.A1(n_355),
.A2(n_315),
.B1(n_338),
.B2(n_327),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_388),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_424),
.B(n_377),
.Y(n_434)
);

O2A1O1Ixp33_ASAP7_75t_L g425 ( 
.A1(n_359),
.A2(n_338),
.B(n_319),
.C(n_322),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_374),
.A2(n_334),
.B1(n_336),
.B2(n_293),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_427),
.B(n_428),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_386),
.B(n_309),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_382),
.B(n_340),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_430),
.B(n_363),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_359),
.B(n_299),
.Y(n_431)
);

INVx13_ASAP7_75t_L g433 ( 
.A(n_421),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_433),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_434),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_396),
.A2(n_392),
.B1(n_379),
.B2(n_390),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_435),
.A2(n_450),
.B1(n_459),
.B2(n_404),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_401),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_436),
.B(n_443),
.Y(n_472)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_438),
.Y(n_477)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_411),
.Y(n_441)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_441),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_428),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_432),
.B(n_356),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_444),
.B(n_448),
.Y(n_494)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_411),
.Y(n_445)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_445),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_426),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_446),
.B(n_452),
.Y(n_479)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_408),
.Y(n_447)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_447),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_412),
.B(n_341),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_431),
.B(n_385),
.Y(n_449)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_449),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_410),
.A2(n_392),
.B1(n_357),
.B2(n_373),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_451),
.A2(n_461),
.B1(n_422),
.B2(n_446),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_412),
.B(n_341),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_306),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_454),
.B(n_465),
.Y(n_486)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_414),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_455),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_456),
.B(n_462),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_398),
.B(n_372),
.C(n_393),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_464),
.C(n_415),
.Y(n_473)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_414),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_458),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_406),
.A2(n_368),
.B1(n_366),
.B2(n_369),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_SL g460 ( 
.A(n_399),
.B(n_387),
.C(n_376),
.Y(n_460)
);

FAx1_ASAP7_75t_SL g491 ( 
.A(n_460),
.B(n_367),
.CI(n_365),
.CON(n_491),
.SN(n_491)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_416),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_430),
.B(n_358),
.Y(n_463)
);

OAI21xp33_ASAP7_75t_L g483 ( 
.A1(n_463),
.A2(n_467),
.B(n_403),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_418),
.B(n_306),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_413),
.B(n_327),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_416),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_466),
.B(n_417),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_406),
.B(n_361),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_439),
.A2(n_422),
.B1(n_429),
.B2(n_404),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_469),
.A2(n_488),
.B1(n_435),
.B2(n_461),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_470),
.A2(n_476),
.B1(n_493),
.B2(n_405),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_442),
.B(n_415),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_471),
.B(n_489),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_473),
.B(n_449),
.C(n_440),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_456),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_474),
.B(n_485),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_475),
.A2(n_451),
.B1(n_455),
.B2(n_441),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_439),
.A2(n_404),
.B1(n_425),
.B2(n_399),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_453),
.A2(n_399),
.B(n_395),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_478),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_436),
.A2(n_397),
.B1(n_423),
.B2(n_420),
.Y(n_480)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_480),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_483),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_453),
.A2(n_423),
.B(n_407),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_461),
.A2(n_419),
.B1(n_400),
.B2(n_417),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_442),
.B(n_316),
.Y(n_489)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_490),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_459),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_450),
.A2(n_400),
.B1(n_419),
.B2(n_405),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_443),
.B(n_343),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_496),
.B(n_500),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_464),
.B(n_457),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_497),
.B(n_317),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_440),
.B(n_343),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_472),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_502),
.B(n_521),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_504),
.B(n_507),
.C(n_508),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_489),
.B(n_449),
.C(n_437),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_471),
.B(n_437),
.C(n_460),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_509),
.A2(n_514),
.B1(n_518),
.B2(n_476),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_510),
.A2(n_491),
.B(n_490),
.Y(n_535)
);

NAND2xp67_ASAP7_75t_SL g512 ( 
.A(n_485),
.B(n_467),
.Y(n_512)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_512),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_SL g513 ( 
.A1(n_499),
.A2(n_466),
.B1(n_462),
.B2(n_458),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_513),
.A2(n_477),
.B1(n_433),
.B2(n_384),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_492),
.B(n_463),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g544 ( 
.A(n_515),
.B(n_527),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_473),
.B(n_445),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_516),
.B(n_526),
.Y(n_550)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_472),
.Y(n_517)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_517),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_469),
.A2(n_447),
.B1(n_438),
.B2(n_403),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_519),
.B(n_529),
.C(n_498),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_486),
.B(n_362),
.Y(n_521)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_495),
.Y(n_523)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_523),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_524),
.A2(n_488),
.B1(n_481),
.B2(n_498),
.Y(n_530)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_495),
.Y(n_525)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_525),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_497),
.B(n_378),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_478),
.B(n_317),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_479),
.B(n_421),
.Y(n_528)
);

CKINVDCx14_ASAP7_75t_R g541 ( 
.A(n_528),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_492),
.B(n_321),
.C(n_303),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_530),
.A2(n_518),
.B1(n_512),
.B2(n_529),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_506),
.B(n_481),
.Y(n_532)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_532),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_534),
.B(n_543),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_535),
.A2(n_507),
.B(n_504),
.Y(n_555)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_536),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_516),
.B(n_493),
.C(n_470),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_537),
.B(n_540),
.Y(n_564)
);

XNOR2x1_ASAP7_75t_L g538 ( 
.A(n_508),
.B(n_491),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_538),
.B(n_310),
.Y(n_572)
);

AOI21xp33_ASAP7_75t_L g540 ( 
.A1(n_522),
.A2(n_484),
.B(n_482),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_520),
.B(n_484),
.Y(n_542)
);

CKINVDCx14_ASAP7_75t_R g559 ( 
.A(n_542),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_522),
.A2(n_482),
.B1(n_468),
.B2(n_487),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_514),
.A2(n_509),
.B1(n_503),
.B2(n_510),
.Y(n_545)
);

INVxp33_ASAP7_75t_SL g563 ( 
.A(n_545),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_511),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_546),
.B(n_549),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_501),
.B(n_487),
.C(n_468),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_552),
.B(n_433),
.Y(n_566)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_505),
.Y(n_553)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_553),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_554),
.A2(n_545),
.B1(n_536),
.B2(n_547),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_555),
.A2(n_565),
.B(n_535),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_548),
.B(n_526),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_556),
.B(n_560),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_549),
.B(n_501),
.C(n_519),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_542),
.B(n_527),
.Y(n_562)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_562),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_SL g565 ( 
.A1(n_531),
.A2(n_515),
.B(n_477),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_566),
.B(n_572),
.Y(n_586)
);

CKINVDCx14_ASAP7_75t_R g568 ( 
.A(n_532),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_568),
.B(n_551),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_541),
.B(n_553),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_569),
.B(n_571),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_533),
.B(n_323),
.C(n_321),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_533),
.B(n_375),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_573),
.B(n_534),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_567),
.B(n_537),
.Y(n_574)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_574),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_575),
.A2(n_587),
.B1(n_559),
.B2(n_557),
.Y(n_597)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_576),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_571),
.B(n_550),
.C(n_530),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_577),
.B(n_580),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_560),
.B(n_561),
.C(n_564),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_555),
.B(n_550),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_581),
.B(n_584),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_582),
.B(n_565),
.Y(n_596)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_558),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_583),
.B(n_585),
.Y(n_592)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_558),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_561),
.A2(n_543),
.B(n_551),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_563),
.B(n_538),
.C(n_544),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_589),
.B(n_590),
.C(n_562),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_570),
.B(n_544),
.C(n_539),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_591),
.B(n_596),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_577),
.B(n_570),
.C(n_566),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_593),
.B(n_594),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_574),
.B(n_572),
.C(n_557),
.Y(n_594)
);

INVx6_ASAP7_75t_L g595 ( 
.A(n_588),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_595),
.B(n_580),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_597),
.B(n_575),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_578),
.B(n_539),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_599),
.A2(n_600),
.B(n_586),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_590),
.B(n_381),
.Y(n_600)
);

OAI21x1_ASAP7_75t_SL g614 ( 
.A1(n_604),
.A2(n_608),
.B(n_592),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_605),
.B(n_607),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_603),
.B(n_579),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_606),
.B(n_611),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_SL g607 ( 
.A1(n_601),
.A2(n_589),
.B1(n_586),
.B2(n_383),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_591),
.B(n_331),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_610),
.B(n_613),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_602),
.B(n_331),
.C(n_310),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_598),
.B(n_593),
.C(n_594),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_614),
.A2(n_607),
.B(n_610),
.Y(n_621)
);

AOI322xp5_ASAP7_75t_L g616 ( 
.A1(n_609),
.A2(n_595),
.A3(n_596),
.B1(n_323),
.B2(n_330),
.C1(n_332),
.C2(n_297),
.Y(n_616)
);

OAI321xp33_ASAP7_75t_L g623 ( 
.A1(n_616),
.A2(n_330),
.A3(n_14),
.B1(n_4),
.B2(n_6),
.C(n_8),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_605),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_618),
.B(n_619),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_612),
.B(n_332),
.Y(n_619)
);

AOI31xp67_ASAP7_75t_SL g625 ( 
.A1(n_621),
.A2(n_623),
.A3(n_2),
.B(n_3),
.Y(n_625)
);

AOI21xp33_ASAP7_75t_L g622 ( 
.A1(n_617),
.A2(n_615),
.B(n_620),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_622),
.B(n_624),
.Y(n_626)
);

OAI21x1_ASAP7_75t_SL g627 ( 
.A1(n_625),
.A2(n_626),
.B(n_4),
.Y(n_627)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_627),
.B(n_8),
.Y(n_628)
);

OAI221xp5_ASAP7_75t_L g629 ( 
.A1(n_628),
.A2(n_10),
.B1(n_12),
.B2(n_297),
.C(n_583),
.Y(n_629)
);

XOR2xp5_ASAP7_75t_L g630 ( 
.A(n_629),
.B(n_10),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_630),
.B(n_12),
.Y(n_631)
);


endmodule