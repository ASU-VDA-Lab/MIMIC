module fake_jpeg_3468_n_180 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_180);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_63),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_18),
.C(n_36),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_48),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_66),
.A2(n_65),
.B1(n_60),
.B2(n_58),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

CKINVDCx9p33_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_57),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_58),
.B1(n_42),
.B2(n_53),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_54),
.B1(n_56),
.B2(n_50),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_42),
.B1(n_46),
.B2(n_48),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_79),
.A2(n_56),
.B(n_62),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_91),
.Y(n_104)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g103 ( 
.A(n_83),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_68),
.B(n_64),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_84),
.Y(n_111)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_49),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_73),
.B(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_74),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_55),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_69),
.B1(n_50),
.B2(n_3),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_97),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_112),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_69),
.B1(n_54),
.B2(n_49),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_102),
.B1(n_3),
.B2(n_4),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_1),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_119),
.Y(n_133)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_21),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_SL g150 ( 
.A(n_117),
.B(n_16),
.C(n_17),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_2),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_87),
.B1(n_86),
.B2(n_5),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_123),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

OA21x2_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_87),
.B(n_4),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_11),
.B(n_12),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_131),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_7),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_24),
.C(n_34),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_145),
.C(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_130),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_146),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_121),
.C(n_128),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_9),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_114),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_150),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_12),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_149),
.B(n_19),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_142),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_154),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_133),
.B(n_22),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_145),
.B(n_26),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_140),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_29),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_134),
.B(n_27),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_28),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_139),
.B1(n_141),
.B2(n_144),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_166),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_168),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_136),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_153),
.A2(n_148),
.B(n_135),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_167),
.Y(n_172)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_152),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_174),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_160),
.B(n_155),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_163),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_171),
.B(n_164),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_172),
.B(n_160),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_30),
.B(n_32),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_33),
.Y(n_180)
);


endmodule