module fake_jpeg_16166_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_43),
.Y(n_58)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_22),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_18),
.Y(n_60)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_26),
.B1(n_24),
.B2(n_30),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_46),
.A2(n_19),
.B1(n_17),
.B2(n_27),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_48),
.B(n_55),
.Y(n_81)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_40),
.Y(n_50)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_60),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_30),
.Y(n_55)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_44),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_26),
.B1(n_29),
.B2(n_21),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_44),
.B1(n_29),
.B2(n_38),
.Y(n_80)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_35),
.Y(n_88)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_26),
.B1(n_39),
.B2(n_42),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_71),
.A2(n_82),
.B1(n_86),
.B2(n_49),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_42),
.B1(n_41),
.B2(n_32),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_72),
.A2(n_74),
.B1(n_65),
.B2(n_53),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_42),
.B1(n_32),
.B2(n_23),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_76),
.B(n_84),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_58),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_79),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_80),
.A2(n_94),
.B1(n_27),
.B2(n_17),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_43),
.B1(n_38),
.B2(n_32),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_61),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_43),
.B1(n_32),
.B2(n_23),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_68),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_52),
.B(n_22),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_95),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_47),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_59),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_103),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_50),
.B(n_35),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_69),
.B(n_31),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_70),
.B(n_81),
.C(n_83),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_51),
.B1(n_54),
.B2(n_57),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_77),
.B1(n_69),
.B2(n_96),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_54),
.B1(n_51),
.B2(n_18),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_9),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_119),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_78),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_110),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_114),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_122),
.B1(n_16),
.B2(n_86),
.Y(n_140)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_120),
.B1(n_125),
.B2(n_72),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_59),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_71),
.A2(n_67),
.B1(n_35),
.B2(n_28),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_80),
.A2(n_67),
.B1(n_21),
.B2(n_19),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_74),
.A2(n_35),
.B1(n_28),
.B2(n_36),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_104),
.B(n_90),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_139),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_16),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_135),
.B(n_148),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_140),
.B1(n_144),
.B2(n_145),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_104),
.B(n_95),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_142),
.A2(n_143),
.B(n_151),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_101),
.A2(n_69),
.B1(n_96),
.B2(n_91),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_123),
.A2(n_77),
.B1(n_85),
.B2(n_73),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_85),
.B1(n_73),
.B2(n_77),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_36),
.C(n_93),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_31),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_28),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_36),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_102),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_93),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_150),
.B(n_122),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_109),
.A2(n_33),
.B1(n_25),
.B2(n_2),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_152),
.A2(n_107),
.B1(n_120),
.B2(n_116),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_117),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_165),
.Y(n_181)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_156),
.B(n_158),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_128),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_159),
.A2(n_172),
.B1(n_145),
.B2(n_129),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_133),
.A2(n_101),
.B1(n_119),
.B2(n_115),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_111),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_171),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_167),
.A2(n_170),
.B(n_142),
.Y(n_184)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_105),
.Y(n_169)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

AOI322xp5_ASAP7_75t_L g170 ( 
.A1(n_127),
.A2(n_114),
.A3(n_125),
.B1(n_33),
.B2(n_126),
.C1(n_121),
.C2(n_124),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_113),
.A3(n_126),
.B1(n_98),
.B2(n_100),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_133),
.A2(n_100),
.B1(n_126),
.B2(n_116),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_132),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_175),
.Y(n_201)
);

OA21x2_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_25),
.B(n_33),
.Y(n_174)
);

AO22x1_ASAP7_75t_SL g187 ( 
.A1(n_174),
.A2(n_176),
.B1(n_152),
.B2(n_136),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_150),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g176 ( 
.A1(n_141),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_178),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_178),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_182),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_164),
.B1(n_167),
.B2(n_151),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_183),
.A2(n_184),
.B1(n_187),
.B2(n_191),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_154),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_189),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_188),
.A2(n_195),
.B1(n_176),
.B2(n_159),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_162),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_129),
.B(n_147),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_163),
.A2(n_151),
.B(n_139),
.Y(n_194)
);

AOI21xp33_ASAP7_75t_L g229 ( 
.A1(n_194),
.A2(n_204),
.B(n_157),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_171),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_146),
.C(n_137),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_199),
.C(n_173),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_151),
.B(n_143),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_203),
.B1(n_174),
.B2(n_176),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_146),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_134),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_164),
.A2(n_175),
.B1(n_169),
.B2(n_161),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_160),
.A2(n_148),
.B(n_135),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_153),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_211),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_228),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_203),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_213),
.C(n_218),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_171),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_166),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_227),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_216),
.B(n_187),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_217),
.A2(n_221),
.B1(n_223),
.B2(n_179),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_158),
.C(n_156),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_190),
.A2(n_176),
.B1(n_170),
.B2(n_140),
.Y(n_220)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_190),
.B1(n_185),
.B2(n_205),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_183),
.C(n_200),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_224),
.C(n_226),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_205),
.A2(n_172),
.B1(n_174),
.B2(n_165),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_174),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_225),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_204),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_181),
.B(n_157),
.C(n_144),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_SL g233 ( 
.A(n_229),
.B(n_187),
.C(n_196),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_210),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_251),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_236),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_226),
.B(n_219),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_241),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_213),
.B(n_186),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_218),
.A2(n_192),
.B1(n_189),
.B2(n_179),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_237),
.A2(n_243),
.B1(n_0),
.B2(n_1),
.Y(n_257)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_223),
.A2(n_202),
.B(n_196),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_240),
.A2(n_237),
.B(n_243),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_202),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_209),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_224),
.C(n_13),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_180),
.B1(n_138),
.B2(n_2),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_15),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_250),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_14),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_14),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_208),
.B1(n_211),
.B2(n_215),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_253),
.A2(n_261),
.B1(n_265),
.B2(n_269),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_10),
.C(n_11),
.Y(n_284)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_257),
.Y(n_282)
);

O2A1O1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_260),
.A2(n_4),
.B(n_6),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_234),
.A2(n_232),
.B1(n_230),
.B2(n_248),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_262),
.A2(n_247),
.B(n_242),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_1),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_264),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_3),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_249),
.B1(n_236),
.B2(n_247),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_270),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_274),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_264),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_275),
.A2(n_253),
.B(n_262),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_255),
.Y(n_276)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_244),
.B1(n_5),
.B2(n_6),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_277),
.A2(n_279),
.B1(n_284),
.B2(n_258),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_244),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_258),
.C(n_12),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_263),
.B(n_273),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_261),
.B(n_9),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_260),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_254),
.B(n_10),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_283),
.B(n_284),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_288),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_286),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_267),
.Y(n_288)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_267),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_297),
.C(n_12),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_257),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_293),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_266),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_296),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_269),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_298),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_281),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_304),
.C(n_308),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_294),
.A2(n_277),
.B1(n_8),
.B2(n_7),
.Y(n_303)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_303),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_285),
.A2(n_12),
.B(n_13),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_7),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_291),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_306),
.A2(n_287),
.B1(n_290),
.B2(n_297),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_313),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_298),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_288),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_316),
.Y(n_323)
);

OR2x6_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_13),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_7),
.B(n_8),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_309),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_7),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_304),
.C(n_305),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_315),
.Y(n_319)
);

OAI21x1_ASAP7_75t_SL g326 ( 
.A1(n_319),
.A2(n_320),
.B(n_321),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_323),
.A2(n_302),
.B(n_315),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_310),
.C(n_324),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

AOI32xp33_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_322),
.A3(n_326),
.B1(n_301),
.B2(n_300),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_318),
.Y(n_330)
);


endmodule