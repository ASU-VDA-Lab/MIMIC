module fake_ariane_781_n_1858 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_543, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_558, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_531, n_1858);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_558;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;
input n_531;

output n_1858;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_1383;
wire n_603;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_1853;
wire n_764;
wire n_1503;
wire n_1196;
wire n_1181;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_813;
wire n_995;
wire n_1184;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_1751;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1716;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_1819;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_632;
wire n_650;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1674;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_670;
wire n_1826;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1467;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_604;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_1726;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_887;
wire n_729;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_1156;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_1402;
wire n_957;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_1005;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_1708;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_832;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_1854;
wire n_666;
wire n_1747;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_805;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_1137;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1208;
wire n_802;
wire n_1151;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_748;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_576;
wire n_843;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_673;
wire n_1038;
wire n_571;
wire n_1521;
wire n_1694;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_1166;
wire n_1056;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_1789;
wire n_763;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_621;
wire n_1587;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_1679;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_917;
wire n_1271;
wire n_1530;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_1813;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1344;
wire n_1390;
wire n_1792;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_904;
wire n_1696;
wire n_1059;
wire n_684;
wire n_1039;
wire n_1150;
wire n_977;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_1063;
wire n_991;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_1126;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_946;
wire n_757;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_937;
wire n_1474;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_1434;
wire n_1569;
wire n_1662;
wire n_1299;
wire n_782;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_849;
wire n_1820;
wire n_1251;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_573;
wire n_796;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_282),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_119),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_531),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_533),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_413),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_483),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_477),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_414),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_302),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_463),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_507),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_361),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_545),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_468),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_474),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_557),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_45),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_522),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_315),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_526),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_141),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_503),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_24),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_540),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_524),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_115),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_319),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_491),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_146),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_559),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_255),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_46),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_550),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_365),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_80),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_389),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_549),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_363),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_515),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_362),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_269),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_539),
.Y(n_601)
);

BUFx10_ASAP7_75t_L g602 ( 
.A(n_223),
.Y(n_602)
);

BUFx5_ASAP7_75t_L g603 ( 
.A(n_516),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_520),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_354),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_355),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_525),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_95),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_270),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_489),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_490),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_498),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_558),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_466),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_122),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_450),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_312),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_18),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_91),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_50),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_209),
.Y(n_621)
);

BUFx5_ASAP7_75t_L g622 ( 
.A(n_227),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_128),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_453),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_396),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_3),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_324),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_231),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_514),
.Y(n_629)
);

BUFx8_ASAP7_75t_SL g630 ( 
.A(n_187),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_102),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_215),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_178),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_298),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_118),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_145),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_94),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_118),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_39),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_84),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_494),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_554),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_282),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_242),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_510),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_470),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_197),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_504),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_497),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_521),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_480),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_467),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_20),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_190),
.Y(n_654)
);

BUFx10_ASAP7_75t_L g655 ( 
.A(n_293),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_348),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_374),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_543),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_523),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_415),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_383),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_328),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_148),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_186),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_541),
.Y(n_665)
);

BUFx10_ASAP7_75t_L g666 ( 
.A(n_551),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_127),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_418),
.Y(n_668)
);

CKINVDCx14_ASAP7_75t_R g669 ( 
.A(n_333),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_127),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_500),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_204),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_339),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_534),
.Y(n_674)
);

CKINVDCx16_ASAP7_75t_R g675 ( 
.A(n_82),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_335),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_381),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_517),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_495),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_86),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_41),
.Y(n_681)
);

CKINVDCx16_ASAP7_75t_R g682 ( 
.A(n_139),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_511),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_488),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_536),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_320),
.Y(n_686)
);

BUFx10_ASAP7_75t_L g687 ( 
.A(n_260),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_49),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_409),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_221),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_464),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_230),
.Y(n_692)
);

CKINVDCx16_ASAP7_75t_R g693 ( 
.A(n_513),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_538),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_155),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_179),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_258),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_125),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_532),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_60),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_528),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_527),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_492),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_116),
.Y(n_704)
);

CKINVDCx14_ASAP7_75t_R g705 ( 
.A(n_486),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_281),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_519),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_499),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_87),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_461),
.Y(n_710)
);

BUFx10_ASAP7_75t_L g711 ( 
.A(n_493),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_509),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_518),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_150),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_395),
.Y(n_715)
);

BUFx10_ASAP7_75t_L g716 ( 
.A(n_471),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_473),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_512),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_535),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_555),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_68),
.Y(n_721)
);

INVxp67_ASAP7_75t_SL g722 ( 
.A(n_196),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_151),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_113),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_484),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_347),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_546),
.Y(n_727)
);

BUFx10_ASAP7_75t_L g728 ( 
.A(n_478),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_482),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_505),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_176),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_530),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_29),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_508),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_553),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_496),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_292),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_387),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_506),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_529),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_188),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_175),
.Y(n_742)
);

BUFx5_ASAP7_75t_L g743 ( 
.A(n_277),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_401),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_537),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_544),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_481),
.Y(n_747)
);

BUFx5_ASAP7_75t_L g748 ( 
.A(n_501),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_547),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_218),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_161),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_476),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_487),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_458),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_542),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_465),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_280),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_438),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_94),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_126),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_556),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_399),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_154),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_502),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_552),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_343),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_48),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_448),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_469),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_257),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_344),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_485),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_462),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_265),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_29),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_13),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_548),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_19),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_84),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_239),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_108),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_39),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_136),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_168),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_263),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_261),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_197),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_43),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_472),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_114),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_128),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_675),
.B(n_0),
.Y(n_792)
);

CKINVDCx14_ASAP7_75t_R g793 ( 
.A(n_669),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_622),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_622),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_R g796 ( 
.A(n_573),
.B(n_284),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_682),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_630),
.Y(n_798)
);

NOR2xp67_ASAP7_75t_L g799 ( 
.A(n_637),
.B(n_0),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_622),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_566),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_622),
.Y(n_802)
);

INVxp67_ASAP7_75t_SL g803 ( 
.A(n_791),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_567),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_743),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_576),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_577),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_743),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_612),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_743),
.Y(n_810)
);

INVxp67_ASAP7_75t_SL g811 ( 
.A(n_780),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_743),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_743),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_582),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_649),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_614),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_609),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_615),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_794),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_816),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_793),
.B(n_693),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_795),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_800),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_811),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_802),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_805),
.B(n_564),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_808),
.B(n_565),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_810),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_812),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_813),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_797),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_814),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_803),
.B(n_570),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_817),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_803),
.B(n_574),
.Y(n_835)
);

OA21x2_ASAP7_75t_L g836 ( 
.A1(n_818),
.A2(n_596),
.B(n_587),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_806),
.B(n_705),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_792),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_806),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_801),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_799),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_804),
.Y(n_842)
);

OA21x2_ASAP7_75t_L g843 ( 
.A1(n_796),
.A2(n_604),
.B(n_599),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_809),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_815),
.B(n_655),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_798),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_831),
.B(n_618),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_820),
.Y(n_848)
);

OR2x6_ASAP7_75t_L g849 ( 
.A(n_840),
.B(n_653),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_831),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_828),
.B(n_659),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_838),
.B(n_807),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_846),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_829),
.B(n_830),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_832),
.Y(n_855)
);

NOR2x1p5_ASAP7_75t_L g856 ( 
.A(n_846),
.B(n_722),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_839),
.B(n_684),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_819),
.Y(n_858)
);

AND2x2_ASAP7_75t_SL g859 ( 
.A(n_840),
.B(n_844),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_819),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_822),
.B(n_715),
.Y(n_861)
);

INVx8_ASAP7_75t_L g862 ( 
.A(n_845),
.Y(n_862)
);

INVx5_ASAP7_75t_L g863 ( 
.A(n_842),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_841),
.B(n_713),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_833),
.B(n_670),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_821),
.B(n_560),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_824),
.B(n_606),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_832),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_834),
.Y(n_869)
);

INVxp67_ASAP7_75t_SL g870 ( 
.A(n_826),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_835),
.B(n_823),
.Y(n_871)
);

OR2x6_ASAP7_75t_L g872 ( 
.A(n_827),
.B(n_608),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_825),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_843),
.A2(n_741),
.B1(n_776),
.B2(n_700),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_843),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_836),
.B(n_602),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_820),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_837),
.B(n_561),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_837),
.B(n_673),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_832),
.Y(n_880)
);

BUFx6f_ASAP7_75t_SL g881 ( 
.A(n_846),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_837),
.B(n_702),
.Y(n_882)
);

BUFx10_ASAP7_75t_L g883 ( 
.A(n_846),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_855),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_868),
.Y(n_885)
);

AO22x2_ASAP7_75t_L g886 ( 
.A1(n_847),
.A2(n_770),
.B1(n_785),
.B2(n_709),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_850),
.Y(n_887)
);

NAND2xp33_ASAP7_75t_L g888 ( 
.A(n_862),
.B(n_580),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_870),
.A2(n_752),
.B1(n_744),
.B2(n_588),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_873),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_852),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_880),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_871),
.B(n_780),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_854),
.A2(n_590),
.B1(n_591),
.B2(n_585),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_869),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_883),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_853),
.B(n_619),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_858),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_858),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_860),
.Y(n_900)
);

AO22x2_ASAP7_75t_L g901 ( 
.A1(n_857),
.A2(n_697),
.B1(n_698),
.B2(n_667),
.Y(n_901)
);

NOR2xp67_ASAP7_75t_L g902 ( 
.A(n_863),
.B(n_718),
.Y(n_902)
);

AO22x2_ASAP7_75t_L g903 ( 
.A1(n_864),
.A2(n_723),
.B1(n_628),
.B2(n_632),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_881),
.Y(n_904)
);

AO22x2_ASAP7_75t_L g905 ( 
.A1(n_878),
.A2(n_631),
.B1(n_644),
.B2(n_635),
.Y(n_905)
);

OAI221xp5_ASAP7_75t_L g906 ( 
.A1(n_867),
.A2(n_690),
.B1(n_692),
.B2(n_681),
.C(n_664),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_862),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_860),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_859),
.B(n_602),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_875),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_861),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_851),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_849),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_866),
.B(n_848),
.Y(n_914)
);

NOR2xp67_ASAP7_75t_L g915 ( 
.A(n_863),
.B(n_624),
.Y(n_915)
);

BUFx8_ASAP7_75t_L g916 ( 
.A(n_856),
.Y(n_916)
);

BUFx8_ASAP7_75t_L g917 ( 
.A(n_849),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_877),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_872),
.B(n_687),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_879),
.B(n_782),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_882),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_874),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_855),
.Y(n_923)
);

NAND2x1p5_ASAP7_75t_L g924 ( 
.A(n_853),
.B(n_757),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_855),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_870),
.B(n_780),
.Y(n_926)
);

OAI221xp5_ASAP7_75t_L g927 ( 
.A1(n_865),
.A2(n_786),
.B1(n_787),
.B2(n_778),
.C(n_774),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_855),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_870),
.B(n_788),
.Y(n_929)
);

NAND2x1p5_ASAP7_75t_L g930 ( 
.A(n_853),
.B(n_648),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_850),
.B(n_687),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_855),
.Y(n_932)
);

NOR2xp67_ASAP7_75t_L g933 ( 
.A(n_863),
.B(n_627),
.Y(n_933)
);

AO22x2_ASAP7_75t_L g934 ( 
.A1(n_847),
.A2(n_645),
.B1(n_679),
.B2(n_629),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_855),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_853),
.B(n_594),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_881),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_855),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_881),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_850),
.B(n_600),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_855),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_870),
.B(n_788),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_870),
.B(n_788),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_870),
.A2(n_650),
.B1(n_651),
.B2(n_646),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_870),
.A2(n_621),
.B1(n_623),
.B2(n_620),
.Y(n_945)
);

OR2x6_ASAP7_75t_L g946 ( 
.A(n_853),
.B(n_671),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_850),
.B(n_626),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_873),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_855),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_873),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_850),
.B(n_633),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_855),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_873),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_881),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_855),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_876),
.A2(n_666),
.B1(n_711),
.B2(n_655),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_883),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_855),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_873),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_883),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_855),
.Y(n_961)
);

AO22x2_ASAP7_75t_L g962 ( 
.A1(n_847),
.A2(n_737),
.B1(n_730),
.B2(n_668),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_870),
.B(n_783),
.Y(n_963)
);

NAND2x1p5_ASAP7_75t_L g964 ( 
.A(n_853),
.B(n_755),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_873),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_873),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_855),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_855),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_883),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_855),
.Y(n_970)
);

OAI221xp5_ASAP7_75t_L g971 ( 
.A1(n_865),
.A2(n_639),
.B1(n_640),
.B2(n_638),
.C(n_636),
.Y(n_971)
);

NOR2xp67_ASAP7_75t_L g972 ( 
.A(n_863),
.B(n_660),
.Y(n_972)
);

NOR2xp67_ASAP7_75t_L g973 ( 
.A(n_863),
.B(n_694),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_853),
.B(n_643),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_912),
.B(n_647),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_969),
.B(n_654),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_969),
.B(n_663),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_963),
.B(n_672),
.Y(n_978)
);

NAND2xp33_ASAP7_75t_SL g979 ( 
.A(n_896),
.B(n_680),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_887),
.B(n_688),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_921),
.B(n_695),
.Y(n_981)
);

NAND2xp33_ASAP7_75t_SL g982 ( 
.A(n_957),
.B(n_696),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_911),
.B(n_704),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_909),
.B(n_701),
.Y(n_984)
);

NAND2xp33_ASAP7_75t_SL g985 ( 
.A(n_960),
.B(n_706),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_891),
.B(n_714),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_914),
.B(n_721),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_889),
.B(n_944),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_892),
.B(n_724),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_920),
.B(n_731),
.Y(n_990)
);

NAND2xp33_ASAP7_75t_SL g991 ( 
.A(n_918),
.B(n_733),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_918),
.B(n_703),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_895),
.B(n_742),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_898),
.B(n_707),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_884),
.B(n_750),
.Y(n_995)
);

NAND2xp33_ASAP7_75t_SL g996 ( 
.A(n_885),
.B(n_751),
.Y(n_996)
);

NAND2xp33_ASAP7_75t_SL g997 ( 
.A(n_923),
.B(n_759),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_925),
.B(n_760),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_928),
.B(n_763),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_932),
.B(n_767),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_935),
.B(n_775),
.Y(n_1001)
);

NAND2xp33_ASAP7_75t_SL g1002 ( 
.A(n_938),
.B(n_941),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_949),
.B(n_779),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_899),
.B(n_717),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_952),
.B(n_781),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_955),
.B(n_784),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_958),
.B(n_790),
.Y(n_1007)
);

NAND2xp33_ASAP7_75t_SL g1008 ( 
.A(n_961),
.B(n_773),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_967),
.B(n_789),
.Y(n_1009)
);

NAND2xp33_ASAP7_75t_SL g1010 ( 
.A(n_968),
.B(n_777),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_970),
.B(n_666),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_931),
.B(n_711),
.Y(n_1012)
);

NAND2xp33_ASAP7_75t_SL g1013 ( 
.A(n_904),
.B(n_754),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_922),
.B(n_756),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_940),
.B(n_716),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_947),
.B(n_951),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_962),
.B(n_716),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_926),
.B(n_728),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_893),
.B(n_890),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_929),
.B(n_728),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_942),
.B(n_562),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_962),
.B(n_1),
.Y(n_1022)
);

NAND2xp33_ASAP7_75t_SL g1023 ( 
.A(n_937),
.B(n_761),
.Y(n_1023)
);

NAND2xp33_ASAP7_75t_SL g1024 ( 
.A(n_939),
.B(n_563),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_943),
.B(n_915),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_933),
.B(n_571),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_897),
.B(n_1),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_972),
.B(n_572),
.Y(n_1028)
);

NAND2xp33_ASAP7_75t_SL g1029 ( 
.A(n_954),
.B(n_575),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_973),
.B(n_578),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_936),
.B(n_579),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_974),
.B(n_581),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_913),
.B(n_2),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_SL g1034 ( 
.A(n_894),
.B(n_749),
.Y(n_1034)
);

XNOR2x2_ASAP7_75t_L g1035 ( 
.A(n_901),
.B(n_725),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_948),
.B(n_753),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_950),
.B(n_762),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_953),
.B(n_772),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_902),
.B(n_586),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_900),
.B(n_589),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_908),
.B(n_592),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_946),
.B(n_726),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_924),
.B(n_593),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_959),
.B(n_965),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_945),
.B(n_595),
.Y(n_1045)
);

NAND2xp33_ASAP7_75t_SL g1046 ( 
.A(n_966),
.B(n_768),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_956),
.B(n_597),
.Y(n_1047)
);

NAND2xp33_ASAP7_75t_SL g1048 ( 
.A(n_919),
.B(n_598),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_905),
.B(n_729),
.Y(n_1049)
);

NAND2xp33_ASAP7_75t_SL g1050 ( 
.A(n_888),
.B(n_745),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_917),
.B(n_601),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_930),
.B(n_605),
.Y(n_1052)
);

NAND2xp33_ASAP7_75t_SL g1053 ( 
.A(n_971),
.B(n_607),
.Y(n_1053)
);

NAND2xp33_ASAP7_75t_SL g1054 ( 
.A(n_910),
.B(n_610),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_964),
.B(n_611),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_916),
.B(n_613),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_934),
.B(n_616),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_946),
.B(n_739),
.Y(n_1058)
);

NAND2xp33_ASAP7_75t_SL g1059 ( 
.A(n_927),
.B(n_766),
.Y(n_1059)
);

NAND2xp33_ASAP7_75t_SL g1060 ( 
.A(n_906),
.B(n_617),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_903),
.B(n_625),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_886),
.B(n_634),
.Y(n_1062)
);

NAND2xp33_ASAP7_75t_SL g1063 ( 
.A(n_907),
.B(n_738),
.Y(n_1063)
);

NAND2xp33_ASAP7_75t_SL g1064 ( 
.A(n_907),
.B(n_740),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_963),
.B(n_642),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_912),
.B(n_656),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_912),
.B(n_657),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_912),
.B(n_658),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_912),
.B(n_661),
.Y(n_1069)
);

NAND2xp33_ASAP7_75t_SL g1070 ( 
.A(n_907),
.B(n_765),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_912),
.B(n_662),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_912),
.B(n_665),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_912),
.B(n_676),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_912),
.B(n_677),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_912),
.B(n_678),
.Y(n_1075)
);

AND2x2_ASAP7_75t_SL g1076 ( 
.A(n_888),
.B(n_583),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_912),
.B(n_683),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_912),
.B(n_685),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_912),
.B(n_691),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_887),
.B(n_699),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_912),
.B(n_708),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_963),
.B(n_710),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_912),
.B(n_712),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_912),
.B(n_719),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_912),
.B(n_720),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_912),
.B(n_727),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_963),
.B(n_732),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_963),
.B(n_734),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_912),
.B(n_735),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_912),
.B(n_736),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_912),
.B(n_746),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_963),
.B(n_747),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_912),
.B(n_758),
.Y(n_1093)
);

NAND2xp33_ASAP7_75t_SL g1094 ( 
.A(n_907),
.B(n_771),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_912),
.B(n_641),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_940),
.B(n_2),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_912),
.B(n_652),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_912),
.B(n_674),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_963),
.B(n_3),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_912),
.B(n_689),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1044),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_984),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_984),
.B(n_769),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1019),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1002),
.A2(n_584),
.B(n_569),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1036),
.Y(n_1106)
);

AOI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1025),
.A2(n_686),
.B(n_603),
.Y(n_1107)
);

AND2x2_ASAP7_75t_SL g1108 ( 
.A(n_1076),
.B(n_568),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1037),
.A2(n_748),
.B(n_603),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1038),
.A2(n_748),
.B(n_603),
.Y(n_1110)
);

O2A1O1Ixp5_ASAP7_75t_SL g1111 ( 
.A1(n_1057),
.A2(n_603),
.B(n_748),
.C(n_568),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1099),
.A2(n_748),
.B(n_603),
.Y(n_1112)
);

OA22x2_ASAP7_75t_L g1113 ( 
.A1(n_1016),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_992),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_SL g1115 ( 
.A1(n_1065),
.A2(n_7),
.B(n_4),
.C(n_6),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_978),
.A2(n_9),
.B(n_7),
.C(n_8),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1009),
.A2(n_286),
.B(n_285),
.Y(n_1117)
);

BUFx12f_ASAP7_75t_L g1118 ( 
.A(n_1042),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_988),
.B(n_9),
.Y(n_1119)
);

INVxp67_ASAP7_75t_SL g1120 ( 
.A(n_994),
.Y(n_1120)
);

CKINVDCx11_ASAP7_75t_R g1121 ( 
.A(n_1042),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_1063),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_990),
.B(n_10),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1096),
.B(n_11),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1014),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1095),
.A2(n_288),
.B(n_287),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1082),
.A2(n_15),
.B(n_12),
.C(n_14),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1087),
.A2(n_12),
.B(n_14),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1088),
.B(n_1092),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_994),
.Y(n_1130)
);

AND2x2_ASAP7_75t_SL g1131 ( 
.A(n_1022),
.B(n_764),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1001),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1004),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1080),
.B(n_16),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1060),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1004),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1021),
.A2(n_290),
.B(n_289),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_989),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1097),
.A2(n_294),
.B(n_291),
.Y(n_1139)
);

INVx4_ASAP7_75t_L g1140 ( 
.A(n_1058),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_987),
.A2(n_296),
.B(n_295),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_980),
.B(n_21),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_975),
.B(n_22),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1098),
.A2(n_299),
.B(n_297),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1059),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_1027),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1100),
.A2(n_301),
.B(n_300),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_SL g1148 ( 
.A1(n_1018),
.A2(n_304),
.B(n_303),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1017),
.B(n_23),
.Y(n_1149)
);

AO31x2_ASAP7_75t_L g1150 ( 
.A1(n_1049),
.A2(n_306),
.A3(n_307),
.B(n_305),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_983),
.B(n_25),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1053),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_1152)
);

NAND2x1p5_ASAP7_75t_L g1153 ( 
.A(n_1056),
.B(n_308),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1033),
.Y(n_1154)
);

AO21x2_ASAP7_75t_L g1155 ( 
.A1(n_1020),
.A2(n_310),
.B(n_309),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_981),
.B(n_27),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1026),
.A2(n_313),
.B(n_311),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1035),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1012),
.B(n_28),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_1064),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_SL g1161 ( 
.A(n_1070),
.B(n_28),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_995),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_996),
.B(n_30),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1028),
.A2(n_316),
.B(n_314),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_997),
.B(n_30),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_1051),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_998),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_999),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1066),
.A2(n_31),
.B(n_32),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1067),
.B(n_32),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1068),
.B(n_33),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1030),
.A2(n_318),
.B(n_317),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1069),
.B(n_33),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1040),
.A2(n_322),
.B(n_321),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1000),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1071),
.A2(n_325),
.B(n_323),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1072),
.B(n_34),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1041),
.A2(n_327),
.B(n_326),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1073),
.A2(n_330),
.B(n_329),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1074),
.A2(n_332),
.B(n_331),
.Y(n_1180)
);

NOR4xp25_ASAP7_75t_L g1181 ( 
.A(n_1061),
.B(n_37),
.C(n_35),
.D(n_36),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1039),
.A2(n_336),
.B(n_334),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1052),
.A2(n_338),
.B(n_337),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1075),
.A2(n_341),
.B(n_340),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1077),
.B(n_37),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1078),
.A2(n_38),
.B(n_40),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1079),
.A2(n_41),
.B1(n_38),
.B2(n_40),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1055),
.A2(n_345),
.B(n_342),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1054),
.A2(n_349),
.A3(n_350),
.B(n_346),
.Y(n_1189)
);

NAND2xp33_ASAP7_75t_L g1190 ( 
.A(n_1008),
.B(n_42),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1081),
.A2(n_352),
.B(n_351),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1031),
.B(n_42),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1048),
.B(n_43),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1062),
.B(n_44),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1046),
.A2(n_356),
.A3(n_357),
.B(n_353),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1003),
.A2(n_359),
.B(n_358),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1083),
.B(n_44),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1084),
.A2(n_45),
.B(n_46),
.Y(n_1198)
);

NAND3xp33_ASAP7_75t_SL g1199 ( 
.A(n_1034),
.B(n_55),
.C(n_47),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1109),
.A2(n_1006),
.B(n_1005),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1102),
.B(n_986),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1131),
.A2(n_1094),
.B1(n_1010),
.B2(n_985),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1104),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1125),
.B(n_1047),
.Y(n_1204)
);

AO21x2_ASAP7_75t_L g1205 ( 
.A1(n_1112),
.A2(n_1086),
.B(n_1085),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1110),
.A2(n_1007),
.B(n_993),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_1114),
.Y(n_1207)
);

AND2x2_ASAP7_75t_SL g1208 ( 
.A(n_1108),
.B(n_1050),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1107),
.A2(n_1117),
.B(n_1126),
.Y(n_1209)
);

AO21x2_ASAP7_75t_L g1210 ( 
.A1(n_1129),
.A2(n_1090),
.B(n_1089),
.Y(n_1210)
);

OR2x6_ASAP7_75t_L g1211 ( 
.A(n_1118),
.B(n_1032),
.Y(n_1211)
);

INVx4_ASAP7_75t_L g1212 ( 
.A(n_1121),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1101),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1119),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_1130),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_SL g1216 ( 
.A1(n_1158),
.A2(n_1015),
.B1(n_1043),
.B2(n_1011),
.Y(n_1216)
);

NAND3xp33_ASAP7_75t_L g1217 ( 
.A(n_1190),
.B(n_1045),
.C(n_1091),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1133),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1139),
.A2(n_1093),
.B(n_977),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1144),
.A2(n_976),
.B(n_991),
.Y(n_1220)
);

AOI221xp5_ASAP7_75t_L g1221 ( 
.A1(n_1181),
.A2(n_982),
.B1(n_979),
.B2(n_1023),
.C(n_1013),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1134),
.A2(n_1029),
.B(n_1024),
.C(n_50),
.Y(n_1222)
);

OAI221xp5_ASAP7_75t_L g1223 ( 
.A1(n_1142),
.A2(n_51),
.B1(n_48),
.B2(n_49),
.C(n_52),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1166),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1147),
.A2(n_364),
.B(n_360),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1157),
.A2(n_367),
.B(n_366),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1123),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_1227)
);

AO21x2_ASAP7_75t_L g1228 ( 
.A1(n_1105),
.A2(n_369),
.B(n_368),
.Y(n_1228)
);

AO21x1_ASAP7_75t_L g1229 ( 
.A1(n_1128),
.A2(n_54),
.B(n_55),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1106),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1164),
.A2(n_371),
.B(n_370),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1172),
.A2(n_373),
.B(n_372),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1124),
.A2(n_376),
.B(n_375),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1176),
.A2(n_378),
.B(n_377),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1111),
.A2(n_380),
.B(n_379),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_SL g1236 ( 
.A1(n_1149),
.A2(n_57),
.B1(n_54),
.B2(n_56),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1143),
.A2(n_1156),
.B(n_1151),
.C(n_1138),
.Y(n_1237)
);

AOI211xp5_ASAP7_75t_SL g1238 ( 
.A1(n_1115),
.A2(n_59),
.B(n_60),
.C(n_58),
.Y(n_1238)
);

NAND2x1p5_ASAP7_75t_L g1239 ( 
.A(n_1160),
.B(n_382),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1167),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1175),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1136),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1196),
.A2(n_385),
.B(n_384),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1174),
.A2(n_388),
.B(n_386),
.Y(n_1244)
);

OAI211xp5_ASAP7_75t_L g1245 ( 
.A1(n_1135),
.A2(n_1152),
.B(n_1159),
.C(n_1186),
.Y(n_1245)
);

NOR2x1_ASAP7_75t_SL g1246 ( 
.A(n_1155),
.B(n_59),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1162),
.Y(n_1247)
);

NOR2xp67_ASAP7_75t_L g1248 ( 
.A(n_1122),
.B(n_390),
.Y(n_1248)
);

OAI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1161),
.A2(n_69),
.B1(n_77),
.B2(n_61),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1166),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1146),
.B(n_61),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1178),
.A2(n_392),
.B(n_391),
.Y(n_1252)
);

AO21x2_ASAP7_75t_L g1253 ( 
.A1(n_1179),
.A2(n_394),
.B(n_393),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1169),
.A2(n_62),
.B(n_63),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1154),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1168),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1182),
.A2(n_398),
.B(n_397),
.Y(n_1257)
);

OA21x2_ASAP7_75t_L g1258 ( 
.A1(n_1183),
.A2(n_402),
.B(n_400),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1192),
.B(n_63),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1188),
.A2(n_404),
.B(n_403),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1120),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1137),
.A2(n_406),
.B(n_405),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_SL g1263 ( 
.A1(n_1198),
.A2(n_66),
.B(n_65),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1103),
.Y(n_1264)
);

AO21x2_ASAP7_75t_L g1265 ( 
.A1(n_1180),
.A2(n_408),
.B(n_407),
.Y(n_1265)
);

OA21x2_ASAP7_75t_L g1266 ( 
.A1(n_1141),
.A2(n_411),
.B(n_410),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1150),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1113),
.A2(n_68),
.B1(n_64),
.B2(n_67),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1194),
.B(n_67),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1184),
.A2(n_416),
.B(n_412),
.Y(n_1270)
);

AOI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1191),
.A2(n_419),
.B(n_417),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1199),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1272)
);

AO21x2_ASAP7_75t_L g1273 ( 
.A1(n_1170),
.A2(n_421),
.B(n_420),
.Y(n_1273)
);

NOR2x1p5_ASAP7_75t_L g1274 ( 
.A(n_1171),
.B(n_71),
.Y(n_1274)
);

BUFx12f_ASAP7_75t_L g1275 ( 
.A(n_1153),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1148),
.A2(n_423),
.B(n_422),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1127),
.A2(n_1116),
.B(n_1173),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1177),
.A2(n_425),
.B(n_424),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1185),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1145),
.A2(n_427),
.B(n_426),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_SL g1281 ( 
.A(n_1187),
.B(n_428),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1197),
.A2(n_430),
.B(n_429),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1163),
.A2(n_432),
.B(n_431),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1132),
.A2(n_72),
.B(n_73),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1193),
.Y(n_1285)
);

AO21x1_ASAP7_75t_L g1286 ( 
.A1(n_1165),
.A2(n_73),
.B(n_74),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1150),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1195),
.A2(n_434),
.B(n_433),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1195),
.A2(n_436),
.B(n_435),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_1189),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1104),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1125),
.B(n_74),
.Y(n_1292)
);

NOR2xp67_ASAP7_75t_L g1293 ( 
.A(n_1140),
.B(n_437),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1109),
.A2(n_440),
.B(n_439),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1121),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1102),
.B(n_75),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1109),
.A2(n_442),
.B(n_441),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1125),
.B(n_75),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1129),
.A2(n_78),
.B(n_79),
.C(n_77),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1104),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1129),
.A2(n_444),
.B(n_443),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1104),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1104),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1125),
.B(n_76),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1125),
.B(n_76),
.Y(n_1305)
);

OA21x2_ASAP7_75t_L g1306 ( 
.A1(n_1112),
.A2(n_446),
.B(n_445),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1118),
.Y(n_1307)
);

INVx2_ASAP7_75t_SL g1308 ( 
.A(n_1224),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1207),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1213),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1203),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1242),
.B(n_79),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1208),
.A2(n_83),
.B1(n_80),
.B2(n_81),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1251),
.B(n_1296),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1215),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1209),
.A2(n_449),
.B(n_447),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1291),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1300),
.Y(n_1318)
);

INVxp67_ASAP7_75t_SL g1319 ( 
.A(n_1218),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1302),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1250),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1303),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1269),
.B(n_85),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1230),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1255),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1264),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1307),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1201),
.B(n_86),
.Y(n_1328)
);

AOI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1287),
.A2(n_452),
.B(n_451),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1274),
.B(n_87),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1275),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1256),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1240),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1241),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1247),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1237),
.B(n_88),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1239),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1214),
.Y(n_1338)
);

INVx4_ASAP7_75t_L g1339 ( 
.A(n_1295),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1211),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1285),
.Y(n_1341)
);

CKINVDCx11_ASAP7_75t_R g1342 ( 
.A(n_1295),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1279),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_1212),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1292),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1298),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1285),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1304),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1204),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1305),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1293),
.B(n_89),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1210),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1277),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1236),
.B(n_1259),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1229),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1220),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1273),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1202),
.B(n_90),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1286),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1254),
.A2(n_90),
.B(n_91),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1200),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1283),
.Y(n_1362)
);

BUFx12f_ASAP7_75t_L g1363 ( 
.A(n_1290),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1206),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_SL g1365 ( 
.A1(n_1246),
.A2(n_92),
.B(n_93),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1263),
.Y(n_1366)
);

NAND2x1_ASAP7_75t_L g1367 ( 
.A(n_1280),
.B(n_1266),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1219),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1227),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1278),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1205),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1284),
.B(n_92),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_R g1373 ( 
.A(n_1342),
.B(n_1281),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1332),
.Y(n_1374)
);

INVxp67_ASAP7_75t_L g1375 ( 
.A(n_1309),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_R g1376 ( 
.A(n_1344),
.B(n_1268),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1319),
.B(n_1249),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1325),
.B(n_1248),
.Y(n_1378)
);

INVxp67_ASAP7_75t_L g1379 ( 
.A(n_1314),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1326),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1341),
.B(n_1217),
.Y(n_1381)
);

CKINVDCx11_ASAP7_75t_R g1382 ( 
.A(n_1339),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1308),
.B(n_1222),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1335),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_1339),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1310),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_R g1387 ( 
.A(n_1331),
.B(n_1337),
.Y(n_1387)
);

XNOR2xp5_ASAP7_75t_L g1388 ( 
.A(n_1340),
.B(n_1216),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_R g1389 ( 
.A(n_1337),
.B(n_1321),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_R g1390 ( 
.A(n_1347),
.B(n_1271),
.Y(n_1390)
);

XNOR2xp5_ASAP7_75t_L g1391 ( 
.A(n_1328),
.B(n_1261),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1323),
.B(n_1238),
.Y(n_1392)
);

XNOR2xp5_ASAP7_75t_L g1393 ( 
.A(n_1327),
.B(n_1330),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1315),
.B(n_1349),
.Y(n_1394)
);

NAND2xp33_ASAP7_75t_R g1395 ( 
.A(n_1312),
.B(n_1306),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_1363),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1343),
.B(n_1299),
.Y(n_1397)
);

NAND2xp33_ASAP7_75t_R g1398 ( 
.A(n_1347),
.B(n_1266),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1348),
.B(n_1245),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_R g1400 ( 
.A(n_1345),
.B(n_1272),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1358),
.B(n_93),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1346),
.B(n_1223),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1350),
.B(n_95),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_R g1404 ( 
.A(n_1354),
.B(n_96),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1338),
.B(n_1267),
.Y(n_1405)
);

AND2x2_ASAP7_75t_SL g1406 ( 
.A(n_1372),
.B(n_1221),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1324),
.B(n_1282),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1333),
.Y(n_1408)
);

OR2x6_ASAP7_75t_L g1409 ( 
.A(n_1351),
.B(n_1233),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1336),
.B(n_97),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1317),
.B(n_98),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1394),
.B(n_1353),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1375),
.B(n_1352),
.Y(n_1413)
);

NOR2x1p5_ASAP7_75t_L g1414 ( 
.A(n_1380),
.B(n_1369),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1406),
.A2(n_1313),
.B1(n_1360),
.B2(n_1351),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1374),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1373),
.B(n_1359),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1399),
.B(n_1386),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_SL g1419 ( 
.A(n_1387),
.B(n_1355),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1379),
.B(n_1318),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1384),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1377),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1405),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1407),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1408),
.Y(n_1425)
);

NOR2x1p5_ASAP7_75t_L g1426 ( 
.A(n_1402),
.B(n_1366),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1404),
.A2(n_1334),
.B1(n_1320),
.B2(n_1322),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1385),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1392),
.B(n_1371),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1397),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1381),
.B(n_1371),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1403),
.B(n_1361),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1395),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1382),
.Y(n_1434)
);

OAI221xp5_ASAP7_75t_L g1435 ( 
.A1(n_1401),
.A2(n_1367),
.B1(n_1301),
.B2(n_1370),
.C(n_1234),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1393),
.B(n_1356),
.Y(n_1436)
);

INVxp67_ASAP7_75t_SL g1437 ( 
.A(n_1398),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1411),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1383),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1410),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1409),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1389),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1378),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1409),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1400),
.B(n_1311),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1391),
.A2(n_1367),
.B1(n_1362),
.B2(n_1356),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1396),
.B(n_1364),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1388),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1390),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1376),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1428),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1416),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1430),
.B(n_1368),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1436),
.B(n_1362),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1422),
.B(n_1357),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1449),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1413),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1429),
.B(n_1316),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1413),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1412),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1418),
.B(n_1288),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1432),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1447),
.B(n_1253),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1444),
.B(n_1329),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1420),
.B(n_1289),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1441),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1423),
.Y(n_1467)
);

AND2x2_ASAP7_75t_SL g1468 ( 
.A(n_1442),
.B(n_1258),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1421),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1434),
.Y(n_1470)
);

OR2x6_ASAP7_75t_L g1471 ( 
.A(n_1414),
.B(n_1365),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1426),
.B(n_1438),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1425),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1439),
.B(n_99),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_SL g1475 ( 
.A(n_1450),
.B(n_1276),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1443),
.B(n_1265),
.Y(n_1476)
);

AND4x1_ASAP7_75t_L g1477 ( 
.A(n_1415),
.B(n_101),
.C(n_99),
.D(n_100),
.Y(n_1477)
);

INVx1_ASAP7_75t_SL g1478 ( 
.A(n_1443),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1440),
.B(n_1258),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1431),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1431),
.B(n_1228),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1437),
.A2(n_1262),
.B(n_1270),
.Y(n_1482)
);

OAI222xp33_ASAP7_75t_L g1483 ( 
.A1(n_1427),
.A2(n_1243),
.B1(n_104),
.B2(n_106),
.C1(n_102),
.C2(n_103),
.Y(n_1483)
);

NOR2x1p5_ASAP7_75t_L g1484 ( 
.A(n_1445),
.B(n_103),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1424),
.B(n_1243),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1446),
.B(n_104),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1448),
.A2(n_1226),
.B1(n_1232),
.B2(n_1231),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1417),
.B(n_105),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1435),
.B(n_1257),
.Y(n_1489)
);

NOR2x1_ASAP7_75t_L g1490 ( 
.A(n_1414),
.B(n_105),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1415),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1433),
.A2(n_1244),
.B1(n_1252),
.B2(n_1260),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1413),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1414),
.Y(n_1494)
);

AO21x2_ASAP7_75t_L g1495 ( 
.A1(n_1437),
.A2(n_1297),
.B(n_1294),
.Y(n_1495)
);

AND2x2_ASAP7_75t_SL g1496 ( 
.A(n_1442),
.B(n_109),
.Y(n_1496)
);

NAND4xp75_ASAP7_75t_L g1497 ( 
.A(n_1419),
.B(n_111),
.C(n_109),
.D(n_110),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1416),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1413),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1416),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1416),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1442),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1442),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1456),
.B(n_1225),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1498),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1500),
.B(n_112),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1501),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1462),
.B(n_113),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1460),
.B(n_114),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1452),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1503),
.B(n_1494),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1467),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1473),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1466),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1478),
.B(n_1454),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1480),
.B(n_1472),
.Y(n_1516)
);

NOR2x1_ASAP7_75t_R g1517 ( 
.A(n_1451),
.B(n_116),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1455),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1469),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_SL g1520 ( 
.A(n_1502),
.B(n_1235),
.Y(n_1520)
);

AND2x2_ASAP7_75t_SL g1521 ( 
.A(n_1496),
.B(n_117),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1457),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1476),
.B(n_1471),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1459),
.Y(n_1524)
);

NOR2xp67_ASAP7_75t_L g1525 ( 
.A(n_1486),
.B(n_120),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1463),
.B(n_120),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1493),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1499),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1458),
.B(n_121),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1465),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1479),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1461),
.B(n_1468),
.Y(n_1532)
);

CKINVDCx16_ASAP7_75t_R g1533 ( 
.A(n_1490),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1488),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1471),
.B(n_123),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1489),
.B(n_123),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1474),
.B(n_124),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1484),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1485),
.B(n_129),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1464),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1464),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1481),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1475),
.B(n_1482),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1495),
.B(n_130),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1477),
.B(n_130),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1497),
.B(n_1483),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1492),
.B(n_1487),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1498),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1453),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1503),
.B(n_131),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1491),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1453),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1498),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1498),
.B(n_132),
.Y(n_1554)
);

AND2x4_ASAP7_75t_SL g1555 ( 
.A(n_1470),
.B(n_133),
.Y(n_1555)
);

INVx3_ASAP7_75t_L g1556 ( 
.A(n_1470),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1498),
.Y(n_1557)
);

AND2x4_ASAP7_75t_SL g1558 ( 
.A(n_1470),
.B(n_134),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1462),
.B(n_134),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1498),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1502),
.B(n_135),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1460),
.B(n_137),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1557),
.B(n_138),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1505),
.B(n_139),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1507),
.B(n_1548),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1518),
.Y(n_1566)
);

AO221x2_ASAP7_75t_L g1567 ( 
.A1(n_1554),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.C(n_143),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1546),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1510),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1553),
.B(n_147),
.Y(n_1570)
);

NOR2xp67_ASAP7_75t_L g1571 ( 
.A(n_1541),
.B(n_148),
.Y(n_1571)
);

OAI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1543),
.A2(n_150),
.B1(n_151),
.B2(n_149),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1540),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1515),
.B(n_152),
.Y(n_1574)
);

CKINVDCx20_ASAP7_75t_R g1575 ( 
.A(n_1555),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1556),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1523),
.B(n_153),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1558),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1523),
.B(n_156),
.Y(n_1579)
);

OAI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1536),
.A2(n_159),
.B1(n_160),
.B2(n_158),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1560),
.B(n_157),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1544),
.B(n_162),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1512),
.Y(n_1583)
);

OR2x6_ASAP7_75t_L g1584 ( 
.A(n_1550),
.B(n_163),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1530),
.B(n_163),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1526),
.B(n_164),
.Y(n_1586)
);

NAND2xp33_ASAP7_75t_R g1587 ( 
.A(n_1535),
.B(n_165),
.Y(n_1587)
);

AO221x1_ASAP7_75t_L g1588 ( 
.A1(n_1542),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.C(n_169),
.Y(n_1588)
);

INVxp67_ASAP7_75t_SL g1589 ( 
.A(n_1525),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1547),
.B(n_170),
.Y(n_1590)
);

AO221x2_ASAP7_75t_L g1591 ( 
.A1(n_1517),
.A2(n_1514),
.B1(n_1521),
.B2(n_1539),
.C(n_1549),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1516),
.Y(n_1592)
);

NOR2x1_ASAP7_75t_L g1593 ( 
.A(n_1508),
.B(n_171),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1538),
.B(n_172),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1529),
.B(n_173),
.Y(n_1595)
);

AO221x2_ASAP7_75t_L g1596 ( 
.A1(n_1552),
.A2(n_177),
.B1(n_174),
.B2(n_176),
.C(n_178),
.Y(n_1596)
);

OAI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1534),
.A2(n_180),
.B1(n_177),
.B2(n_179),
.Y(n_1597)
);

NOR2x1_ASAP7_75t_L g1598 ( 
.A(n_1559),
.B(n_181),
.Y(n_1598)
);

INVxp33_ASAP7_75t_SL g1599 ( 
.A(n_1561),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1562),
.B(n_182),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1513),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1531),
.B(n_183),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1545),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1504),
.B(n_189),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1537),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1519),
.B(n_1522),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1524),
.B(n_191),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1527),
.B(n_192),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_SL g1609 ( 
.A1(n_1551),
.A2(n_1528),
.B1(n_1520),
.B2(n_194),
.Y(n_1609)
);

AO221x2_ASAP7_75t_L g1610 ( 
.A1(n_1506),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.C(n_196),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1557),
.B(n_193),
.Y(n_1611)
);

CKINVDCx20_ASAP7_75t_R g1612 ( 
.A(n_1533),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_1511),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1557),
.B(n_198),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1557),
.B(n_199),
.Y(n_1615)
);

NAND2xp33_ASAP7_75t_SL g1616 ( 
.A(n_1509),
.B(n_199),
.Y(n_1616)
);

NOR2x1_ASAP7_75t_L g1617 ( 
.A(n_1556),
.B(n_200),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_R g1618 ( 
.A(n_1535),
.B(n_201),
.Y(n_1618)
);

NOR2xp67_ASAP7_75t_L g1619 ( 
.A(n_1532),
.B(n_202),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1557),
.B(n_203),
.Y(n_1620)
);

INVx6_ASAP7_75t_L g1621 ( 
.A(n_1584),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1583),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1575),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1566),
.B(n_204),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1587),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1569),
.Y(n_1626)
);

CKINVDCx16_ASAP7_75t_R g1627 ( 
.A(n_1618),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1590),
.B(n_205),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1592),
.B(n_205),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1565),
.B(n_206),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1601),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1604),
.B(n_206),
.Y(n_1632)
);

NOR3xp33_ASAP7_75t_SL g1633 ( 
.A(n_1609),
.B(n_1576),
.C(n_1572),
.Y(n_1633)
);

CKINVDCx16_ASAP7_75t_R g1634 ( 
.A(n_1578),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1599),
.B(n_207),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1584),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1606),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1574),
.B(n_208),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1589),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1585),
.B(n_209),
.Y(n_1640)
);

NAND2x1p5_ASAP7_75t_L g1641 ( 
.A(n_1617),
.B(n_210),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1563),
.B(n_210),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1607),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1577),
.B(n_211),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1602),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1611),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1605),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1614),
.Y(n_1648)
);

OAI31xp33_ASAP7_75t_SL g1649 ( 
.A1(n_1593),
.A2(n_214),
.A3(n_212),
.B(n_213),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1615),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1564),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1608),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1620),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1570),
.B(n_215),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1598),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1581),
.B(n_216),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1582),
.B(n_1595),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1579),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1596),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1600),
.B(n_217),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1571),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1596),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1586),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1619),
.B(n_1603),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1594),
.B(n_219),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1616),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1610),
.B(n_220),
.Y(n_1667)
);

OAI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1568),
.A2(n_225),
.B1(n_222),
.B2(n_224),
.C(n_226),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1597),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1567),
.B(n_226),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1580),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1588),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1583),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1583),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1587),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1613),
.B(n_228),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1573),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1566),
.B(n_229),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1599),
.B(n_232),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1573),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1583),
.Y(n_1681)
);

NOR2x1_ASAP7_75t_L g1682 ( 
.A(n_1612),
.B(n_233),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1591),
.A2(n_234),
.B(n_235),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1565),
.B(n_235),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1583),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1583),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1583),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1583),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1583),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1573),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1583),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1583),
.Y(n_1692)
);

INVx1_ASAP7_75t_SL g1693 ( 
.A(n_1612),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1583),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1583),
.Y(n_1695)
);

NOR2x1_ASAP7_75t_L g1696 ( 
.A(n_1612),
.B(n_236),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1583),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1566),
.B(n_237),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1591),
.A2(n_241),
.B1(n_238),
.B2(n_240),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1583),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1566),
.B(n_241),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1573),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1612),
.Y(n_1703)
);

INVx2_ASAP7_75t_SL g1704 ( 
.A(n_1612),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1599),
.B(n_243),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1566),
.B(n_243),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1683),
.A2(n_244),
.B(n_245),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1621),
.Y(n_1708)
);

OAI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1699),
.A2(n_247),
.B1(n_245),
.B2(n_246),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1651),
.B(n_246),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1674),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1634),
.B(n_247),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1633),
.A2(n_248),
.B(n_249),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1692),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1622),
.Y(n_1715)
);

INVxp67_ASAP7_75t_L g1716 ( 
.A(n_1704),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1639),
.Y(n_1717)
);

OR4x1_ASAP7_75t_L g1718 ( 
.A(n_1672),
.B(n_252),
.C(n_250),
.D(n_251),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1626),
.Y(n_1719)
);

OR2x6_ASAP7_75t_L g1720 ( 
.A(n_1636),
.B(n_252),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1659),
.B(n_253),
.Y(n_1721)
);

AOI21xp33_ASAP7_75t_SL g1722 ( 
.A1(n_1627),
.A2(n_254),
.B(n_256),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1673),
.Y(n_1723)
);

XOR2x2_ASAP7_75t_L g1724 ( 
.A(n_1682),
.B(n_256),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1681),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1693),
.B(n_259),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1662),
.B(n_262),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1646),
.B(n_262),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1685),
.Y(n_1729)
);

INVx2_ASAP7_75t_SL g1730 ( 
.A(n_1623),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1686),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1663),
.B(n_1643),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1687),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1688),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1637),
.B(n_264),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1689),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1691),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1676),
.B(n_1703),
.Y(n_1738)
);

NOR2xp67_ASAP7_75t_L g1739 ( 
.A(n_1666),
.B(n_266),
.Y(n_1739)
);

NOR2x1_ASAP7_75t_L g1740 ( 
.A(n_1696),
.B(n_267),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_L g1741 ( 
.A(n_1649),
.B(n_268),
.C(n_269),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1694),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1664),
.A2(n_273),
.B1(n_271),
.B2(n_272),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1695),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1697),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1664),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_1746)
);

NOR2x1p5_ASAP7_75t_SL g1747 ( 
.A(n_1631),
.B(n_276),
.Y(n_1747)
);

INVxp67_ASAP7_75t_L g1748 ( 
.A(n_1657),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1648),
.B(n_1650),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1700),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1653),
.B(n_277),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1625),
.A2(n_278),
.B(n_279),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1675),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1647),
.Y(n_1754)
);

AND2x2_ASAP7_75t_SL g1755 ( 
.A(n_1667),
.B(n_283),
.Y(n_1755)
);

INVxp67_ASAP7_75t_SL g1756 ( 
.A(n_1655),
.Y(n_1756)
);

AOI222xp33_ASAP7_75t_L g1757 ( 
.A1(n_1670),
.A2(n_456),
.B1(n_459),
.B2(n_454),
.C1(n_455),
.C2(n_457),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1645),
.B(n_460),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1624),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1678),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1698),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1701),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1661),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1671),
.Y(n_1764)
);

INVxp67_ASAP7_75t_SL g1765 ( 
.A(n_1641),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1706),
.Y(n_1766)
);

AOI21xp33_ASAP7_75t_L g1767 ( 
.A1(n_1668),
.A2(n_1669),
.B(n_1684),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1652),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1658),
.B(n_475),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1730),
.B(n_1754),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1748),
.B(n_1629),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1732),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1738),
.B(n_1705),
.Y(n_1773)
);

INVxp67_ASAP7_75t_SL g1774 ( 
.A(n_1739),
.Y(n_1774)
);

CKINVDCx20_ASAP7_75t_R g1775 ( 
.A(n_1724),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1716),
.B(n_1635),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1749),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1764),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1710),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1717),
.Y(n_1780)
);

NAND2x1_ASAP7_75t_SL g1781 ( 
.A(n_1740),
.B(n_1638),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1759),
.B(n_1630),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1712),
.B(n_1665),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1760),
.B(n_1642),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1728),
.B(n_1751),
.Y(n_1785)
);

NOR2x1_ASAP7_75t_L g1786 ( 
.A(n_1713),
.B(n_1679),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1715),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1765),
.B(n_1644),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1741),
.A2(n_1628),
.B1(n_1660),
.B2(n_1654),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1719),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1761),
.B(n_1632),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1762),
.B(n_1766),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1747),
.B(n_1656),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1735),
.B(n_1640),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1723),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1768),
.B(n_1677),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1755),
.B(n_1680),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1763),
.B(n_1690),
.Y(n_1798)
);

NAND2xp33_ASAP7_75t_SL g1799 ( 
.A(n_1711),
.B(n_1702),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1720),
.B(n_479),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1714),
.B(n_1756),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1725),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1729),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1731),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1733),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1734),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1780),
.Y(n_1807)
);

BUFx4f_ASAP7_75t_SL g1808 ( 
.A(n_1788),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1792),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1778),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1770),
.B(n_1722),
.Y(n_1811)
);

CKINVDCx20_ASAP7_75t_R g1812 ( 
.A(n_1775),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1784),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1781),
.Y(n_1814)
);

INVxp33_ASAP7_75t_SL g1815 ( 
.A(n_1776),
.Y(n_1815)
);

INVxp33_ASAP7_75t_SL g1816 ( 
.A(n_1773),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1787),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1783),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1790),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1795),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1802),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1803),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1799),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1804),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1785),
.B(n_1708),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1805),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1806),
.Y(n_1827)
);

OAI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1812),
.A2(n_1786),
.B(n_1707),
.Y(n_1828)
);

NAND2xp33_ASAP7_75t_L g1829 ( 
.A(n_1814),
.B(n_1771),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_SL g1830 ( 
.A(n_1816),
.B(n_1774),
.Y(n_1830)
);

OAI211xp5_ASAP7_75t_L g1831 ( 
.A1(n_1823),
.A2(n_1801),
.B(n_1772),
.C(n_1777),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1815),
.B(n_1789),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1808),
.B(n_1811),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1825),
.A2(n_1793),
.B(n_1752),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1818),
.B(n_1794),
.Y(n_1835)
);

NOR4xp25_ASAP7_75t_L g1836 ( 
.A(n_1807),
.B(n_1779),
.C(n_1721),
.D(n_1727),
.Y(n_1836)
);

AOI221xp5_ASAP7_75t_L g1837 ( 
.A1(n_1813),
.A2(n_1718),
.B1(n_1767),
.B2(n_1709),
.C(n_1797),
.Y(n_1837)
);

NOR3x1_ASAP7_75t_L g1838 ( 
.A(n_1810),
.B(n_1791),
.C(n_1782),
.Y(n_1838)
);

NAND4xp25_ASAP7_75t_L g1839 ( 
.A(n_1830),
.B(n_1809),
.C(n_1819),
.D(n_1817),
.Y(n_1839)
);

NAND3xp33_ASAP7_75t_SL g1840 ( 
.A(n_1828),
.B(n_1743),
.C(n_1757),
.Y(n_1840)
);

AOI221xp5_ASAP7_75t_L g1841 ( 
.A1(n_1836),
.A2(n_1821),
.B1(n_1824),
.B2(n_1822),
.C(n_1820),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1835),
.Y(n_1842)
);

O2A1O1Ixp33_ASAP7_75t_L g1843 ( 
.A1(n_1829),
.A2(n_1827),
.B(n_1826),
.C(n_1726),
.Y(n_1843)
);

BUFx6f_ASAP7_75t_L g1844 ( 
.A(n_1842),
.Y(n_1844)
);

XNOR2x1_ASAP7_75t_L g1845 ( 
.A(n_1840),
.B(n_1832),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1839),
.Y(n_1846)
);

HB1xp67_ASAP7_75t_L g1847 ( 
.A(n_1841),
.Y(n_1847)
);

NAND3xp33_ASAP7_75t_L g1848 ( 
.A(n_1847),
.B(n_1845),
.C(n_1844),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_R g1849 ( 
.A(n_1846),
.B(n_1833),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1848),
.Y(n_1850)
);

INVx3_ASAP7_75t_L g1851 ( 
.A(n_1850),
.Y(n_1851)
);

A2O1A1Ixp33_ASAP7_75t_L g1852 ( 
.A1(n_1851),
.A2(n_1843),
.B(n_1834),
.C(n_1837),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1852),
.A2(n_1798),
.B1(n_1849),
.B2(n_1796),
.Y(n_1853)
);

XNOR2xp5_ASAP7_75t_L g1854 ( 
.A(n_1853),
.B(n_1831),
.Y(n_1854)
);

AOI222xp33_ASAP7_75t_SL g1855 ( 
.A1(n_1854),
.A2(n_1838),
.B1(n_1737),
.B2(n_1742),
.C1(n_1745),
.C2(n_1744),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1855),
.Y(n_1856)
);

OAI221xp5_ASAP7_75t_R g1857 ( 
.A1(n_1856),
.A2(n_1753),
.B1(n_1746),
.B2(n_1736),
.C(n_1750),
.Y(n_1857)
);

AOI211xp5_ASAP7_75t_L g1858 ( 
.A1(n_1857),
.A2(n_1800),
.B(n_1758),
.C(n_1769),
.Y(n_1858)
);


endmodule