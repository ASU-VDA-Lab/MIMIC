module fake_jpeg_5369_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_4),
.B(n_3),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_8),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

AOI21xp33_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_0),
.B(n_1),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_23),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_2),
.B(n_3),
.C(n_5),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_2),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_27),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_27),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_29),
.B(n_31),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_34),
.A2(n_23),
.B1(n_26),
.B2(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_40),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_16),
.B1(n_14),
.B2(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_12),
.B(n_25),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_11),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_13),
.B1(n_11),
.B2(n_3),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_11),
.B1(n_13),
.B2(n_5),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_11),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_53),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_47),
.C(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_56),
.B(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_62),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_43),
.C(n_41),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_61),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_54),
.B1(n_47),
.B2(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_49),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_49),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_47),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_70),
.C(n_69),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_66),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_72),
.C(n_73),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_64),
.B(n_51),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_75),
.A2(n_74),
.B1(n_45),
.B2(n_7),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_40),
.Y(n_77)
);


endmodule