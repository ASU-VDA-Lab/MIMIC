module fake_jpeg_4210_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_12),
.B(n_10),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_SL g25 ( 
.A(n_14),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_6),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_43),
.B(n_19),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_26),
.Y(n_44)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_50),
.Y(n_93)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_65),
.Y(n_96)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_21),
.B(n_6),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_24),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVxp67_ASAP7_75t_SL g56 ( 
.A(n_25),
.Y(n_56)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_66),
.Y(n_72)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_63),
.A2(n_64),
.B1(n_68),
.B2(n_35),
.Y(n_83)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_29),
.Y(n_99)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_69),
.B(n_75),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_39),
.B1(n_42),
.B2(n_41),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_70),
.A2(n_74),
.B1(n_30),
.B2(n_28),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_39),
.B1(n_22),
.B2(n_41),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_73),
.A2(n_95),
.B1(n_97),
.B2(n_102),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_41),
.B1(n_22),
.B2(n_24),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_44),
.B(n_38),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_94),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_22),
.B(n_35),
.C(n_29),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_18),
.B1(n_31),
.B2(n_27),
.Y(n_121)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_84),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_82),
.B(n_110),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_36),
.B(n_34),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_85),
.A2(n_106),
.B(n_4),
.C(n_11),
.Y(n_145)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_89),
.Y(n_133)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_20),
.B1(n_19),
.B2(n_27),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_59),
.A2(n_35),
.B1(n_36),
.B2(n_28),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_38),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_103),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_99),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_60),
.A2(n_35),
.B1(n_36),
.B2(n_34),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_67),
.A2(n_34),
.B1(n_30),
.B2(n_28),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_4),
.B1(n_11),
.B2(n_9),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_45),
.B(n_18),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_43),
.B(n_32),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_115),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_101),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_116),
.Y(n_180)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_124),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_121),
.A2(n_77),
.B1(n_78),
.B2(n_84),
.Y(n_164)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_128),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_32),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_130),
.Y(n_155)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_72),
.B(n_30),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_75),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_88),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_82),
.A2(n_31),
.B1(n_20),
.B2(n_33),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_88),
.A2(n_33),
.B1(n_29),
.B2(n_8),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_140),
.Y(n_170)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_141),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_76),
.B(n_4),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_142),
.B(n_77),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_15),
.B(n_1),
.C(n_3),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_105),
.B1(n_91),
.B2(n_100),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_113),
.A2(n_8),
.B1(n_11),
.B2(n_9),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_91),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_96),
.B(n_8),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_147),
.B(n_15),
.Y(n_161)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_83),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_149),
.A2(n_151),
.B1(n_102),
.B2(n_97),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_104),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_151)
);

NAND2xp33_ASAP7_75t_SL g207 ( 
.A(n_153),
.B(n_185),
.Y(n_207)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_154),
.B(n_161),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_93),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_159),
.C(n_146),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_80),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_158),
.B(n_163),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_113),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_162),
.A2(n_165),
.B1(n_149),
.B2(n_150),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_78),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_L g218 ( 
.A(n_164),
.B(n_172),
.C(n_184),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_92),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_168),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_0),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_0),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_175),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_123),
.A2(n_15),
.B(n_3),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_186),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_3),
.Y(n_175)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_89),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_107),
.Y(n_181)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_122),
.B(n_107),
.Y(n_182)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_129),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_136),
.B(n_105),
.Y(n_187)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_149),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_185),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_189),
.B(n_195),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_187),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_197),
.B(n_206),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_219),
.B1(n_169),
.B2(n_157),
.Y(n_222)
);

XOR2x2_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_150),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_202),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_179),
.A2(n_118),
.B(n_133),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_216),
.B(n_171),
.Y(n_229)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_205),
.Y(n_237)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_209),
.B(n_211),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_214),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_152),
.A2(n_114),
.B1(n_128),
.B2(n_141),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_115),
.B1(n_163),
.B2(n_177),
.Y(n_234)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_155),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_217),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_155),
.A2(n_131),
.B(n_125),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_162),
.A2(n_158),
.B(n_157),
.C(n_163),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_158),
.A2(n_115),
.B1(n_140),
.B2(n_138),
.Y(n_219)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_180),
.Y(n_244)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_226),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_196),
.Y(n_224)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_200),
.A2(n_159),
.B1(n_169),
.B2(n_154),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_227),
.A2(n_241),
.B1(n_191),
.B2(n_196),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_208),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_233),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_236),
.B(n_193),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_180),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_232),
.B(n_205),
.Y(n_258)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_201),
.Y(n_235)
);

INVx13_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

AO22x1_ASAP7_75t_L g236 ( 
.A1(n_188),
.A2(n_165),
.B1(n_125),
.B2(n_168),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_246),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_186),
.C(n_175),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_202),
.C(n_216),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_217),
.A2(n_173),
.B1(n_177),
.B2(n_124),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_244),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_206),
.A2(n_194),
.B1(n_214),
.B2(n_212),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_245),
.A2(n_199),
.B1(n_190),
.B2(n_204),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_211),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_198),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_225),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_250),
.A2(n_251),
.B(n_260),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_194),
.B(n_203),
.Y(n_251)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_222),
.B1(n_232),
.B2(n_223),
.Y(n_273)
);

AOI21xp33_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_207),
.B(n_210),
.Y(n_255)
);

AOI321xp33_ASAP7_75t_L g284 ( 
.A1(n_255),
.A2(n_258),
.A3(n_259),
.B1(n_238),
.B2(n_246),
.C(n_170),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_268),
.C(n_241),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_230),
.A2(n_199),
.B(n_210),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_237),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_226),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_233),
.A2(n_195),
.B(n_189),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_234),
.B1(n_236),
.B2(n_221),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_239),
.B(n_218),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_232),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_235),
.B(n_148),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_278),
.C(n_281),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_284),
.B(n_252),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_227),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_277),
.C(n_285),
.Y(n_296)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_262),
.B(n_228),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_274),
.B(n_252),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_261),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_276),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_224),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_229),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_268),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_248),
.A2(n_236),
.B1(n_240),
.B2(n_245),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_SL g291 ( 
.A1(n_280),
.A2(n_254),
.B(n_257),
.C(n_248),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_266),
.B1(n_257),
.B2(n_285),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_183),
.C(n_231),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_286),
.A2(n_291),
.B(n_294),
.Y(n_306)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_288),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_247),
.Y(n_304)
);

BUFx12f_ASAP7_75t_SL g294 ( 
.A(n_278),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_282),
.B1(n_273),
.B2(n_280),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_263),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_297),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_270),
.B(n_264),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_299),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_250),
.C(n_267),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_271),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_309),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_282),
.B(n_266),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_265),
.B(n_251),
.Y(n_317)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_304),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_247),
.Y(n_305)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_305),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_308),
.A2(n_292),
.B1(n_298),
.B2(n_291),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_277),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_281),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_289),
.C(n_299),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_301),
.B(n_260),
.Y(n_311)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_311),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_314),
.B(n_318),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_291),
.B1(n_302),
.B2(n_303),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_317),
.A2(n_306),
.B(n_264),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_261),
.C(n_291),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_324),
.B(n_316),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_323),
.C(n_318),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_315),
.A2(n_306),
.B1(n_307),
.B2(n_284),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_312),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_312),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_327),
.B(n_328),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_324),
.A2(n_314),
.B(n_307),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_300),
.C(n_320),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_329),
.C(n_309),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_117),
.Y(n_333)
);


endmodule