module fake_jpeg_10755_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_3),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx8_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx4_ASAP7_75t_SL g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_10),
.B(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_16),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_0),
.Y(n_17)
);

FAx1_ASAP7_75t_SL g25 ( 
.A(n_17),
.B(n_13),
.CI(n_12),
.CON(n_25),
.SN(n_25)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_19),
.Y(n_24)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_7),
.B(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_27),
.B(n_26),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_29),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_34),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_32),
.B(n_25),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_16),
.C(n_17),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_24),
.C(n_23),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_26),
.A2(n_20),
.B1(n_14),
.B2(n_19),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_33),
.A2(n_29),
.B1(n_11),
.B2(n_25),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_11),
.B(n_21),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_12),
.B1(n_1),
.B2(n_6),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_43),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_5),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_5),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_48),
.B1(n_45),
.B2(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_42),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_12),
.Y(n_50)
);


endmodule