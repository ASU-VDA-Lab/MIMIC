module fake_jpeg_29760_n_45 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_45);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_45;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_23),
.B1(n_19),
.B2(n_2),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_23)
);

AOI222xp33_ASAP7_75t_L g24 ( 
.A1(n_17),
.A2(n_21),
.B1(n_20),
.B2(n_19),
.C1(n_3),
.C2(n_4),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_25),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_29),
.B1(n_32),
.B2(n_6),
.Y(n_37)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_1),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_8),
.C(n_2),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_27),
.C(n_5),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_37),
.Y(n_40)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_33),
.B1(n_36),
.B2(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_40),
.Y(n_43)
);

NOR3xp33_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_41),
.C(n_7),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_4),
.Y(n_45)
);


endmodule