module fake_jpeg_2712_n_563 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_563);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_563;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_54),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_55),
.B(n_57),
.Y(n_121)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_56),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_20),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_58),
.B(n_62),
.Y(n_128)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_59),
.Y(n_165)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_0),
.Y(n_61)
);

NAND2x1p5_ASAP7_75t_L g132 ( 
.A(n_61),
.B(n_37),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_26),
.B(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_9),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_63),
.B(n_64),
.Y(n_155)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

OR2x2_ASAP7_75t_SL g66 ( 
.A(n_23),
.B(n_10),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_66),
.B(n_102),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_68),
.Y(n_159)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_69),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_72),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_22),
.B(n_52),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_73),
.B(n_74),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_19),
.B(n_10),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_20),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_76),
.B(n_85),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_34),
.Y(n_77)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_27),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_86),
.B(n_87),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_10),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g134 ( 
.A(n_95),
.B(n_97),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_101),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_31),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_33),
.B(n_0),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_33),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_104),
.Y(n_116)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_25),
.B1(n_51),
.B2(n_49),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_119),
.A2(n_130),
.B1(n_135),
.B2(n_137),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_47),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_28),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_61),
.A2(n_40),
.B1(n_48),
.B2(n_45),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_123),
.B(n_142),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_41),
.B1(n_33),
.B2(n_48),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_143),
.B1(n_144),
.B2(n_146),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_77),
.A2(n_94),
.B1(n_99),
.B2(n_95),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_132),
.B(n_81),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_75),
.A2(n_25),
.B1(n_51),
.B2(n_52),
.Y(n_135)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_80),
.A2(n_25),
.B1(n_105),
.B2(n_97),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_61),
.A2(n_41),
.B1(n_48),
.B2(n_45),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_79),
.A2(n_45),
.B1(n_40),
.B2(n_48),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_90),
.A2(n_52),
.B1(n_51),
.B2(n_47),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_106),
.A2(n_21),
.B1(n_42),
.B2(n_32),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_73),
.A2(n_45),
.B1(n_44),
.B2(n_36),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_152),
.A2(n_158),
.B1(n_162),
.B2(n_40),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_82),
.A2(n_44),
.B1(n_36),
.B2(n_41),
.Y(n_153)
);

AO22x1_ASAP7_75t_L g177 ( 
.A1(n_153),
.A2(n_37),
.B1(n_84),
.B2(n_44),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_66),
.A2(n_34),
.B(n_37),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_154),
.Y(n_176)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_83),
.A2(n_29),
.B1(n_42),
.B2(n_32),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_104),
.A2(n_29),
.B1(n_28),
.B2(n_98),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_167),
.B(n_180),
.Y(n_234)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx3_ASAP7_75t_SL g241 ( 
.A(n_169),
.Y(n_241)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

INVx3_ASAP7_75t_SL g257 ( 
.A(n_171),
.Y(n_257)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_172),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_112),
.B(n_122),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_173),
.B(n_178),
.Y(n_275)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_174),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_175),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_177),
.A2(n_125),
.B1(n_153),
.B2(n_143),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_65),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_181),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_59),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_182),
.B(n_186),
.Y(n_239)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_183),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_114),
.B(n_56),
.C(n_71),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_132),
.C(n_151),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_128),
.B(n_78),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_121),
.B(n_68),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_187),
.B(n_191),
.Y(n_267)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_188),
.Y(n_253)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_189),
.Y(n_264)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_190),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_120),
.B(n_91),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_192),
.B(n_210),
.Y(n_246)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_193),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_117),
.B(n_60),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_199),
.Y(n_235)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_196),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_197),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_120),
.B(n_67),
.Y(n_199)
);

INVx4_ASAP7_75t_SL g200 ( 
.A(n_160),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_200),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_111),
.B(n_67),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_201),
.Y(n_249)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_111),
.Y(n_202)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_202),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_114),
.B(n_88),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_203),
.B(n_208),
.Y(n_260)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_133),
.Y(n_204)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_204),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_139),
.B(n_89),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_205),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_147),
.Y(n_206)
);

NAND2xp33_ASAP7_75t_SL g229 ( 
.A(n_206),
.B(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_116),
.B(n_89),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_139),
.B(n_72),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_209),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_118),
.Y(n_210)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_110),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_211),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_150),
.Y(n_212)
);

NAND2xp33_ASAP7_75t_SL g231 ( 
.A(n_212),
.B(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_150),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_145),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_214),
.B(n_215),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_124),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_259)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_138),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_140),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_126),
.B(n_72),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_220),
.B(n_223),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_221),
.A2(n_148),
.B1(n_34),
.B2(n_113),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_116),
.A2(n_40),
.B1(n_44),
.B2(n_41),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_123),
.B1(n_142),
.B2(n_156),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_132),
.B(n_36),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_126),
.B(n_36),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_224),
.B(n_213),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_225),
.A2(n_232),
.B1(n_243),
.B2(n_252),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_168),
.A2(n_147),
.B1(n_154),
.B2(n_141),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_227),
.A2(n_244),
.B1(n_251),
.B2(n_254),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_228),
.B(n_247),
.C(n_250),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_176),
.A2(n_134),
.B(n_149),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_233),
.A2(n_4),
.B(n_5),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_L g243 ( 
.A1(n_176),
.A2(n_140),
.B1(n_107),
.B2(n_115),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_170),
.A2(n_203),
.B1(n_223),
.B2(n_177),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_184),
.B(n_127),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_208),
.B(n_127),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_170),
.A2(n_141),
.B1(n_129),
.B2(n_165),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_192),
.A2(n_129),
.B1(n_138),
.B2(n_107),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_198),
.A2(n_115),
.B1(n_136),
.B2(n_166),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_192),
.B(n_165),
.C(n_166),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_256),
.B(n_265),
.C(n_24),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_262),
.A2(n_24),
.B1(n_35),
.B2(n_175),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_172),
.B(n_159),
.C(n_124),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_177),
.A2(n_134),
.B1(n_148),
.B2(n_159),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_271),
.A2(n_273),
.B1(n_189),
.B2(n_163),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_167),
.A2(n_163),
.B1(n_92),
.B2(n_54),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_274),
.B(n_200),
.Y(n_292)
);

OA22x2_ASAP7_75t_L g276 ( 
.A1(n_181),
.A2(n_69),
.B1(n_24),
.B2(n_113),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_212),
.Y(n_278)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_226),
.Y(n_277)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_277),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_278),
.B(n_282),
.Y(n_366)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_226),
.Y(n_279)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_190),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_280),
.B(n_296),
.Y(n_350)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_281),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_246),
.A2(n_188),
.B1(n_202),
.B2(n_215),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_244),
.A2(n_207),
.B1(n_211),
.B2(n_174),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_283),
.A2(n_284),
.B1(n_288),
.B2(n_307),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_227),
.A2(n_185),
.B1(n_179),
.B2(n_219),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_239),
.B(n_195),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_286),
.B(n_291),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_260),
.A2(n_179),
.B1(n_185),
.B2(n_219),
.Y(n_288)
);

OR2x6_ASAP7_75t_SL g289 ( 
.A(n_233),
.B(n_69),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_289),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_230),
.B(n_193),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g343 ( 
.A(n_290),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_230),
.B(n_218),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_292),
.B(n_297),
.Y(n_334)
);

A2O1A1O1Ixp25_ASAP7_75t_L g293 ( 
.A1(n_266),
.A2(n_169),
.B(n_171),
.C(n_204),
.D(n_196),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_293),
.A2(n_295),
.B(n_310),
.Y(n_328)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_242),
.Y(n_294)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_294),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_229),
.A2(n_217),
.B(n_216),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_247),
.B(n_183),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_263),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_298),
.B(n_276),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_210),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_300),
.B(n_308),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_238),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_301),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_SL g357 ( 
.A(n_302),
.B(n_306),
.Y(n_357)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_253),
.Y(n_303)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_303),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_248),
.B(n_210),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_304),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_248),
.B(n_235),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_305),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_275),
.B(n_234),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_275),
.B(n_175),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_249),
.B(n_267),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_309),
.B(n_314),
.Y(n_352)
);

OAI21xp33_ASAP7_75t_L g310 ( 
.A1(n_246),
.A2(n_2),
.B(n_4),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_253),
.Y(n_311)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_311),
.Y(n_363)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_258),
.Y(n_312)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_312),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_228),
.B(n_17),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_323),
.C(n_237),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_250),
.B(n_2),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_258),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_315),
.B(n_316),
.Y(n_362)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_241),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_225),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_232),
.B1(n_252),
.B2(n_257),
.Y(n_335)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_268),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_318),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_319),
.A2(n_263),
.B(n_265),
.Y(n_336)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_268),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_320),
.Y(n_338)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_241),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_321),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_246),
.A2(n_274),
.B(n_231),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_322),
.A2(n_324),
.B(n_231),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_256),
.B(n_4),
.Y(n_323)
);

NOR2x1_ASAP7_75t_L g324 ( 
.A(n_271),
.B(n_273),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_287),
.B(n_251),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_325),
.B(n_346),
.C(n_347),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_332),
.A2(n_339),
.B(n_353),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_333),
.B(n_298),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_335),
.B(n_283),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_336),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_285),
.A2(n_254),
.B1(n_269),
.B2(n_238),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_337),
.A2(n_345),
.B1(n_349),
.B2(n_356),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_322),
.A2(n_259),
.B(n_245),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_285),
.A2(n_269),
.B1(n_276),
.B2(n_261),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_287),
.B(n_270),
.C(n_272),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_297),
.A2(n_272),
.B1(n_261),
.B2(n_276),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_348),
.A2(n_360),
.B1(n_361),
.B2(n_321),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_280),
.A2(n_257),
.B1(n_241),
.B2(n_245),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_289),
.A2(n_264),
.B(n_255),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_313),
.B(n_264),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_355),
.B(n_365),
.C(n_295),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_299),
.A2(n_257),
.B1(n_236),
.B2(n_255),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_299),
.A2(n_236),
.B1(n_240),
.B2(n_7),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_286),
.A2(n_240),
.B1(n_6),
.B2(n_7),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_296),
.B(n_5),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_300),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_370),
.B(n_372),
.Y(n_414)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_340),
.Y(n_371)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_371),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_358),
.B(n_279),
.Y(n_372)
);

AOI22x1_ASAP7_75t_L g373 ( 
.A1(n_366),
.A2(n_278),
.B1(n_289),
.B2(n_284),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_373),
.A2(n_376),
.B1(n_403),
.B2(n_405),
.Y(n_411)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_340),
.Y(n_377)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_377),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_378),
.B(n_384),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_282),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_379),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_325),
.B(n_323),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_380),
.B(n_387),
.C(n_398),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_334),
.B(n_314),
.Y(n_381)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_381),
.Y(n_413)
);

AO22x1_ASAP7_75t_L g382 ( 
.A1(n_341),
.A2(n_302),
.B1(n_317),
.B2(n_288),
.Y(n_382)
);

OA21x2_ASAP7_75t_L g428 ( 
.A1(n_382),
.A2(n_349),
.B(n_363),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_362),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_383),
.B(n_385),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_362),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_351),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_386),
.B(n_388),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_312),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_358),
.B(n_281),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_315),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_397),
.Y(n_407)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_326),
.Y(n_390)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_390),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_329),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_391),
.B(n_402),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_343),
.B(n_277),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_392),
.B(n_395),
.Y(n_430)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_326),
.Y(n_393)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_393),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_332),
.A2(n_319),
.B(n_324),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_394),
.A2(n_399),
.B(n_404),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_351),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_331),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_396),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_350),
.B(n_311),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_355),
.B(n_294),
.C(n_320),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_341),
.A2(n_324),
.B(n_293),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_367),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_400),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_318),
.Y(n_401)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_401),
.Y(n_434)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_327),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_366),
.A2(n_303),
.B(n_316),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_331),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_374),
.A2(n_345),
.B1(n_366),
.B2(n_337),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_408),
.A2(n_382),
.B1(n_369),
.B2(n_373),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_380),
.B(n_346),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_412),
.B(n_423),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_374),
.A2(n_335),
.B1(n_330),
.B2(n_356),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_415),
.A2(n_425),
.B1(n_431),
.B2(n_432),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_368),
.B(n_333),
.C(n_365),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_422),
.B(n_384),
.C(n_398),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_368),
.B(n_336),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_387),
.B(n_352),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_424),
.B(n_429),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_376),
.A2(n_330),
.B1(n_328),
.B2(n_339),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_401),
.A2(n_329),
.B1(n_338),
.B2(n_328),
.Y(n_426)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_426),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_375),
.A2(n_338),
.B(n_363),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_427),
.A2(n_436),
.B(n_404),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_428),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_378),
.B(n_352),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_394),
.A2(n_359),
.B1(n_354),
.B2(n_344),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_379),
.A2(n_359),
.B1(n_354),
.B2(n_344),
.Y(n_432)
);

OAI32xp33_ASAP7_75t_L g435 ( 
.A1(n_379),
.A2(n_327),
.A3(n_342),
.B1(n_301),
.B2(n_367),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_435),
.B(n_391),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_375),
.A2(n_342),
.B(n_301),
.Y(n_436)
);

BUFx24_ASAP7_75t_SL g440 ( 
.A(n_414),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_440),
.B(n_466),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_413),
.B(n_381),
.Y(n_441)
);

NAND3xp33_ASAP7_75t_L g480 ( 
.A(n_441),
.B(n_463),
.C(n_464),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_443),
.A2(n_421),
.B(n_436),
.Y(n_476)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_420),
.Y(n_444)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_444),
.Y(n_477)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_438),
.Y(n_445)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_445),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_446),
.B(n_422),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_447),
.A2(n_458),
.B1(n_428),
.B2(n_434),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_448),
.A2(n_459),
.B1(n_428),
.B2(n_431),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_420),
.B(n_389),
.Y(n_449)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_449),
.Y(n_486)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_419),
.Y(n_450)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_450),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_423),
.B(n_409),
.C(n_418),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_451),
.B(n_454),
.C(n_468),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_417),
.B(n_397),
.Y(n_452)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_452),
.Y(n_491)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_438),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_453),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_409),
.B(n_373),
.C(n_369),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_411),
.A2(n_382),
.B1(n_390),
.B2(n_402),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_408),
.A2(n_399),
.B1(n_393),
.B2(n_377),
.Y(n_459)
);

FAx1_ASAP7_75t_SL g460 ( 
.A(n_427),
.B(n_371),
.CI(n_400),
.CON(n_460),
.SN(n_460)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_460),
.B(n_465),
.Y(n_469)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_430),
.Y(n_462)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_462),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_413),
.B(n_5),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_429),
.B(n_6),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_406),
.B(n_6),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_437),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_412),
.B(n_6),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_467),
.B(n_407),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_418),
.B(n_7),
.C(n_8),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_433),
.Y(n_471)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_471),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_473),
.B(n_478),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_424),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_479),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_476),
.A2(n_483),
.B(n_443),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_451),
.B(n_407),
.C(n_439),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_461),
.B(n_439),
.Y(n_479)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_481),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_447),
.A2(n_434),
.B(n_425),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_484),
.B(n_455),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_485),
.A2(n_488),
.B1(n_460),
.B2(n_459),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_456),
.A2(n_458),
.B1(n_442),
.B2(n_457),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_454),
.B(n_432),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_467),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_455),
.B(n_433),
.C(n_415),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_490),
.B(n_446),
.C(n_468),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_493),
.B(n_498),
.Y(n_520)
);

OAI221xp5_ASAP7_75t_L g495 ( 
.A1(n_486),
.A2(n_444),
.B1(n_456),
.B2(n_452),
.C(n_448),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_495),
.Y(n_511)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_496),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_483),
.A2(n_435),
.B(n_460),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_499),
.B(n_504),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_500),
.B(n_482),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_471),
.Y(n_501)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_501),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_491),
.B(n_465),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g524 ( 
.A(n_502),
.B(n_505),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_453),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_473),
.B(n_416),
.C(n_410),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_508),
.C(n_475),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_475),
.B(n_445),
.C(n_10),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_469),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_510),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_470),
.B(n_480),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_512),
.B(n_518),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_503),
.A2(n_485),
.B1(n_477),
.B2(n_469),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_513),
.A2(n_495),
.B1(n_494),
.B2(n_501),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_493),
.A2(n_476),
.B(n_489),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_514),
.A2(n_522),
.B(n_494),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_503),
.A2(n_479),
.B1(n_490),
.B2(n_472),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_517),
.B(n_523),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_499),
.B(n_478),
.C(n_474),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_484),
.C(n_472),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_519),
.B(n_525),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_498),
.A2(n_487),
.B(n_482),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_506),
.B(n_7),
.C(n_11),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_497),
.B(n_11),
.C(n_12),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_527),
.B(n_11),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_521),
.B(n_508),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_532),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_530),
.B(n_535),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_511),
.A2(n_502),
.B1(n_497),
.B2(n_500),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_533),
.B(n_536),
.Y(n_548)
);

BUFx24_ASAP7_75t_SL g534 ( 
.A(n_515),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_534),
.B(n_526),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_520),
.A2(n_11),
.B(n_12),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_520),
.A2(n_13),
.B(n_14),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_537),
.B(n_538),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_522),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_512),
.B(n_13),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_540),
.B(n_541),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_518),
.B(n_13),
.C(n_16),
.Y(n_541)
);

O2A1O1Ixp33_ASAP7_75t_SL g542 ( 
.A1(n_538),
.A2(n_524),
.B(n_516),
.C(n_513),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_542),
.A2(n_546),
.B(n_539),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_544),
.B(n_545),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_528),
.B(n_531),
.Y(n_545)
);

O2A1O1Ixp33_ASAP7_75t_SL g546 ( 
.A1(n_539),
.A2(n_514),
.B(n_517),
.C(n_523),
.Y(n_546)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_547),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_551),
.B(n_554),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_543),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_552),
.A2(n_553),
.B(n_541),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_548),
.B(n_540),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_555),
.A2(n_519),
.B(n_547),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_556),
.A2(n_557),
.B(n_558),
.Y(n_559)
);

NOR3xp33_ASAP7_75t_SL g560 ( 
.A(n_557),
.B(n_549),
.C(n_550),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_560),
.B(n_559),
.C(n_527),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_561),
.B(n_525),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_562),
.A2(n_13),
.B(n_16),
.Y(n_563)
);


endmodule