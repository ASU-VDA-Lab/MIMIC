module fake_aes_7865_n_1521 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1521);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1521;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1477;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_641;
wire n_379;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1520;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_799;
wire n_342;
wire n_423;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_606;
wire n_332;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_1455;
wire n_659;
wire n_432;
wire n_386;
wire n_1329;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1518;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1491;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1439;
wire n_374;
wire n_718;
wire n_1484;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g330 ( .A(n_77), .Y(n_330) );
INVxp67_ASAP7_75t_L g331 ( .A(n_221), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_289), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_260), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_44), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_70), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_101), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_182), .Y(n_338) );
CKINVDCx16_ASAP7_75t_R g339 ( .A(n_232), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_65), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_240), .Y(n_341) );
INVxp33_ASAP7_75t_SL g342 ( .A(n_208), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_130), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_193), .Y(n_344) );
CKINVDCx16_ASAP7_75t_R g345 ( .A(n_157), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_298), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_135), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_310), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_263), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_133), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_58), .Y(n_351) );
INVxp33_ASAP7_75t_L g352 ( .A(n_238), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_142), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_236), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_105), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_114), .Y(n_356) );
INVxp67_ASAP7_75t_SL g357 ( .A(n_301), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_108), .Y(n_358) );
INVxp33_ASAP7_75t_L g359 ( .A(n_162), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_322), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_73), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_83), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_152), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_87), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_103), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_227), .Y(n_366) );
CKINVDCx16_ASAP7_75t_R g367 ( .A(n_155), .Y(n_367) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_0), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_147), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_98), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_237), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_244), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_144), .Y(n_373) );
INVxp33_ASAP7_75t_L g374 ( .A(n_54), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_234), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_11), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_73), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_302), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_26), .Y(n_379) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_68), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_156), .Y(n_381) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_317), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_283), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_220), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_292), .Y(n_385) );
INVxp67_ASAP7_75t_SL g386 ( .A(n_318), .Y(n_386) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_204), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_49), .Y(n_388) );
INVxp67_ASAP7_75t_SL g389 ( .A(n_170), .Y(n_389) );
BUFx2_ASAP7_75t_L g390 ( .A(n_269), .Y(n_390) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_117), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_197), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_323), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_249), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_116), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_46), .Y(n_396) );
BUFx2_ASAP7_75t_SL g397 ( .A(n_107), .Y(n_397) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_18), .Y(n_398) );
INVxp67_ASAP7_75t_SL g399 ( .A(n_284), .Y(n_399) );
CKINVDCx16_ASAP7_75t_R g400 ( .A(n_153), .Y(n_400) );
INVxp33_ASAP7_75t_SL g401 ( .A(n_8), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_113), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_6), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_8), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_65), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_68), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_256), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_217), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_313), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_105), .Y(n_410) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_272), .Y(n_411) );
INVxp33_ASAP7_75t_SL g412 ( .A(n_12), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_20), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_69), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_48), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_21), .Y(n_416) );
INVxp33_ASAP7_75t_SL g417 ( .A(n_47), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_45), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_222), .Y(n_419) );
INVxp67_ASAP7_75t_SL g420 ( .A(n_101), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_55), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_51), .Y(n_422) );
INVxp67_ASAP7_75t_L g423 ( .A(n_115), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_178), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_37), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_184), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_306), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_31), .Y(n_428) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_209), .Y(n_429) );
INVxp33_ASAP7_75t_L g430 ( .A(n_5), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_81), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_30), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_199), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_327), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_44), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_18), .Y(n_436) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_201), .Y(n_437) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_250), .Y(n_438) );
INVxp33_ASAP7_75t_L g439 ( .A(n_61), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_90), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_20), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_171), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_320), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_216), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_134), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_11), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_59), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_235), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_48), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_195), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_281), .Y(n_451) );
INVxp33_ASAP7_75t_SL g452 ( .A(n_239), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_102), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_88), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_213), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_258), .Y(n_456) );
INVxp67_ASAP7_75t_SL g457 ( .A(n_56), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_24), .Y(n_458) );
INVxp33_ASAP7_75t_SL g459 ( .A(n_4), .Y(n_459) );
CKINVDCx16_ASAP7_75t_R g460 ( .A(n_128), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_96), .Y(n_461) );
INVxp33_ASAP7_75t_SL g462 ( .A(n_226), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_294), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_38), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_119), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_165), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_84), .Y(n_467) );
BUFx3_ASAP7_75t_L g468 ( .A(n_275), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_1), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_91), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_106), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_50), .Y(n_472) );
CKINVDCx14_ASAP7_75t_R g473 ( .A(n_168), .Y(n_473) );
INVxp67_ASAP7_75t_L g474 ( .A(n_180), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g475 ( .A(n_55), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_111), .Y(n_476) );
INVxp67_ASAP7_75t_SL g477 ( .A(n_129), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_84), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_188), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_169), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_15), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_104), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_161), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_196), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_316), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_47), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_145), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_123), .Y(n_488) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_19), .Y(n_489) );
INVxp33_ASAP7_75t_SL g490 ( .A(n_85), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_69), .Y(n_491) );
NOR2xp67_ASAP7_75t_L g492 ( .A(n_25), .B(n_54), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_360), .Y(n_493) );
INVx3_ASAP7_75t_L g494 ( .A(n_346), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_381), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_390), .B(n_0), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_360), .Y(n_497) );
INVx2_ASAP7_75t_SL g498 ( .A(n_390), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_391), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_363), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_362), .B(n_1), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_363), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_374), .B(n_2), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_366), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_366), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_372), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_346), .Y(n_507) );
BUFx8_ASAP7_75t_L g508 ( .A(n_391), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_372), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_373), .Y(n_510) );
INVx5_ASAP7_75t_L g511 ( .A(n_391), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_373), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_375), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_375), .Y(n_514) );
INVx3_ASAP7_75t_L g515 ( .A(n_347), .Y(n_515) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_391), .Y(n_516) );
OAI21x1_ASAP7_75t_L g517 ( .A1(n_347), .A2(n_110), .B(n_109), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_362), .B(n_2), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_391), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_378), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_378), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_438), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_430), .B(n_3), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_439), .B(n_3), .Y(n_524) );
XNOR2xp5_ASAP7_75t_L g525 ( .A(n_398), .B(n_4), .Y(n_525) );
NOR2x1_ASAP7_75t_L g526 ( .A(n_332), .B(n_5), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_438), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_371), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_438), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_480), .Y(n_530) );
BUFx3_ASAP7_75t_L g531 ( .A(n_508), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_493), .B(n_371), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_494), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_493), .B(n_393), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_511), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_511), .Y(n_536) );
NOR2xp33_ASAP7_75t_SL g537 ( .A(n_493), .B(n_339), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_495), .Y(n_538) );
BUFx4f_ASAP7_75t_L g539 ( .A(n_496), .Y(n_539) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_516), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_498), .B(n_475), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_496), .B(n_351), .Y(n_542) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_517), .A2(n_480), .B(n_338), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_503), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_498), .B(n_345), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_496), .B(n_351), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_494), .Y(n_547) );
BUFx2_ASAP7_75t_L g548 ( .A(n_496), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_496), .A2(n_412), .B1(n_417), .B2(n_401), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_497), .B(n_502), .Y(n_550) );
OAI22xp33_ASAP7_75t_L g551 ( .A1(n_498), .A2(n_489), .B1(n_425), .B2(n_403), .Y(n_551) );
INVx6_ASAP7_75t_L g552 ( .A(n_508), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_511), .Y(n_553) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_516), .Y(n_554) );
OR2x2_ASAP7_75t_SL g555 ( .A(n_525), .B(n_432), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_511), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_496), .A2(n_370), .B1(n_376), .B2(n_365), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_497), .B(n_388), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_503), .B(n_367), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_494), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_503), .B(n_400), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_511), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_497), .B(n_388), .Y(n_563) );
BUFx2_ASAP7_75t_L g564 ( .A(n_524), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_511), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_502), .B(n_431), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_511), .Y(n_567) );
AND2x6_ASAP7_75t_L g568 ( .A(n_526), .B(n_392), .Y(n_568) );
AND2x6_ASAP7_75t_L g569 ( .A(n_526), .B(n_392), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_494), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_511), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_524), .B(n_460), .Y(n_572) );
INVx4_ASAP7_75t_L g573 ( .A(n_511), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_502), .B(n_431), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_504), .B(n_446), .Y(n_575) );
INVx4_ASAP7_75t_L g576 ( .A(n_494), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_504), .B(n_446), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_550), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_576), .Y(n_579) );
INVx3_ASAP7_75t_L g580 ( .A(n_576), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_550), .Y(n_581) );
INVx4_ASAP7_75t_L g582 ( .A(n_552), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_576), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_576), .Y(n_584) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_531), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_544), .B(n_524), .Y(n_586) );
AOI22xp5_ASAP7_75t_SL g587 ( .A1(n_538), .A2(n_525), .B1(n_491), .B2(n_412), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_544), .Y(n_588) );
INVx5_ASAP7_75t_L g589 ( .A(n_552), .Y(n_589) );
BUFx12f_ASAP7_75t_L g590 ( .A(n_541), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_533), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_558), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_558), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_564), .B(n_523), .Y(n_594) );
AND2x4_ASAP7_75t_L g595 ( .A(n_548), .B(n_501), .Y(n_595) );
NAND2x1p5_ASAP7_75t_L g596 ( .A(n_539), .B(n_517), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_558), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_564), .B(n_500), .Y(n_598) );
INVx5_ASAP7_75t_L g599 ( .A(n_552), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_533), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_559), .B(n_523), .Y(n_601) );
INVx5_ASAP7_75t_L g602 ( .A(n_552), .Y(n_602) );
NOR2x1_ASAP7_75t_L g603 ( .A(n_541), .B(n_424), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_548), .B(n_500), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_542), .B(n_501), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_547), .Y(n_606) );
AND2x6_ASAP7_75t_SL g607 ( .A(n_559), .B(n_525), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g608 ( .A1(n_537), .A2(n_518), .B(n_520), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_547), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_560), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_559), .B(n_520), .Y(n_611) );
INVx2_ASAP7_75t_SL g612 ( .A(n_539), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_560), .Y(n_613) );
A2O1A1Ixp33_ASAP7_75t_L g614 ( .A1(n_539), .A2(n_504), .B(n_506), .C(n_505), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_570), .Y(n_615) );
AO21x2_ASAP7_75t_L g616 ( .A1(n_543), .A2(n_517), .B(n_506), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_539), .A2(n_506), .B1(n_509), .B2(n_505), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_558), .Y(n_618) );
INVx2_ASAP7_75t_SL g619 ( .A(n_552), .Y(n_619) );
CKINVDCx5p33_ASAP7_75t_R g620 ( .A(n_561), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_561), .A2(n_417), .B1(n_459), .B2(n_401), .Y(n_621) );
AND2x4_ASAP7_75t_L g622 ( .A(n_542), .B(n_518), .Y(n_622) );
INVx3_ASAP7_75t_L g623 ( .A(n_558), .Y(n_623) );
INVx3_ASAP7_75t_L g624 ( .A(n_563), .Y(n_624) );
INVx6_ASAP7_75t_L g625 ( .A(n_563), .Y(n_625) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_561), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_570), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_543), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_563), .Y(n_629) );
BUFx2_ASAP7_75t_L g630 ( .A(n_572), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_572), .B(n_521), .Y(n_631) );
INVxp67_ASAP7_75t_L g632 ( .A(n_537), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_572), .A2(n_490), .B1(n_459), .B2(n_334), .Y(n_633) );
BUFx2_ASAP7_75t_L g634 ( .A(n_531), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_563), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_563), .Y(n_636) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_531), .Y(n_637) );
NOR2x1p5_ASAP7_75t_SL g638 ( .A(n_535), .B(n_505), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_542), .B(n_521), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_542), .B(n_509), .Y(n_640) );
AND3x1_ASAP7_75t_SL g641 ( .A(n_555), .B(n_336), .C(n_330), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_549), .A2(n_490), .B1(n_355), .B2(n_361), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_566), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_557), .B(n_509), .Y(n_644) );
BUFx3_ASAP7_75t_L g645 ( .A(n_542), .Y(n_645) );
INVx2_ASAP7_75t_SL g646 ( .A(n_546), .Y(n_646) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_551), .Y(n_647) );
INVx1_ASAP7_75t_SL g648 ( .A(n_532), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_545), .B(n_352), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_543), .Y(n_650) );
CKINVDCx6p67_ASAP7_75t_R g651 ( .A(n_568), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_543), .Y(n_652) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_566), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_535), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_566), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_546), .B(n_510), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_546), .A2(n_512), .B1(n_513), .B2(n_510), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_546), .B(n_510), .Y(n_658) );
AND2x6_ASAP7_75t_SL g659 ( .A(n_555), .B(n_365), .Y(n_659) );
NOR2xp67_ASAP7_75t_L g660 ( .A(n_549), .B(n_512), .Y(n_660) );
BUFx2_ASAP7_75t_L g661 ( .A(n_568), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_566), .Y(n_662) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_566), .Y(n_663) );
INVx2_ASAP7_75t_SL g664 ( .A(n_546), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_532), .A2(n_456), .B1(n_479), .B2(n_451), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_574), .B(n_530), .Y(n_666) );
OR2x4_ASAP7_75t_L g667 ( .A(n_534), .B(n_512), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_574), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_574), .Y(n_669) );
INVxp67_ASAP7_75t_SL g670 ( .A(n_578), .Y(n_670) );
INVx2_ASAP7_75t_SL g671 ( .A(n_667), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_578), .Y(n_672) );
NAND2x1p5_ASAP7_75t_L g673 ( .A(n_648), .B(n_574), .Y(n_673) );
BUFx12f_ASAP7_75t_L g674 ( .A(n_607), .Y(n_674) );
INVx1_ASAP7_75t_SL g675 ( .A(n_634), .Y(n_675) );
NOR2xp67_ASAP7_75t_L g676 ( .A(n_642), .B(n_574), .Y(n_676) );
AOI21x1_ASAP7_75t_L g677 ( .A1(n_628), .A2(n_534), .B(n_517), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_646), .Y(n_678) );
OR2x6_ASAP7_75t_L g679 ( .A(n_665), .B(n_575), .Y(n_679) );
A2O1A1Ixp33_ASAP7_75t_L g680 ( .A1(n_581), .A2(n_577), .B(n_575), .C(n_514), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_605), .B(n_575), .Y(n_681) );
BUFx4f_ASAP7_75t_SL g682 ( .A(n_590), .Y(n_682) );
BUFx2_ASAP7_75t_L g683 ( .A(n_590), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_645), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_645), .Y(n_685) );
NAND2x1p5_ASAP7_75t_L g686 ( .A(n_623), .B(n_575), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_605), .B(n_575), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_626), .B(n_551), .Y(n_688) );
AOI222xp33_ASAP7_75t_L g689 ( .A1(n_630), .A2(n_464), .B1(n_461), .B2(n_457), .C1(n_380), .C2(n_420), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_601), .A2(n_569), .B1(n_568), .B2(n_577), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_646), .Y(n_691) );
BUFx6f_ASAP7_75t_L g692 ( .A(n_585), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_625), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_605), .B(n_577), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g695 ( .A1(n_611), .A2(n_631), .B(n_608), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_622), .B(n_577), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_622), .B(n_577), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_587), .B(n_334), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_622), .B(n_568), .Y(n_699) );
AND2x4_ASAP7_75t_L g700 ( .A(n_588), .B(n_368), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_630), .B(n_355), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_625), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g703 ( .A1(n_628), .A2(n_514), .B(n_513), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_625), .Y(n_704) );
CKINVDCx5p33_ASAP7_75t_R g705 ( .A(n_659), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_664), .Y(n_706) );
AND2x4_ASAP7_75t_L g707 ( .A(n_660), .B(n_492), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_625), .Y(n_708) );
OR2x6_ASAP7_75t_SL g709 ( .A(n_620), .B(n_361), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_620), .A2(n_569), .B1(n_568), .B2(n_364), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_667), .Y(n_711) );
INVx3_ASAP7_75t_L g712 ( .A(n_653), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_667), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_664), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_623), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_601), .A2(n_569), .B1(n_568), .B2(n_364), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_623), .Y(n_717) );
BUFx5_ASAP7_75t_L g718 ( .A(n_583), .Y(n_718) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_585), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_621), .A2(n_569), .B1(n_568), .B2(n_410), .Y(n_720) );
INVx4_ASAP7_75t_L g721 ( .A(n_653), .Y(n_721) );
AOI33xp33_ASAP7_75t_L g722 ( .A1(n_594), .A2(n_514), .A3(n_530), .B1(n_513), .B2(n_404), .B3(n_337), .Y(n_722) );
INVx6_ASAP7_75t_L g723 ( .A(n_653), .Y(n_723) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_585), .Y(n_724) );
CKINVDCx5p33_ASAP7_75t_R g725 ( .A(n_633), .Y(n_725) );
OAI21x1_ASAP7_75t_SL g726 ( .A1(n_640), .A2(n_530), .B(n_466), .Y(n_726) );
BUFx2_ASAP7_75t_L g727 ( .A(n_632), .Y(n_727) );
OR2x2_ASAP7_75t_L g728 ( .A(n_647), .B(n_410), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_603), .A2(n_569), .B1(n_568), .B2(n_421), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_579), .Y(n_730) );
INVx3_ASAP7_75t_L g731 ( .A(n_653), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_579), .Y(n_732) );
AND2x4_ASAP7_75t_L g733 ( .A(n_612), .B(n_340), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_650), .A2(n_536), .B(n_535), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_624), .Y(n_735) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_634), .Y(n_736) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_585), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_595), .A2(n_569), .B1(n_568), .B2(n_452), .Y(n_738) );
INVx6_ASAP7_75t_L g739 ( .A(n_653), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_663), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_624), .Y(n_741) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_580), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_650), .A2(n_553), .B(n_536), .Y(n_743) );
INVx1_ASAP7_75t_SL g744 ( .A(n_580), .Y(n_744) );
AND2x2_ASAP7_75t_SL g745 ( .A(n_661), .B(n_370), .Y(n_745) );
BUFx6f_ASAP7_75t_L g746 ( .A(n_585), .Y(n_746) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_637), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_663), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_663), .Y(n_749) );
BUFx3_ASAP7_75t_L g750 ( .A(n_663), .Y(n_750) );
INVxp67_ASAP7_75t_SL g751 ( .A(n_663), .Y(n_751) );
INVx5_ASAP7_75t_L g752 ( .A(n_637), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_641), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_624), .Y(n_754) );
BUFx2_ASAP7_75t_L g755 ( .A(n_595), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_656), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_595), .B(n_569), .Y(n_757) );
AND2x4_ASAP7_75t_L g758 ( .A(n_612), .B(n_396), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_594), .A2(n_569), .B1(n_421), .B2(n_436), .Y(n_759) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_637), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_584), .Y(n_761) );
INVx1_ASAP7_75t_SL g762 ( .A(n_580), .Y(n_762) );
BUFx3_ASAP7_75t_L g763 ( .A(n_592), .Y(n_763) );
AND2x4_ASAP7_75t_L g764 ( .A(n_586), .B(n_405), .Y(n_764) );
NAND2x1p5_ASAP7_75t_L g765 ( .A(n_593), .B(n_376), .Y(n_765) );
INVx4_ASAP7_75t_L g766 ( .A(n_651), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_658), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_591), .Y(n_768) );
NOR2x1_ASAP7_75t_SL g769 ( .A(n_582), .B(n_397), .Y(n_769) );
BUFx4f_ASAP7_75t_L g770 ( .A(n_651), .Y(n_770) );
CKINVDCx5p33_ASAP7_75t_R g771 ( .A(n_649), .Y(n_771) );
AOI22xp33_ASAP7_75t_SL g772 ( .A1(n_598), .A2(n_569), .B1(n_452), .B2(n_462), .Y(n_772) );
A2O1A1Ixp33_ASAP7_75t_L g773 ( .A1(n_614), .A2(n_507), .B(n_515), .C(n_494), .Y(n_773) );
INVxp67_ASAP7_75t_L g774 ( .A(n_639), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_597), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_657), .B(n_428), .Y(n_776) );
INVx3_ASAP7_75t_L g777 ( .A(n_637), .Y(n_777) );
INVx3_ASAP7_75t_L g778 ( .A(n_637), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_618), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_629), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_614), .B(n_428), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_617), .B(n_436), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_604), .B(n_467), .Y(n_783) );
BUFx3_ASAP7_75t_L g784 ( .A(n_635), .Y(n_784) );
BUFx6f_ASAP7_75t_L g785 ( .A(n_589), .Y(n_785) );
BUFx6f_ASAP7_75t_L g786 ( .A(n_589), .Y(n_786) );
AND2x4_ASAP7_75t_L g787 ( .A(n_636), .B(n_406), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_643), .Y(n_788) );
INVx1_ASAP7_75t_SL g789 ( .A(n_661), .Y(n_789) );
OR2x6_ASAP7_75t_L g790 ( .A(n_655), .B(n_397), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_662), .Y(n_791) );
AND2x4_ASAP7_75t_L g792 ( .A(n_668), .B(n_413), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_669), .Y(n_793) );
BUFx6f_ASAP7_75t_L g794 ( .A(n_589), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_591), .Y(n_795) );
INVx3_ASAP7_75t_L g796 ( .A(n_600), .Y(n_796) );
HB1xp67_ASAP7_75t_L g797 ( .A(n_666), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_644), .A2(n_462), .B1(n_342), .B2(n_473), .Y(n_798) );
BUFx2_ASAP7_75t_L g799 ( .A(n_600), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_606), .Y(n_800) );
INVx4_ASAP7_75t_L g801 ( .A(n_589), .Y(n_801) );
BUFx2_ASAP7_75t_SL g802 ( .A(n_589), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_644), .A2(n_342), .B1(n_415), .B2(n_414), .Y(n_803) );
CKINVDCx11_ASAP7_75t_R g804 ( .A(n_652), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_606), .Y(n_805) );
AND2x4_ASAP7_75t_L g806 ( .A(n_638), .B(n_416), .Y(n_806) );
OAI22xp33_ASAP7_75t_L g807 ( .A1(n_670), .A2(n_467), .B1(n_471), .B2(n_469), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_670), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_701), .B(n_469), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_688), .A2(n_666), .B1(n_609), .B2(n_652), .Y(n_810) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_673), .Y(n_811) );
INVxp67_ASAP7_75t_L g812 ( .A(n_709), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_672), .Y(n_813) );
INVx2_ASAP7_75t_L g814 ( .A(n_768), .Y(n_814) );
O2A1O1Ixp33_ASAP7_75t_L g815 ( .A1(n_680), .A2(n_609), .B(n_422), .C(n_435), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_745), .A2(n_613), .B1(n_615), .B2(n_610), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_755), .B(n_610), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_795), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_774), .A2(n_615), .B1(n_627), .B2(n_613), .Y(n_819) );
CKINVDCx14_ASAP7_75t_R g820 ( .A(n_804), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_765), .Y(n_821) );
OR2x2_ASAP7_75t_L g822 ( .A(n_698), .B(n_471), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_774), .A2(n_627), .B1(n_596), .B2(n_359), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_800), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_783), .B(n_486), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_805), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_728), .B(n_486), .Y(n_827) );
CKINVDCx8_ASAP7_75t_R g828 ( .A(n_683), .Y(n_828) );
OAI22xp33_ASAP7_75t_L g829 ( .A1(n_679), .A2(n_682), .B1(n_759), .B2(n_676), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_796), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_679), .A2(n_515), .B1(n_528), .B2(n_507), .Y(n_831) );
INVx3_ASAP7_75t_L g832 ( .A(n_721), .Y(n_832) );
BUFx12f_ASAP7_75t_L g833 ( .A(n_674), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_679), .B(n_654), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_753), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_765), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_673), .A2(n_596), .B1(n_582), .B2(n_654), .Y(n_837) );
OAI21xp5_ASAP7_75t_L g838 ( .A1(n_703), .A2(n_596), .B(n_619), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_722), .B(n_638), .Y(n_839) );
OAI211xp5_ASAP7_75t_L g840 ( .A1(n_772), .A2(n_379), .B(n_441), .C(n_377), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_764), .B(n_377), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_796), .Y(n_842) );
OAI22xp33_ASAP7_75t_L g843 ( .A1(n_725), .A2(n_582), .B1(n_441), .B2(n_478), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_764), .A2(n_515), .B1(n_528), .B2(n_507), .Y(n_844) );
CKINVDCx5p33_ASAP7_75t_R g845 ( .A(n_705), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_799), .A2(n_675), .B1(n_687), .B2(n_681), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_797), .Y(n_847) );
INVx1_ASAP7_75t_SL g848 ( .A(n_675), .Y(n_848) );
O2A1O1Ixp33_ASAP7_75t_SL g849 ( .A1(n_773), .A2(n_335), .B(n_344), .C(n_341), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_681), .A2(n_619), .B1(n_602), .B2(n_599), .Y(n_850) );
AOI22x1_ASAP7_75t_L g851 ( .A1(n_726), .A2(n_519), .B1(n_522), .B2(n_499), .Y(n_851) );
INVx1_ASAP7_75t_SL g852 ( .A(n_806), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_756), .B(n_616), .Y(n_853) );
NOR2xp67_ASAP7_75t_SL g854 ( .A(n_802), .B(n_599), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_730), .Y(n_855) );
OAI22xp33_ASAP7_75t_L g856 ( .A1(n_720), .A2(n_478), .B1(n_481), .B2(n_379), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_689), .B(n_700), .Y(n_857) );
INVx4_ASAP7_75t_L g858 ( .A(n_752), .Y(n_858) );
INVx2_ASAP7_75t_L g859 ( .A(n_732), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_797), .Y(n_860) );
BUFx4_ASAP7_75t_SL g861 ( .A(n_790), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_787), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_689), .B(n_481), .Y(n_863) );
OR2x2_ASAP7_75t_L g864 ( .A(n_776), .B(n_482), .Y(n_864) );
OAI22xp33_ASAP7_75t_L g865 ( .A1(n_790), .A2(n_482), .B1(n_333), .B2(n_358), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_767), .A2(n_515), .B1(n_528), .B2(n_507), .Y(n_866) );
INVx2_ASAP7_75t_SL g867 ( .A(n_671), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_687), .B(n_616), .Y(n_868) );
INVxp67_ASAP7_75t_SL g869 ( .A(n_736), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_787), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_692), .Y(n_871) );
INVx2_ASAP7_75t_L g872 ( .A(n_692), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_694), .A2(n_602), .B1(n_599), .B2(n_333), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_772), .A2(n_515), .B1(n_528), .B2(n_507), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_771), .A2(n_343), .B1(n_369), .B2(n_358), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_792), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_806), .A2(n_515), .B1(n_528), .B2(n_507), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g878 ( .A(n_711), .B(n_418), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_792), .Y(n_879) );
AND2x4_ASAP7_75t_L g880 ( .A(n_713), .B(n_599), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_686), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_781), .A2(n_528), .B1(n_449), .B2(n_454), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_781), .A2(n_458), .B1(n_470), .B2(n_440), .Y(n_883) );
INVx1_ASAP7_75t_SL g884 ( .A(n_736), .Y(n_884) );
BUFx3_ASAP7_75t_L g885 ( .A(n_752), .Y(n_885) );
AOI21xp5_ASAP7_75t_L g886 ( .A1(n_734), .A2(n_602), .B(n_599), .Y(n_886) );
BUFx6f_ASAP7_75t_L g887 ( .A(n_692), .Y(n_887) );
AOI21xp5_ASAP7_75t_L g888 ( .A1(n_734), .A2(n_602), .B(n_616), .Y(n_888) );
BUFx3_ASAP7_75t_L g889 ( .A(n_752), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_694), .A2(n_602), .B1(n_343), .B2(n_385), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_719), .Y(n_891) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_790), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_686), .Y(n_893) );
AOI22xp5_ASAP7_75t_L g894 ( .A1(n_757), .A2(n_385), .B1(n_395), .B2(n_369), .Y(n_894) );
NAND2x1p5_ASAP7_75t_L g895 ( .A(n_752), .B(n_447), .Y(n_895) );
OAI22xp33_ASAP7_75t_L g896 ( .A1(n_696), .A2(n_395), .B1(n_448), .B2(n_444), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_695), .A2(n_472), .B1(n_453), .B2(n_447), .Y(n_897) );
INVx2_ASAP7_75t_L g898 ( .A(n_719), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_696), .A2(n_448), .B1(n_455), .B2(n_444), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_700), .B(n_453), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_697), .A2(n_455), .B1(n_423), .B2(n_331), .Y(n_901) );
OAI22xp33_ASAP7_75t_L g902 ( .A1(n_697), .A2(n_474), .B1(n_382), .B2(n_386), .Y(n_902) );
CKINVDCx5p33_ASAP7_75t_R g903 ( .A(n_727), .Y(n_903) );
NAND3xp33_ASAP7_75t_L g904 ( .A(n_695), .B(n_508), .C(n_349), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_733), .Y(n_905) );
OAI22x1_ASAP7_75t_L g906 ( .A1(n_729), .A2(n_387), .B1(n_389), .B2(n_357), .Y(n_906) );
AND2x4_ASAP7_75t_L g907 ( .A(n_684), .B(n_399), .Y(n_907) );
INVx2_ASAP7_75t_L g908 ( .A(n_719), .Y(n_908) );
BUFx6f_ASAP7_75t_L g909 ( .A(n_724), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g910 ( .A(n_776), .B(n_348), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_733), .Y(n_911) );
OAI22xp33_ASAP7_75t_L g912 ( .A1(n_710), .A2(n_429), .B1(n_437), .B2(n_411), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_758), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_724), .Y(n_914) );
OR2x6_ASAP7_75t_L g915 ( .A(n_766), .B(n_393), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_758), .A2(n_353), .B1(n_354), .B2(n_350), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_690), .A2(n_383), .B1(n_384), .B2(n_356), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_738), .A2(n_402), .B1(n_407), .B2(n_394), .Y(n_918) );
INVx2_ASAP7_75t_L g919 ( .A(n_724), .Y(n_919) );
AOI221xp5_ASAP7_75t_L g920 ( .A1(n_707), .A2(n_477), .B1(n_408), .B2(n_483), .C(n_409), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_775), .Y(n_921) );
AOI21xp33_ASAP7_75t_L g922 ( .A1(n_782), .A2(n_426), .B(n_419), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_779), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g924 ( .A(n_803), .B(n_427), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_780), .A2(n_434), .B1(n_442), .B2(n_433), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_788), .A2(n_443), .B1(n_450), .B2(n_445), .Y(n_926) );
AOI221xp5_ASAP7_75t_L g927 ( .A1(n_707), .A2(n_476), .B1(n_463), .B2(n_465), .C(n_487), .Y(n_927) );
BUFx3_ASAP7_75t_L g928 ( .A(n_785), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_791), .Y(n_929) );
AO21x1_ASAP7_75t_L g930 ( .A1(n_743), .A2(n_519), .B(n_499), .Y(n_930) );
NOR2xp33_ASAP7_75t_L g931 ( .A(n_757), .B(n_484), .Y(n_931) );
INVx2_ASAP7_75t_L g932 ( .A(n_737), .Y(n_932) );
HB1xp67_ASAP7_75t_L g933 ( .A(n_721), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_782), .B(n_6), .Y(n_934) );
AO31x2_ASAP7_75t_L g935 ( .A1(n_703), .A2(n_519), .A3(n_522), .B(n_499), .Y(n_935) );
CKINVDCx20_ASAP7_75t_R g936 ( .A(n_716), .Y(n_936) );
NOR2xp67_ASAP7_75t_SL g937 ( .A(n_766), .B(n_468), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g938 ( .A1(n_699), .A2(n_488), .B1(n_466), .B2(n_485), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_793), .Y(n_939) );
BUFx3_ASAP7_75t_L g940 ( .A(n_785), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_763), .A2(n_508), .B1(n_468), .B2(n_485), .Y(n_941) );
INVx2_ASAP7_75t_L g942 ( .A(n_737), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_798), .B(n_7), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_784), .A2(n_508), .B1(n_438), .B2(n_499), .Y(n_944) );
AOI22xp5_ASAP7_75t_L g945 ( .A1(n_699), .A2(n_508), .B1(n_438), .B2(n_536), .Y(n_945) );
INVx3_ASAP7_75t_L g946 ( .A(n_739), .Y(n_946) );
INVx2_ASAP7_75t_L g947 ( .A(n_737), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_685), .B(n_7), .Y(n_948) );
BUFx3_ASAP7_75t_L g949 ( .A(n_785), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_715), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_717), .A2(n_519), .B1(n_527), .B2(n_522), .Y(n_951) );
AO21x2_ASAP7_75t_L g952 ( .A1(n_677), .A2(n_527), .B(n_522), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_735), .A2(n_527), .B1(n_529), .B2(n_516), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_741), .A2(n_527), .B1(n_529), .B2(n_516), .Y(n_954) );
AOI22xp33_ASAP7_75t_SL g955 ( .A1(n_789), .A2(n_12), .B1(n_9), .B2(n_10), .Y(n_955) );
OAI21xp5_ASAP7_75t_L g956 ( .A1(n_743), .A2(n_761), .B(n_742), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_754), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_714), .A2(n_529), .B1(n_516), .B2(n_553), .Y(n_958) );
OR2x2_ASAP7_75t_L g959 ( .A(n_693), .B(n_9), .Y(n_959) );
OAI22xp33_ASAP7_75t_L g960 ( .A1(n_822), .A2(n_789), .B1(n_770), .B2(n_744), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_831), .A2(n_762), .B1(n_744), .B2(n_751), .Y(n_961) );
INVx2_ASAP7_75t_L g962 ( .A(n_814), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_814), .Y(n_963) );
AND2x2_ASAP7_75t_L g964 ( .A(n_857), .B(n_702), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_831), .A2(n_762), .B1(n_751), .B2(n_770), .Y(n_965) );
OAI22xp33_ASAP7_75t_L g966 ( .A1(n_812), .A2(n_816), .B1(n_848), .B2(n_903), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_916), .A2(n_739), .B1(n_742), .B2(n_723), .Y(n_967) );
AOI221xp5_ASAP7_75t_L g968 ( .A1(n_863), .A2(n_708), .B1(n_704), .B2(n_691), .C(n_706), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_936), .A2(n_750), .B1(n_740), .B2(n_749), .Y(n_969) );
OR2x6_ASAP7_75t_L g970 ( .A(n_915), .B(n_739), .Y(n_970) );
AOI22xp33_ASAP7_75t_SL g971 ( .A1(n_820), .A2(n_769), .B1(n_723), .B2(n_801), .Y(n_971) );
OAI21x1_ASAP7_75t_L g972 ( .A1(n_888), .A2(n_778), .B(n_777), .Y(n_972) );
OAI22xp5_ASAP7_75t_L g973 ( .A1(n_916), .A2(n_874), .B1(n_823), .B2(n_808), .Y(n_973) );
INVx2_ASAP7_75t_L g974 ( .A(n_818), .Y(n_974) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_807), .A2(n_678), .B1(n_731), .B2(n_712), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_825), .B(n_712), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_813), .Y(n_977) );
OAI21xp33_ASAP7_75t_L g978 ( .A1(n_910), .A2(n_748), .B(n_731), .Y(n_978) );
AOI22xp33_ASAP7_75t_SL g979 ( .A1(n_820), .A2(n_801), .B1(n_794), .B2(n_786), .Y(n_979) );
OAI22xp33_ASAP7_75t_L g980 ( .A1(n_884), .A2(n_794), .B1(n_786), .B2(n_746), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_841), .B(n_718), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_883), .B(n_718), .Y(n_982) );
OAI221xp5_ASAP7_75t_L g983 ( .A1(n_920), .A2(n_778), .B1(n_777), .B2(n_794), .C(n_786), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_809), .B(n_10), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_921), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_943), .A2(n_874), .B1(n_910), .B2(n_829), .Y(n_986) );
AOI222xp33_ASAP7_75t_L g987 ( .A1(n_827), .A2(n_529), .B1(n_747), .B2(n_746), .C1(n_760), .C2(n_516), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_934), .A2(n_718), .B1(n_747), .B2(n_746), .Y(n_988) );
AOI21xp33_ASAP7_75t_L g989 ( .A1(n_815), .A2(n_760), .B(n_747), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_922), .A2(n_718), .B1(n_760), .B2(n_516), .Y(n_990) );
OAI21xp33_ASAP7_75t_L g991 ( .A1(n_897), .A2(n_556), .B(n_553), .Y(n_991) );
AOI221xp5_ASAP7_75t_L g992 ( .A1(n_900), .A2(n_516), .B1(n_562), .B2(n_571), .C(n_567), .Y(n_992) );
NOR2x1_ASAP7_75t_SL g993 ( .A(n_915), .B(n_718), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_883), .B(n_13), .Y(n_994) );
OA21x2_ASAP7_75t_L g995 ( .A1(n_930), .A2(n_562), .B(n_556), .Y(n_995) );
BUFx2_ASAP7_75t_L g996 ( .A(n_869), .Y(n_996) );
AOI221xp5_ASAP7_75t_L g997 ( .A1(n_878), .A2(n_516), .B1(n_571), .B2(n_567), .C(n_565), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_846), .A2(n_554), .B1(n_540), .B2(n_15), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_923), .B(n_13), .Y(n_999) );
AOI221xp5_ASAP7_75t_L g1000 ( .A1(n_878), .A2(n_562), .B1(n_571), .B2(n_567), .C(n_565), .Y(n_1000) );
INVx1_ASAP7_75t_SL g1001 ( .A(n_861), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_931), .A2(n_554), .B1(n_540), .B2(n_17), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_844), .B(n_14), .Y(n_1003) );
AOI22xp33_ASAP7_75t_SL g1004 ( .A1(n_892), .A2(n_17), .B1(n_14), .B2(n_16), .Y(n_1004) );
NAND2x1p5_ASAP7_75t_L g1005 ( .A(n_858), .B(n_573), .Y(n_1005) );
INVx2_ASAP7_75t_L g1006 ( .A(n_818), .Y(n_1006) );
HB1xp67_ASAP7_75t_L g1007 ( .A(n_828), .Y(n_1007) );
OAI21xp5_ASAP7_75t_L g1008 ( .A1(n_853), .A2(n_565), .B(n_556), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_931), .A2(n_554), .B1(n_540), .B2(n_21), .Y(n_1009) );
CKINVDCx20_ASAP7_75t_R g1010 ( .A(n_833), .Y(n_1010) );
AOI222xp33_ASAP7_75t_L g1011 ( .A1(n_927), .A2(n_16), .B1(n_19), .B2(n_22), .C1(n_23), .C2(n_24), .Y(n_1011) );
OAI22xp33_ASAP7_75t_L g1012 ( .A1(n_821), .A2(n_25), .B1(n_22), .B2(n_23), .Y(n_1012) );
HB1xp67_ASAP7_75t_L g1013 ( .A(n_836), .Y(n_1013) );
OAI33xp33_ASAP7_75t_L g1014 ( .A1(n_856), .A2(n_26), .A3(n_27), .B1(n_28), .B2(n_29), .B3(n_30), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_844), .B(n_27), .Y(n_1015) );
INVx2_ASAP7_75t_SL g1016 ( .A(n_885), .Y(n_1016) );
AOI22xp33_ASAP7_75t_SL g1017 ( .A1(n_840), .A2(n_31), .B1(n_28), .B2(n_29), .Y(n_1017) );
AOI221xp5_ASAP7_75t_L g1018 ( .A1(n_843), .A2(n_554), .B1(n_540), .B2(n_573), .C(n_35), .Y(n_1018) );
AOI22xp33_ASAP7_75t_SL g1019 ( .A1(n_915), .A2(n_34), .B1(n_32), .B2(n_33), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_875), .B(n_32), .Y(n_1020) );
AOI22xp33_ASAP7_75t_SL g1021 ( .A1(n_811), .A2(n_35), .B1(n_33), .B2(n_34), .Y(n_1021) );
AOI21xp33_ASAP7_75t_L g1022 ( .A1(n_839), .A2(n_36), .B(n_37), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_905), .A2(n_540), .B1(n_554), .B2(n_39), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_929), .Y(n_1024) );
INVx2_ASAP7_75t_SL g1025 ( .A(n_885), .Y(n_1025) );
OR2x2_ASAP7_75t_L g1026 ( .A(n_864), .B(n_36), .Y(n_1026) );
NOR2xp33_ASAP7_75t_L g1027 ( .A(n_862), .B(n_38), .Y(n_1027) );
INVx1_ASAP7_75t_SL g1028 ( .A(n_889), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_939), .B(n_39), .Y(n_1029) );
OAI22xp33_ASAP7_75t_L g1030 ( .A1(n_865), .A2(n_40), .B1(n_41), .B2(n_42), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_870), .B(n_40), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_881), .B(n_41), .Y(n_1032) );
OAI211xp5_ASAP7_75t_L g1033 ( .A1(n_918), .A2(n_554), .B(n_540), .C(n_573), .Y(n_1033) );
BUFx6f_ASAP7_75t_L g1034 ( .A(n_887), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_893), .B(n_42), .Y(n_1035) );
AOI22xp33_ASAP7_75t_SL g1036 ( .A1(n_852), .A2(n_43), .B1(n_45), .B2(n_46), .Y(n_1036) );
HB1xp67_ASAP7_75t_L g1037 ( .A(n_933), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_847), .Y(n_1038) );
OAI21xp5_ASAP7_75t_L g1039 ( .A1(n_868), .A2(n_573), .B(n_43), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_824), .Y(n_1040) );
AOI221xp5_ASAP7_75t_L g1041 ( .A1(n_897), .A2(n_554), .B1(n_540), .B2(n_51), .C(n_52), .Y(n_1041) );
OAI22xp5_ASAP7_75t_L g1042 ( .A1(n_819), .A2(n_49), .B1(n_50), .B2(n_52), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_876), .B(n_53), .Y(n_1043) );
INVx2_ASAP7_75t_L g1044 ( .A(n_824), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_879), .B(n_53), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_860), .Y(n_1046) );
OAI21x1_ASAP7_75t_L g1047 ( .A1(n_851), .A2(n_118), .B(n_112), .Y(n_1047) );
OAI22xp33_ASAP7_75t_L g1048 ( .A1(n_911), .A2(n_56), .B1(n_57), .B2(n_58), .Y(n_1048) );
OAI211xp5_ASAP7_75t_L g1049 ( .A1(n_918), .A2(n_57), .B(n_59), .C(n_60), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_913), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_882), .A2(n_62), .B1(n_63), .B2(n_64), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_948), .Y(n_1052) );
NAND2x1p5_ASAP7_75t_L g1053 ( .A(n_858), .B(n_63), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_899), .B(n_64), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_917), .A2(n_66), .B1(n_67), .B2(n_70), .Y(n_1055) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_889), .Y(n_1056) );
INVx2_ASAP7_75t_L g1057 ( .A(n_826), .Y(n_1057) );
AO21x2_ASAP7_75t_L g1058 ( .A1(n_952), .A2(n_904), .B(n_838), .Y(n_1058) );
OR2x2_ASAP7_75t_L g1059 ( .A(n_901), .B(n_66), .Y(n_1059) );
BUFx3_ASAP7_75t_L g1060 ( .A(n_928), .Y(n_1060) );
NAND3xp33_ASAP7_75t_L g1061 ( .A(n_882), .B(n_67), .C(n_71), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_817), .A2(n_71), .B1(n_72), .B2(n_74), .Y(n_1062) );
OAI211xp5_ASAP7_75t_L g1063 ( .A1(n_955), .A2(n_72), .B(n_74), .C(n_75), .Y(n_1063) );
AOI222xp33_ASAP7_75t_L g1064 ( .A1(n_833), .A2(n_75), .B1(n_76), .B2(n_77), .C1(n_78), .C2(n_79), .Y(n_1064) );
AO21x2_ASAP7_75t_L g1065 ( .A1(n_952), .A2(n_121), .B(n_120), .Y(n_1065) );
OAI22xp33_ASAP7_75t_L g1066 ( .A1(n_959), .A2(n_76), .B1(n_78), .B2(n_79), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_817), .B(n_925), .Y(n_1067) );
AO21x2_ASAP7_75t_L g1068 ( .A1(n_956), .A2(n_124), .B(n_122), .Y(n_1068) );
OAI21x1_ASAP7_75t_L g1069 ( .A1(n_886), .A2(n_126), .B(n_125), .Y(n_1069) );
AOI22xp5_ASAP7_75t_L g1070 ( .A1(n_896), .A2(n_80), .B1(n_81), .B2(n_82), .Y(n_1070) );
AO21x2_ASAP7_75t_L g1071 ( .A1(n_849), .A2(n_131), .B(n_127), .Y(n_1071) );
OAI21xp5_ASAP7_75t_L g1072 ( .A1(n_810), .A2(n_80), .B(n_82), .Y(n_1072) );
INVx2_ASAP7_75t_L g1073 ( .A(n_826), .Y(n_1073) );
HB1xp67_ASAP7_75t_L g1074 ( .A(n_834), .Y(n_1074) );
OR2x2_ASAP7_75t_L g1075 ( .A(n_924), .B(n_83), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_925), .B(n_85), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_950), .Y(n_1077) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_917), .A2(n_810), .B1(n_877), .B2(n_926), .Y(n_1078) );
OAI221xp5_ASAP7_75t_SL g1079 ( .A1(n_926), .A2(n_86), .B1(n_87), .B2(n_88), .C(n_89), .Y(n_1079) );
A2O1A1Ixp33_ASAP7_75t_L g1080 ( .A1(n_855), .A2(n_86), .B(n_89), .C(n_90), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_877), .B(n_91), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_906), .A2(n_92), .B1(n_93), .B2(n_94), .Y(n_1082) );
OAI22xp5_ASAP7_75t_L g1083 ( .A1(n_895), .A2(n_92), .B1(n_93), .B2(n_94), .Y(n_1083) );
AOI221xp5_ASAP7_75t_L g1084 ( .A1(n_912), .A2(n_95), .B1(n_96), .B2(n_97), .C(n_98), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_938), .A2(n_95), .B1(n_97), .B2(n_99), .Y(n_1085) );
INVx3_ASAP7_75t_L g1086 ( .A(n_928), .Y(n_1086) );
OAI221xp5_ASAP7_75t_SL g1087 ( .A1(n_902), .A2(n_99), .B1(n_100), .B2(n_102), .C(n_103), .Y(n_1087) );
CKINVDCx5p33_ASAP7_75t_R g1088 ( .A(n_845), .Y(n_1088) );
AOI221xp5_ASAP7_75t_L g1089 ( .A1(n_849), .A2(n_100), .B1(n_104), .B2(n_106), .C(n_132), .Y(n_1089) );
BUFx2_ASAP7_75t_L g1090 ( .A(n_895), .Y(n_1090) );
INVx2_ASAP7_75t_L g1091 ( .A(n_935), .Y(n_1091) );
INVx2_ASAP7_75t_L g1092 ( .A(n_935), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_957), .B(n_136), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_866), .A2(n_137), .B1(n_138), .B2(n_139), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_907), .Y(n_1095) );
NOR4xp25_ASAP7_75t_L g1096 ( .A(n_866), .B(n_140), .C(n_141), .D(n_143), .Y(n_1096) );
AND2x4_ASAP7_75t_L g1097 ( .A(n_940), .B(n_949), .Y(n_1097) );
BUFx4f_ASAP7_75t_SL g1098 ( .A(n_835), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_907), .A2(n_146), .B1(n_148), .B2(n_149), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_941), .A2(n_150), .B1(n_151), .B2(n_154), .Y(n_1100) );
INVx2_ASAP7_75t_L g1101 ( .A(n_935), .Y(n_1101) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_996), .B(n_832), .Y(n_1102) );
AOI22xp33_ASAP7_75t_SL g1103 ( .A1(n_993), .A2(n_832), .B1(n_837), .B2(n_940), .Y(n_1103) );
HB1xp67_ASAP7_75t_L g1104 ( .A(n_1037), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_985), .Y(n_1105) );
INVx4_ASAP7_75t_L g1106 ( .A(n_970), .Y(n_1106) );
INVx2_ASAP7_75t_L g1107 ( .A(n_962), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_962), .B(n_855), .Y(n_1108) );
AO21x2_ASAP7_75t_L g1109 ( .A1(n_1039), .A2(n_945), .B(n_872), .Y(n_1109) );
OAI33xp33_ASAP7_75t_L g1110 ( .A1(n_1030), .A2(n_890), .A3(n_873), .B1(n_850), .B2(n_830), .B3(n_842), .Y(n_1110) );
OR2x2_ASAP7_75t_L g1111 ( .A(n_1026), .B(n_859), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1024), .Y(n_1112) );
INVx3_ASAP7_75t_L g1113 ( .A(n_1034), .Y(n_1113) );
OA21x2_ASAP7_75t_L g1114 ( .A1(n_1091), .A2(n_954), .B(n_953), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_977), .Y(n_1115) );
AOI221xp5_ASAP7_75t_L g1116 ( .A1(n_1087), .A2(n_867), .B1(n_941), .B2(n_937), .C(n_944), .Y(n_1116) );
AOI211xp5_ASAP7_75t_L g1117 ( .A1(n_966), .A2(n_894), .B(n_880), .C(n_946), .Y(n_1117) );
OAI21x1_ASAP7_75t_L g1118 ( .A1(n_972), .A2(n_872), .B(n_871), .Y(n_1118) );
INVxp67_ASAP7_75t_L g1119 ( .A(n_1013), .Y(n_1119) );
INVx2_ASAP7_75t_L g1120 ( .A(n_963), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_986), .A2(n_830), .B1(n_842), .B2(n_859), .Y(n_1121) );
AOI221xp5_ASAP7_75t_L g1122 ( .A1(n_1079), .A2(n_944), .B1(n_951), .B2(n_953), .C(n_954), .Y(n_1122) );
INVx3_ASAP7_75t_L g1123 ( .A(n_1034), .Y(n_1123) );
OAI221xp5_ASAP7_75t_L g1124 ( .A1(n_986), .A2(n_951), .B1(n_958), .B2(n_946), .C(n_949), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_964), .B(n_935), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_963), .B(n_871), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1077), .Y(n_1127) );
INVx2_ASAP7_75t_L g1128 ( .A(n_974), .Y(n_1128) );
NAND3xp33_ASAP7_75t_L g1129 ( .A(n_1082), .B(n_958), .C(n_880), .Y(n_1129) );
INVx2_ASAP7_75t_L g1130 ( .A(n_974), .Y(n_1130) );
OAI22xp33_ASAP7_75t_L g1131 ( .A1(n_1053), .A2(n_887), .B1(n_909), .B2(n_947), .Y(n_1131) );
AOI211xp5_ASAP7_75t_SL g1132 ( .A1(n_960), .A2(n_880), .B(n_942), .C(n_932), .Y(n_1132) );
AOI221x1_ASAP7_75t_SL g1133 ( .A1(n_1012), .A2(n_947), .B1(n_942), .B2(n_932), .C(n_919), .Y(n_1133) );
OR2x2_ASAP7_75t_L g1134 ( .A(n_1028), .B(n_891), .Y(n_1134) );
AOI22xp33_ASAP7_75t_SL g1135 ( .A1(n_1053), .A2(n_1067), .B1(n_973), .B2(n_1076), .Y(n_1135) );
BUFx3_ASAP7_75t_L g1136 ( .A(n_1090), .Y(n_1136) );
AOI22xp5_ASAP7_75t_L g1137 ( .A1(n_1078), .A2(n_854), .B1(n_914), .B2(n_908), .Y(n_1137) );
AOI221xp5_ASAP7_75t_L g1138 ( .A1(n_1084), .A2(n_919), .B1(n_914), .B2(n_908), .C(n_898), .Y(n_1138) );
OAI211xp5_ASAP7_75t_SL g1139 ( .A1(n_1064), .A2(n_898), .B(n_891), .C(n_160), .Y(n_1139) );
OR2x2_ASAP7_75t_L g1140 ( .A(n_984), .B(n_887), .Y(n_1140) );
OAI221xp5_ASAP7_75t_L g1141 ( .A1(n_1019), .A2(n_909), .B1(n_887), .B2(n_163), .C(n_164), .Y(n_1141) );
INVx2_ASAP7_75t_L g1142 ( .A(n_1006), .Y(n_1142) );
AOI21xp5_ASAP7_75t_L g1143 ( .A1(n_1058), .A2(n_909), .B(n_159), .Y(n_1143) );
AOI221xp5_ASAP7_75t_L g1144 ( .A1(n_1014), .A2(n_909), .B1(n_166), .B2(n_167), .C(n_172), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_1081), .A2(n_158), .B1(n_173), .B2(n_174), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1146 ( .A(n_1038), .B(n_329), .Y(n_1146) );
AOI21xp5_ASAP7_75t_SL g1147 ( .A1(n_1072), .A2(n_175), .B(n_176), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1006), .B(n_177), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1046), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1040), .B(n_179), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_999), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1029), .Y(n_1152) );
OAI221xp5_ASAP7_75t_L g1153 ( .A1(n_1017), .A2(n_181), .B1(n_183), .B2(n_185), .C(n_186), .Y(n_1153) );
OA21x2_ASAP7_75t_L g1154 ( .A1(n_1091), .A2(n_187), .B(n_189), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_1003), .A2(n_190), .B1(n_191), .B2(n_192), .Y(n_1155) );
BUFx3_ASAP7_75t_L g1156 ( .A(n_1060), .Y(n_1156) );
AOI221xp5_ASAP7_75t_L g1157 ( .A1(n_1027), .A2(n_1048), .B1(n_1066), .B2(n_1055), .C(n_1095), .Y(n_1157) );
OAI31xp33_ASAP7_75t_L g1158 ( .A1(n_1063), .A2(n_194), .A3(n_198), .B(n_200), .Y(n_1158) );
OAI33xp33_ASAP7_75t_L g1159 ( .A1(n_1083), .A2(n_202), .A3(n_203), .B1(n_205), .B2(n_206), .B3(n_207), .Y(n_1159) );
HB1xp67_ASAP7_75t_L g1160 ( .A(n_1056), .Y(n_1160) );
OAI221xp5_ASAP7_75t_L g1161 ( .A1(n_1082), .A2(n_210), .B1(n_211), .B2(n_212), .C(n_214), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1043), .Y(n_1162) );
OAI22xp5_ASAP7_75t_L g1163 ( .A1(n_1002), .A2(n_215), .B1(n_218), .B2(n_219), .Y(n_1163) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1040), .Y(n_1164) );
AOI22xp33_ASAP7_75t_L g1165 ( .A1(n_1015), .A2(n_223), .B1(n_224), .B2(n_225), .Y(n_1165) );
HB1xp67_ASAP7_75t_L g1166 ( .A(n_1032), .Y(n_1166) );
BUFx3_ASAP7_75t_L g1167 ( .A(n_1060), .Y(n_1167) );
INVxp67_ASAP7_75t_L g1168 ( .A(n_1007), .Y(n_1168) );
OAI22xp5_ASAP7_75t_L g1169 ( .A1(n_1002), .A2(n_228), .B1(n_229), .B2(n_230), .Y(n_1169) );
BUFx2_ASAP7_75t_L g1170 ( .A(n_1016), .Y(n_1170) );
OA21x2_ASAP7_75t_L g1171 ( .A1(n_1092), .A2(n_231), .B(n_233), .Y(n_1171) );
AO21x2_ASAP7_75t_L g1172 ( .A1(n_1058), .A2(n_241), .B(n_242), .Y(n_1172) );
OR2x2_ASAP7_75t_L g1173 ( .A(n_1074), .B(n_243), .Y(n_1173) );
OAI221xp5_ASAP7_75t_SL g1174 ( .A1(n_1062), .A2(n_245), .B1(n_246), .B2(n_247), .C(n_248), .Y(n_1174) );
AOI221xp5_ASAP7_75t_L g1175 ( .A1(n_1027), .A2(n_251), .B1(n_252), .B2(n_253), .C(n_254), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g1176 ( .A1(n_1052), .A2(n_255), .B1(n_257), .B2(n_259), .Y(n_1176) );
BUFx2_ASAP7_75t_L g1177 ( .A(n_1016), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1020), .B(n_261), .Y(n_1178) );
AOI22xp5_ASAP7_75t_L g1179 ( .A1(n_1054), .A2(n_262), .B1(n_264), .B2(n_265), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1045), .Y(n_1180) );
NOR2xp33_ASAP7_75t_L g1181 ( .A(n_981), .B(n_266), .Y(n_1181) );
AOI21xp33_ASAP7_75t_L g1182 ( .A1(n_987), .A2(n_267), .B(n_268), .Y(n_1182) );
BUFx3_ASAP7_75t_L g1183 ( .A(n_1097), .Y(n_1183) );
AOI22xp33_ASAP7_75t_SL g1184 ( .A1(n_1049), .A2(n_270), .B1(n_271), .B2(n_273), .Y(n_1184) );
NAND3xp33_ASAP7_75t_L g1185 ( .A(n_1011), .B(n_274), .C(n_276), .Y(n_1185) );
NOR2x1_ASAP7_75t_L g1186 ( .A(n_1010), .B(n_277), .Y(n_1186) );
AOI21x1_ASAP7_75t_L g1187 ( .A1(n_995), .A2(n_328), .B(n_279), .Y(n_1187) );
AO21x2_ASAP7_75t_L g1188 ( .A1(n_1092), .A2(n_1101), .B(n_972), .Y(n_1188) );
INVx2_ASAP7_75t_L g1189 ( .A(n_1044), .Y(n_1189) );
OAI221xp5_ASAP7_75t_L g1190 ( .A1(n_1004), .A2(n_278), .B1(n_280), .B2(n_282), .C(n_285), .Y(n_1190) );
HB1xp67_ASAP7_75t_L g1191 ( .A(n_1035), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1031), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1075), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1194 ( .A(n_1001), .B(n_326), .Y(n_1194) );
AO21x2_ASAP7_75t_L g1195 ( .A1(n_1101), .A2(n_286), .B(n_287), .Y(n_1195) );
OAI211xp5_ASAP7_75t_SL g1196 ( .A1(n_1021), .A2(n_288), .B(n_290), .C(n_291), .Y(n_1196) );
AOI33xp33_ASAP7_75t_L g1197 ( .A1(n_1062), .A2(n_1051), .A3(n_1050), .B1(n_1036), .B2(n_1085), .B3(n_976), .Y(n_1197) );
INVx2_ASAP7_75t_L g1198 ( .A(n_1044), .Y(n_1198) );
AOI222xp33_ASAP7_75t_L g1199 ( .A1(n_1098), .A2(n_293), .B1(n_295), .B2(n_296), .C1(n_297), .C2(n_299), .Y(n_1199) );
AOI33xp33_ASAP7_75t_L g1200 ( .A1(n_1051), .A2(n_300), .A3(n_304), .B1(n_305), .B2(n_307), .B3(n_308), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1057), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1057), .Y(n_1202) );
OR2x2_ASAP7_75t_L g1203 ( .A(n_1059), .B(n_325), .Y(n_1203) );
OAI21xp5_ASAP7_75t_L g1204 ( .A1(n_1018), .A2(n_998), .B(n_1009), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1073), .Y(n_1205) );
BUFx2_ASAP7_75t_L g1206 ( .A(n_1025), .Y(n_1206) );
NOR2x1_ASAP7_75t_R g1207 ( .A(n_1088), .B(n_309), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1073), .B(n_311), .Y(n_1208) );
BUFx6f_ASAP7_75t_L g1209 ( .A(n_1034), .Y(n_1209) );
HB1xp67_ASAP7_75t_L g1210 ( .A(n_1025), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1080), .B(n_312), .Y(n_1211) );
AOI22xp33_ASAP7_75t_L g1212 ( .A1(n_994), .A2(n_314), .B1(n_315), .B2(n_319), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1042), .Y(n_1213) );
OAI221xp5_ASAP7_75t_L g1214 ( .A1(n_1085), .A2(n_321), .B1(n_324), .B2(n_1070), .C(n_998), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1061), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1201), .Y(n_1216) );
HB1xp67_ASAP7_75t_L g1217 ( .A(n_1104), .Y(n_1217) );
NAND2xp5_ASAP7_75t_SL g1218 ( .A(n_1131), .B(n_980), .Y(n_1218) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1107), .Y(n_1219) );
OR2x2_ASAP7_75t_L g1220 ( .A(n_1125), .B(n_982), .Y(n_1220) );
AND2x4_ASAP7_75t_L g1221 ( .A(n_1106), .B(n_1086), .Y(n_1221) );
BUFx6f_ASAP7_75t_L g1222 ( .A(n_1209), .Y(n_1222) );
OAI33xp33_ASAP7_75t_L g1223 ( .A1(n_1119), .A2(n_967), .A3(n_1100), .B1(n_961), .B2(n_1093), .B3(n_1088), .Y(n_1223) );
AOI22xp5_ASAP7_75t_L g1224 ( .A1(n_1135), .A2(n_1050), .B1(n_968), .B2(n_983), .Y(n_1224) );
AOI21xp33_ASAP7_75t_L g1225 ( .A1(n_1215), .A2(n_970), .B(n_969), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1108), .B(n_995), .Y(n_1226) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1107), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1108), .B(n_995), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1149), .Y(n_1229) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1120), .Y(n_1230) );
NAND3xp33_ASAP7_75t_L g1231 ( .A(n_1199), .B(n_1080), .C(n_1022), .Y(n_1231) );
NOR3xp33_ASAP7_75t_SL g1232 ( .A(n_1139), .B(n_1010), .C(n_1098), .Y(n_1232) );
AND4x1_ASAP7_75t_L g1233 ( .A(n_1186), .B(n_1089), .C(n_1099), .D(n_1009), .Y(n_1233) );
INVx2_ASAP7_75t_L g1234 ( .A(n_1120), .Y(n_1234) );
INVx2_ASAP7_75t_L g1235 ( .A(n_1128), .Y(n_1235) );
INVx4_ASAP7_75t_L g1236 ( .A(n_1106), .Y(n_1236) );
AOI221xp5_ASAP7_75t_L g1237 ( .A1(n_1193), .A2(n_1041), .B1(n_1096), .B2(n_1023), .C(n_992), .Y(n_1237) );
OR2x2_ASAP7_75t_L g1238 ( .A(n_1160), .B(n_969), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1105), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1128), .B(n_1008), .Y(n_1240) );
INVx2_ASAP7_75t_L g1241 ( .A(n_1130), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1130), .B(n_1086), .Y(n_1242) );
AOI22xp33_ASAP7_75t_L g1243 ( .A1(n_1185), .A2(n_970), .B1(n_978), .B2(n_1023), .Y(n_1243) );
INVx3_ASAP7_75t_L g1244 ( .A(n_1209), .Y(n_1244) );
OR2x2_ASAP7_75t_L g1245 ( .A(n_1111), .B(n_1086), .Y(n_1245) );
INVx2_ASAP7_75t_L g1246 ( .A(n_1142), .Y(n_1246) );
INVx2_ASAP7_75t_SL g1247 ( .A(n_1156), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1142), .B(n_1065), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1164), .B(n_1065), .Y(n_1249) );
INVx2_ASAP7_75t_SL g1250 ( .A(n_1156), .Y(n_1250) );
OAI21xp33_ASAP7_75t_L g1251 ( .A1(n_1211), .A2(n_1099), .B(n_1094), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1164), .B(n_1097), .Y(n_1252) );
OAI21xp5_ASAP7_75t_L g1253 ( .A1(n_1129), .A2(n_975), .B(n_990), .Y(n_1253) );
OR2x2_ASAP7_75t_L g1254 ( .A(n_1102), .B(n_970), .Y(n_1254) );
INVx2_ASAP7_75t_L g1255 ( .A(n_1189), .Y(n_1255) );
HB1xp67_ASAP7_75t_L g1256 ( .A(n_1210), .Y(n_1256) );
AOI221xp5_ASAP7_75t_L g1257 ( .A1(n_1151), .A2(n_979), .B1(n_997), .B2(n_971), .C(n_1000), .Y(n_1257) );
OAI222xp33_ASAP7_75t_L g1258 ( .A1(n_1106), .A2(n_1094), .B1(n_990), .B2(n_965), .C1(n_1097), .C2(n_988), .Y(n_1258) );
OAI221xp5_ASAP7_75t_L g1259 ( .A1(n_1157), .A2(n_988), .B1(n_989), .B2(n_991), .C(n_1033), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1112), .B(n_1071), .Y(n_1260) );
AND2x4_ASAP7_75t_L g1261 ( .A(n_1183), .B(n_1034), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1262 ( .A(n_1189), .B(n_1068), .Y(n_1262) );
NOR2xp33_ASAP7_75t_R g1263 ( .A(n_1136), .B(n_1005), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1202), .Y(n_1264) );
OAI33xp33_ASAP7_75t_L g1265 ( .A1(n_1168), .A2(n_1071), .A3(n_1068), .B1(n_1069), .B2(n_1047), .B3(n_1005), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1198), .B(n_1069), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1115), .B(n_1047), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1198), .B(n_1205), .Y(n_1268) );
AOI221xp5_ASAP7_75t_L g1269 ( .A1(n_1152), .A2(n_1192), .B1(n_1180), .B2(n_1162), .C(n_1213), .Y(n_1269) );
HB1xp67_ASAP7_75t_L g1270 ( .A(n_1170), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1127), .Y(n_1271) );
HB1xp67_ASAP7_75t_L g1272 ( .A(n_1177), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1166), .B(n_1191), .Y(n_1273) );
AOI21x1_ASAP7_75t_L g1274 ( .A1(n_1187), .A2(n_1143), .B(n_1154), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1188), .Y(n_1275) );
OAI33xp33_ASAP7_75t_L g1276 ( .A1(n_1203), .A2(n_1194), .A3(n_1178), .B1(n_1173), .B2(n_1146), .B3(n_1163), .Y(n_1276) );
NOR3xp33_ASAP7_75t_L g1277 ( .A(n_1207), .B(n_1116), .C(n_1141), .Y(n_1277) );
OAI221xp5_ASAP7_75t_L g1278 ( .A1(n_1133), .A2(n_1117), .B1(n_1204), .B2(n_1121), .C(n_1214), .Y(n_1278) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1134), .Y(n_1279) );
INVx2_ASAP7_75t_L g1280 ( .A(n_1188), .Y(n_1280) );
AOI211xp5_ASAP7_75t_SL g1281 ( .A1(n_1147), .A2(n_1174), .B(n_1131), .C(n_1190), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1126), .B(n_1121), .Y(n_1282) );
NOR2x1_ASAP7_75t_L g1283 ( .A(n_1136), .B(n_1167), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1206), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1126), .B(n_1148), .Y(n_1285) );
AO21x2_ASAP7_75t_L g1286 ( .A1(n_1172), .A2(n_1118), .B(n_1137), .Y(n_1286) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1173), .Y(n_1287) );
OAI31xp33_ASAP7_75t_L g1288 ( .A1(n_1132), .A2(n_1211), .A3(n_1161), .B(n_1196), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1148), .B(n_1150), .Y(n_1289) );
OAI22xp5_ASAP7_75t_L g1290 ( .A1(n_1145), .A2(n_1165), .B1(n_1155), .B2(n_1176), .Y(n_1290) );
AOI22xp33_ASAP7_75t_L g1291 ( .A1(n_1110), .A2(n_1124), .B1(n_1159), .B2(n_1122), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1150), .B(n_1208), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1208), .B(n_1183), .Y(n_1293) );
INVx2_ASAP7_75t_SL g1294 ( .A(n_1167), .Y(n_1294) );
AOI211xp5_ASAP7_75t_L g1295 ( .A1(n_1147), .A2(n_1153), .B(n_1182), .C(n_1169), .Y(n_1295) );
AOI22xp33_ASAP7_75t_L g1296 ( .A1(n_1181), .A2(n_1175), .B1(n_1109), .B2(n_1145), .Y(n_1296) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1140), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1113), .B(n_1123), .Y(n_1298) );
AOI211xp5_ASAP7_75t_SL g1299 ( .A1(n_1181), .A2(n_1179), .B(n_1144), .C(n_1113), .Y(n_1299) );
NAND3xp33_ASAP7_75t_L g1300 ( .A(n_1200), .B(n_1197), .C(n_1158), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1113), .B(n_1123), .Y(n_1301) );
OAI22xp5_ASAP7_75t_L g1302 ( .A1(n_1155), .A2(n_1165), .B1(n_1176), .B2(n_1103), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1123), .B(n_1209), .Y(n_1303) );
OR2x2_ASAP7_75t_L g1304 ( .A(n_1209), .B(n_1109), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1226), .B(n_1118), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1226), .B(n_1172), .Y(n_1306) );
OAI22xp5_ASAP7_75t_L g1307 ( .A1(n_1224), .A2(n_1212), .B1(n_1184), .B2(n_1154), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1228), .B(n_1114), .Y(n_1308) );
NAND3xp33_ASAP7_75t_L g1309 ( .A(n_1277), .B(n_1200), .C(n_1197), .Y(n_1309) );
AOI22xp33_ASAP7_75t_SL g1310 ( .A1(n_1263), .A2(n_1154), .B1(n_1171), .B2(n_1195), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1228), .B(n_1114), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1282), .B(n_1114), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1282), .B(n_1171), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1285), .B(n_1171), .Y(n_1314) );
INVxp67_ASAP7_75t_L g1315 ( .A(n_1217), .Y(n_1315) );
NOR2x1p5_ASAP7_75t_L g1316 ( .A(n_1236), .B(n_1212), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1216), .Y(n_1317) );
INVx2_ASAP7_75t_L g1318 ( .A(n_1219), .Y(n_1318) );
OR2x2_ASAP7_75t_L g1319 ( .A(n_1220), .B(n_1195), .Y(n_1319) );
NAND2xp5_ASAP7_75t_L g1320 ( .A(n_1279), .B(n_1297), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1269), .B(n_1138), .Y(n_1321) );
NAND2xp5_ASAP7_75t_L g1322 ( .A(n_1229), .B(n_1239), .Y(n_1322) );
OAI21xp33_ASAP7_75t_SL g1323 ( .A1(n_1283), .A2(n_1294), .B(n_1247), .Y(n_1323) );
BUFx2_ASAP7_75t_L g1324 ( .A(n_1247), .Y(n_1324) );
INVx2_ASAP7_75t_SL g1325 ( .A(n_1250), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1271), .B(n_1273), .Y(n_1326) );
OR2x2_ASAP7_75t_L g1327 ( .A(n_1220), .B(n_1256), .Y(n_1327) );
AOI22xp33_ASAP7_75t_L g1328 ( .A1(n_1251), .A2(n_1278), .B1(n_1231), .B2(n_1276), .Y(n_1328) );
OAI21xp5_ASAP7_75t_L g1329 ( .A1(n_1300), .A2(n_1291), .B(n_1232), .Y(n_1329) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_1238), .B(n_1270), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1285), .B(n_1268), .Y(n_1331) );
HB1xp67_ASAP7_75t_L g1332 ( .A(n_1272), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1287), .B(n_1216), .Y(n_1333) );
AOI21xp5_ASAP7_75t_L g1334 ( .A1(n_1290), .A2(n_1218), .B(n_1302), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1264), .Y(n_1335) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1264), .Y(n_1336) );
NAND4xp25_ASAP7_75t_L g1337 ( .A(n_1288), .B(n_1257), .C(n_1281), .D(n_1296), .Y(n_1337) );
INVx1_ASAP7_75t_SL g1338 ( .A(n_1250), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1268), .B(n_1249), .Y(n_1339) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1284), .Y(n_1340) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1227), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1230), .Y(n_1342) );
NAND2x1p5_ASAP7_75t_L g1343 ( .A(n_1236), .B(n_1218), .Y(n_1343) );
OR2x2_ASAP7_75t_L g1344 ( .A(n_1238), .B(n_1255), .Y(n_1344) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1230), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1245), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_1245), .B(n_1294), .Y(n_1347) );
OR2x2_ASAP7_75t_L g1348 ( .A(n_1234), .B(n_1246), .Y(n_1348) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1234), .Y(n_1349) );
HB1xp67_ASAP7_75t_L g1350 ( .A(n_1242), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1252), .B(n_1242), .Y(n_1351) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1248), .B(n_1249), .Y(n_1352) );
HB1xp67_ASAP7_75t_L g1353 ( .A(n_1252), .Y(n_1353) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1235), .Y(n_1354) );
NOR2xp33_ASAP7_75t_R g1355 ( .A(n_1236), .B(n_1293), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1240), .B(n_1254), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1248), .B(n_1241), .Y(n_1357) );
OAI33xp33_ASAP7_75t_L g1358 ( .A1(n_1254), .A2(n_1260), .A3(n_1275), .B1(n_1267), .B2(n_1304), .B3(n_1301), .Y(n_1358) );
OR2x2_ASAP7_75t_L g1359 ( .A(n_1241), .B(n_1255), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1246), .B(n_1289), .Y(n_1360) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1275), .Y(n_1361) );
AND2x2_ASAP7_75t_SL g1362 ( .A(n_1293), .B(n_1292), .Y(n_1362) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1289), .B(n_1292), .Y(n_1363) );
INVx2_ASAP7_75t_SL g1364 ( .A(n_1261), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1280), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1266), .B(n_1240), .Y(n_1366) );
OAI332xp33_ASAP7_75t_L g1367 ( .A1(n_1259), .A2(n_1304), .A3(n_1280), .B1(n_1262), .B2(n_1301), .B3(n_1233), .C1(n_1223), .C2(n_1258), .Y(n_1367) );
INVx2_ASAP7_75t_L g1368 ( .A(n_1266), .Y(n_1368) );
OR2x2_ASAP7_75t_L g1369 ( .A(n_1262), .B(n_1298), .Y(n_1369) );
OR2x2_ASAP7_75t_L g1370 ( .A(n_1327), .B(n_1286), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1363), .B(n_1286), .Y(n_1371) );
NAND4xp25_ASAP7_75t_L g1372 ( .A(n_1328), .B(n_1295), .C(n_1243), .D(n_1225), .Y(n_1372) );
NAND2xp5_ASAP7_75t_L g1373 ( .A(n_1334), .B(n_1221), .Y(n_1373) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1322), .Y(n_1374) );
NOR2x1_ASAP7_75t_L g1375 ( .A(n_1316), .B(n_1221), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1376 ( .A(n_1363), .B(n_1286), .Y(n_1376) );
HB1xp67_ASAP7_75t_L g1377 ( .A(n_1332), .Y(n_1377) );
AND2x4_ASAP7_75t_L g1378 ( .A(n_1360), .B(n_1303), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1317), .Y(n_1379) );
CKINVDCx16_ASAP7_75t_R g1380 ( .A(n_1355), .Y(n_1380) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1317), .Y(n_1381) );
NOR2x1p5_ASAP7_75t_L g1382 ( .A(n_1337), .B(n_1221), .Y(n_1382) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_1331), .B(n_1298), .Y(n_1383) );
INVx2_ASAP7_75t_L g1384 ( .A(n_1368), .Y(n_1384) );
OAI31xp33_ASAP7_75t_L g1385 ( .A1(n_1309), .A2(n_1299), .A3(n_1303), .B(n_1261), .Y(n_1385) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_1331), .B(n_1253), .Y(n_1386) );
INVx2_ASAP7_75t_L g1387 ( .A(n_1368), .Y(n_1387) );
NOR3xp33_ASAP7_75t_SL g1388 ( .A(n_1329), .B(n_1265), .C(n_1237), .Y(n_1388) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1327), .Y(n_1389) );
INVxp67_ASAP7_75t_L g1390 ( .A(n_1324), .Y(n_1390) );
AND2x2_ASAP7_75t_L g1391 ( .A(n_1366), .B(n_1244), .Y(n_1391) );
NAND2xp67_ASAP7_75t_L g1392 ( .A(n_1333), .B(n_1274), .Y(n_1392) );
NOR2xp33_ASAP7_75t_L g1393 ( .A(n_1315), .B(n_1261), .Y(n_1393) );
XOR2x2_ASAP7_75t_L g1394 ( .A(n_1362), .B(n_1274), .Y(n_1394) );
INVx1_ASAP7_75t_SL g1395 ( .A(n_1338), .Y(n_1395) );
INVxp67_ASAP7_75t_L g1396 ( .A(n_1324), .Y(n_1396) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1335), .Y(n_1397) );
NOR3xp33_ASAP7_75t_L g1398 ( .A(n_1367), .B(n_1244), .C(n_1222), .Y(n_1398) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1335), .Y(n_1399) );
INVx2_ASAP7_75t_L g1400 ( .A(n_1348), .Y(n_1400) );
INVx1_ASAP7_75t_SL g1401 ( .A(n_1325), .Y(n_1401) );
INVx2_ASAP7_75t_L g1402 ( .A(n_1348), .Y(n_1402) );
INVx1_ASAP7_75t_SL g1403 ( .A(n_1325), .Y(n_1403) );
OR2x2_ASAP7_75t_L g1404 ( .A(n_1330), .B(n_1244), .Y(n_1404) );
NOR2xp33_ASAP7_75t_R g1405 ( .A(n_1362), .B(n_1222), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1346), .B(n_1222), .Y(n_1406) );
INVx2_ASAP7_75t_L g1407 ( .A(n_1359), .Y(n_1407) );
NAND2xp5_ASAP7_75t_L g1408 ( .A(n_1330), .B(n_1222), .Y(n_1408) );
NAND2xp5_ASAP7_75t_L g1409 ( .A(n_1326), .B(n_1222), .Y(n_1409) );
AOI21xp5_ASAP7_75t_L g1410 ( .A1(n_1307), .A2(n_1323), .B(n_1310), .Y(n_1410) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1336), .Y(n_1411) );
INVxp67_ASAP7_75t_L g1412 ( .A(n_1320), .Y(n_1412) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1336), .Y(n_1413) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_1360), .B(n_1340), .Y(n_1414) );
OR2x2_ASAP7_75t_L g1415 ( .A(n_1369), .B(n_1344), .Y(n_1415) );
NOR2xp33_ASAP7_75t_L g1416 ( .A(n_1347), .B(n_1321), .Y(n_1416) );
INVx2_ASAP7_75t_L g1417 ( .A(n_1384), .Y(n_1417) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1379), .Y(n_1418) );
AND2x2_ASAP7_75t_L g1419 ( .A(n_1371), .B(n_1312), .Y(n_1419) );
HB1xp67_ASAP7_75t_L g1420 ( .A(n_1377), .Y(n_1420) );
INVxp67_ASAP7_75t_L g1421 ( .A(n_1416), .Y(n_1421) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1379), .Y(n_1422) );
INVxp67_ASAP7_75t_L g1423 ( .A(n_1401), .Y(n_1423) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1381), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1381), .Y(n_1425) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1413), .Y(n_1426) );
NAND2xp5_ASAP7_75t_L g1427 ( .A(n_1386), .B(n_1312), .Y(n_1427) );
A2O1A1Ixp33_ASAP7_75t_L g1428 ( .A1(n_1410), .A2(n_1364), .B(n_1353), .C(n_1350), .Y(n_1428) );
NOR2xp33_ASAP7_75t_L g1429 ( .A(n_1380), .B(n_1364), .Y(n_1429) );
AOI21xp5_ASAP7_75t_L g1430 ( .A1(n_1394), .A2(n_1358), .B(n_1343), .Y(n_1430) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1415), .Y(n_1431) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_1389), .B(n_1366), .Y(n_1432) );
INVx1_ASAP7_75t_SL g1433 ( .A(n_1395), .Y(n_1433) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1412), .B(n_1339), .Y(n_1434) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1415), .Y(n_1435) );
NAND2xp5_ASAP7_75t_SL g1436 ( .A(n_1405), .B(n_1343), .Y(n_1436) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_1374), .B(n_1339), .Y(n_1437) );
OAI32xp33_ASAP7_75t_L g1438 ( .A1(n_1373), .A2(n_1343), .A3(n_1319), .B1(n_1369), .B2(n_1344), .Y(n_1438) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1413), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_1371), .B(n_1352), .Y(n_1440) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1376), .B(n_1352), .Y(n_1441) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1414), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1443 ( .A(n_1376), .B(n_1311), .Y(n_1443) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1384), .Y(n_1444) );
OR2x2_ASAP7_75t_L g1445 ( .A(n_1400), .B(n_1356), .Y(n_1445) );
XOR2xp5_ASAP7_75t_L g1446 ( .A(n_1372), .B(n_1351), .Y(n_1446) );
AOI21xp5_ASAP7_75t_L g1447 ( .A1(n_1394), .A2(n_1319), .B(n_1345), .Y(n_1447) );
XNOR2x2_ASAP7_75t_SL g1448 ( .A(n_1405), .B(n_1314), .Y(n_1448) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1397), .Y(n_1449) );
INVxp67_ASAP7_75t_L g1450 ( .A(n_1403), .Y(n_1450) );
AND2x4_ASAP7_75t_L g1451 ( .A(n_1391), .B(n_1305), .Y(n_1451) );
AOI221x1_ASAP7_75t_L g1452 ( .A1(n_1398), .A2(n_1361), .B1(n_1365), .B2(n_1341), .C(n_1354), .Y(n_1452) );
NAND3xp33_ASAP7_75t_L g1453 ( .A(n_1388), .B(n_1361), .C(n_1365), .Y(n_1453) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1399), .Y(n_1454) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1411), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_1400), .B(n_1308), .Y(n_1456) );
INVx2_ASAP7_75t_L g1457 ( .A(n_1387), .Y(n_1457) );
HB1xp67_ASAP7_75t_L g1458 ( .A(n_1402), .Y(n_1458) );
AOI22xp5_ASAP7_75t_L g1459 ( .A1(n_1382), .A2(n_1308), .B1(n_1311), .B2(n_1305), .Y(n_1459) );
OAI22xp5_ASAP7_75t_L g1460 ( .A1(n_1375), .A2(n_1359), .B1(n_1314), .B2(n_1342), .Y(n_1460) );
OAI221xp5_ASAP7_75t_L g1461 ( .A1(n_1385), .A2(n_1393), .B1(n_1370), .B2(n_1390), .C(n_1396), .Y(n_1461) );
XOR2xp5_ASAP7_75t_L g1462 ( .A(n_1378), .B(n_1357), .Y(n_1462) );
OR2x2_ASAP7_75t_L g1463 ( .A(n_1402), .B(n_1357), .Y(n_1463) );
INVxp33_ASAP7_75t_L g1464 ( .A(n_1370), .Y(n_1464) );
NAND2xp5_ASAP7_75t_L g1465 ( .A(n_1407), .B(n_1313), .Y(n_1465) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1383), .Y(n_1466) );
INVx1_ASAP7_75t_SL g1467 ( .A(n_1378), .Y(n_1467) );
INVxp33_ASAP7_75t_SL g1468 ( .A(n_1391), .Y(n_1468) );
OAI211xp5_ASAP7_75t_L g1469 ( .A1(n_1404), .A2(n_1313), .B(n_1306), .C(n_1354), .Y(n_1469) );
OAI21xp33_ASAP7_75t_L g1470 ( .A1(n_1392), .A2(n_1378), .B(n_1407), .Y(n_1470) );
OR2x2_ASAP7_75t_L g1471 ( .A(n_1456), .B(n_1463), .Y(n_1471) );
NAND2x1_ASAP7_75t_L g1472 ( .A(n_1459), .B(n_1448), .Y(n_1472) );
HB1xp67_ASAP7_75t_L g1473 ( .A(n_1420), .Y(n_1473) );
OAI211xp5_ASAP7_75t_SL g1474 ( .A1(n_1461), .A2(n_1428), .B(n_1421), .C(n_1430), .Y(n_1474) );
NAND4xp75_ASAP7_75t_L g1475 ( .A(n_1452), .B(n_1447), .C(n_1429), .D(n_1436), .Y(n_1475) );
AOI221xp5_ASAP7_75t_L g1476 ( .A1(n_1446), .A2(n_1438), .B1(n_1442), .B2(n_1470), .C(n_1453), .Y(n_1476) );
OAI21x1_ASAP7_75t_SL g1477 ( .A1(n_1462), .A2(n_1460), .B(n_1434), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1478 ( .A(n_1435), .B(n_1431), .Y(n_1478) );
AOI21xp33_ASAP7_75t_L g1479 ( .A1(n_1446), .A2(n_1433), .B(n_1438), .Y(n_1479) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1422), .Y(n_1480) );
AOI22xp5_ASAP7_75t_L g1481 ( .A1(n_1468), .A2(n_1466), .B1(n_1450), .B2(n_1423), .Y(n_1481) );
OAI31xp33_ASAP7_75t_L g1482 ( .A1(n_1469), .A2(n_1468), .A3(n_1467), .B(n_1464), .Y(n_1482) );
OAI21xp33_ASAP7_75t_L g1483 ( .A1(n_1464), .A2(n_1427), .B(n_1437), .Y(n_1483) );
AOI21xp5_ASAP7_75t_L g1484 ( .A1(n_1458), .A2(n_1451), .B(n_1444), .Y(n_1484) );
XNOR2xp5_ASAP7_75t_L g1485 ( .A(n_1432), .B(n_1445), .Y(n_1485) );
OAI221xp5_ASAP7_75t_L g1486 ( .A1(n_1472), .A2(n_1449), .B1(n_1455), .B2(n_1454), .C(n_1445), .Y(n_1486) );
AOI21xp5_ASAP7_75t_L g1487 ( .A1(n_1482), .A2(n_1451), .B(n_1444), .Y(n_1487) );
NAND2xp5_ASAP7_75t_L g1488 ( .A(n_1473), .B(n_1443), .Y(n_1488) );
AOI21xp5_ASAP7_75t_L g1489 ( .A1(n_1482), .A2(n_1451), .B(n_1409), .Y(n_1489) );
AOI22xp5_ASAP7_75t_L g1490 ( .A1(n_1474), .A2(n_1443), .B1(n_1419), .B2(n_1441), .Y(n_1490) );
NAND4xp25_ASAP7_75t_L g1491 ( .A(n_1479), .B(n_1404), .C(n_1408), .D(n_1306), .Y(n_1491) );
OAI211xp5_ASAP7_75t_SL g1492 ( .A1(n_1476), .A2(n_1465), .B(n_1418), .C(n_1439), .Y(n_1492) );
BUFx2_ASAP7_75t_L g1493 ( .A(n_1481), .Y(n_1493) );
AOI21xp5_ASAP7_75t_L g1494 ( .A1(n_1477), .A2(n_1417), .B(n_1457), .Y(n_1494) );
AOI21xp5_ASAP7_75t_L g1495 ( .A1(n_1484), .A2(n_1417), .B(n_1457), .Y(n_1495) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1488), .Y(n_1496) );
AOI22xp5_ASAP7_75t_L g1497 ( .A1(n_1493), .A2(n_1475), .B1(n_1483), .B2(n_1478), .Y(n_1497) );
OAI22xp5_ASAP7_75t_L g1498 ( .A1(n_1486), .A2(n_1485), .B1(n_1471), .B2(n_1480), .Y(n_1498) );
OAI211xp5_ASAP7_75t_L g1499 ( .A1(n_1492), .A2(n_1425), .B(n_1422), .C(n_1424), .Y(n_1499) );
INVx2_ASAP7_75t_L g1500 ( .A(n_1490), .Y(n_1500) );
INVx1_ASAP7_75t_L g1501 ( .A(n_1495), .Y(n_1501) );
INVx2_ASAP7_75t_L g1502 ( .A(n_1494), .Y(n_1502) );
XNOR2xp5_ASAP7_75t_L g1503 ( .A(n_1497), .B(n_1491), .Y(n_1503) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1496), .Y(n_1504) );
OAI22xp5_ASAP7_75t_L g1505 ( .A1(n_1497), .A2(n_1487), .B1(n_1489), .B2(n_1463), .Y(n_1505) );
AOI22xp33_ASAP7_75t_L g1506 ( .A1(n_1500), .A2(n_1426), .B1(n_1418), .B2(n_1425), .Y(n_1506) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1501), .Y(n_1507) );
NAND4xp25_ASAP7_75t_L g1508 ( .A(n_1507), .B(n_1498), .C(n_1502), .D(n_1499), .Y(n_1508) );
AOI22xp5_ASAP7_75t_L g1509 ( .A1(n_1503), .A2(n_1419), .B1(n_1441), .B2(n_1440), .Y(n_1509) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1504), .Y(n_1510) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1506), .Y(n_1511) );
XNOR2xp5_ASAP7_75t_L g1512 ( .A(n_1508), .B(n_1505), .Y(n_1512) );
AOI22xp5_ASAP7_75t_L g1513 ( .A1(n_1511), .A2(n_1506), .B1(n_1440), .B2(n_1439), .Y(n_1513) );
INVx2_ASAP7_75t_L g1514 ( .A(n_1510), .Y(n_1514) );
NOR3xp33_ASAP7_75t_L g1515 ( .A(n_1514), .B(n_1509), .C(n_1426), .Y(n_1515) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1512), .Y(n_1516) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1513), .Y(n_1517) );
AOI22xp33_ASAP7_75t_L g1518 ( .A1(n_1516), .A2(n_1424), .B1(n_1387), .B2(n_1406), .Y(n_1518) );
OAI222xp33_ASAP7_75t_L g1519 ( .A1(n_1517), .A2(n_1342), .B1(n_1341), .B2(n_1345), .C1(n_1349), .C2(n_1318), .Y(n_1519) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1515), .Y(n_1520) );
AOI21xp5_ASAP7_75t_L g1521 ( .A1(n_1520), .A2(n_1518), .B(n_1519), .Y(n_1521) );
endmodule