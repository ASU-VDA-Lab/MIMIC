module fake_jpeg_21292_n_298 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_1),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_41),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_45),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_18),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_17),
.B1(n_28),
.B2(n_25),
.Y(n_54)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_59),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_55),
.Y(n_62)
);

AND2x6_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_21),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_31),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_39),
.B1(n_40),
.B2(n_38),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_40),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_74),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_67),
.B(n_71),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_76),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_18),
.B1(n_39),
.B2(n_20),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_73),
.A2(n_84),
.B1(n_94),
.B2(n_97),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_38),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_38),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_75),
.A2(n_77),
.B(n_79),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_43),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_16),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_60),
.B1(n_54),
.B2(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_80),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_18),
.B1(n_24),
.B2(n_20),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_39),
.B1(n_18),
.B2(n_45),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_15),
.B1(n_43),
.B2(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_82),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_45),
.B1(n_43),
.B2(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_19),
.B1(n_20),
.B2(n_24),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_46),
.A2(n_15),
.B1(n_34),
.B2(n_23),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_88),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_22),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_86),
.Y(n_134)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_22),
.B1(n_19),
.B2(n_32),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_22),
.B1(n_15),
.B2(n_23),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_92),
.B(n_62),
.Y(n_104)
);

OAI32xp33_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_92),
.A3(n_21),
.B1(n_31),
.B2(n_16),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_33),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_95),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_25),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_46),
.A2(n_15),
.B1(n_25),
.B2(n_32),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_51),
.A2(n_14),
.B1(n_17),
.B2(n_32),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_26),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_26),
.C(n_16),
.Y(n_113)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_99),
.A2(n_33),
.B1(n_36),
.B2(n_28),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_56),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_101),
.Y(n_136)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_51),
.A2(n_29),
.B1(n_14),
.B2(n_28),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_103),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_51),
.A2(n_29),
.B1(n_26),
.B2(n_16),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_104),
.A2(n_122),
.B(n_125),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_21),
.C(n_29),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_113),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_120),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_65),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_127),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_63),
.A2(n_21),
.B(n_31),
.C(n_14),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_77),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_26),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_83),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_87),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_67),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_63),
.A2(n_9),
.B(n_13),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

AND2x4_ASAP7_75t_SL g138 ( 
.A(n_129),
.B(n_71),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_138),
.A2(n_157),
.B(n_130),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_90),
.C(n_77),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_139),
.B(n_158),
.C(n_159),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_135),
.B(n_76),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_145),
.Y(n_167)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_110),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_149),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_137),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_117),
.A2(n_102),
.B1(n_70),
.B2(n_103),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_160),
.B1(n_118),
.B2(n_125),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_75),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_151),
.B(n_162),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_136),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_165),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_66),
.Y(n_155)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_66),
.B1(n_74),
.B2(n_75),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_156),
.A2(n_112),
.B1(n_129),
.B2(n_113),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_104),
.A2(n_74),
.B(n_72),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_98),
.C(n_82),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_98),
.C(n_80),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_116),
.A2(n_79),
.B1(n_89),
.B2(n_64),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_85),
.C(n_96),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_120),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_61),
.Y(n_162)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_137),
.A2(n_99),
.B1(n_101),
.B2(n_95),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_112),
.B(n_93),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_139),
.B(n_106),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_178),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_169),
.A2(n_190),
.B1(n_119),
.B2(n_110),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_173),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_154),
.A2(n_109),
.B(n_118),
.C(n_105),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_140),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_176),
.B(n_177),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_SL g196 ( 
.A1(n_180),
.A2(n_188),
.B(n_156),
.C(n_144),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_123),
.B1(n_130),
.B2(n_125),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_169),
.B1(n_166),
.B2(n_183),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_184),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_107),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_144),
.B(n_147),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_105),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_187),
.B(n_191),
.Y(n_212)
);

AND2x6_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_126),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_123),
.B1(n_160),
.B2(n_152),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_141),
.B(n_107),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_159),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_134),
.Y(n_193)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_182),
.A2(n_155),
.A3(n_150),
.B1(n_157),
.B2(n_142),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_204),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_196),
.A2(n_173),
.B1(n_168),
.B2(n_167),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_203),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_142),
.C(n_158),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_213),
.C(n_178),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_207),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_161),
.B1(n_153),
.B2(n_149),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_215),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_119),
.B1(n_143),
.B2(n_163),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_214),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_132),
.C(n_108),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_163),
.B1(n_132),
.B2(n_17),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_13),
.B1(n_11),
.B2(n_9),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_176),
.A2(n_13),
.B(n_11),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_175),
.Y(n_225)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_224),
.C(n_229),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_192),
.C(n_183),
.Y(n_224)
);

NOR3xp33_ASAP7_75t_SL g249 ( 
.A(n_225),
.B(n_201),
.C(n_211),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_175),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_232),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_180),
.C(n_174),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_174),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_214),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_167),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_179),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_205),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_234),
.B(n_235),
.Y(n_243)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_191),
.C(n_172),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_208),
.C(n_196),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_227),
.A2(n_217),
.B1(n_215),
.B2(n_206),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_239),
.A2(n_241),
.B1(n_250),
.B2(n_255),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_231),
.A2(n_204),
.B1(n_202),
.B2(n_196),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_247),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_238),
.B(n_201),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_244),
.B(n_249),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_196),
.C(n_210),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_248),
.C(n_254),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_172),
.C(n_194),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_231),
.A2(n_211),
.B1(n_181),
.B2(n_179),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_181),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_253),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_229),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_179),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_230),
.B(n_9),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_220),
.A2(n_237),
.B1(n_221),
.B2(n_223),
.Y(n_255)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_237),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_259),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_243),
.B(n_236),
.Y(n_259)
);

XOR2x1_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_232),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_262),
.A2(n_242),
.B1(n_253),
.B2(n_251),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_232),
.B1(n_33),
.B2(n_4),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_264),
.B(n_267),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_0),
.B(n_3),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_266),
.A2(n_268),
.B(n_3),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_267)
);

OA22x2_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_33),
.B1(n_4),
.B2(n_5),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_240),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_271),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_240),
.Y(n_271)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_256),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_263),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_275),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_257),
.A2(n_254),
.B(n_33),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_269),
.B(n_267),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_276),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_279),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_265),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_268),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_263),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_287),
.Y(n_292)
);

NOR3xp33_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_262),
.C(n_268),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_288),
.Y(n_291)
);

AOI21x1_ASAP7_75t_L g289 ( 
.A1(n_281),
.A2(n_274),
.B(n_261),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_279),
.B(n_284),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_290),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_292),
.B(n_261),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_SL g295 ( 
.A1(n_294),
.A2(n_291),
.B(n_7),
.C(n_8),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_6),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_293),
.B(n_7),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_6),
.Y(n_298)
);


endmodule