module fake_aes_5652_n_18 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_18);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
NOR2xp33_ASAP7_75t_L g10 ( .A(n_2), .B(n_0), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_4), .B(n_3), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_8), .Y(n_12) );
OAI21x1_ASAP7_75t_L g13 ( .A1(n_9), .A2(n_5), .B(n_0), .Y(n_13) );
BUFx3_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_14), .Y(n_15) );
NAND3xp33_ASAP7_75t_L g16 ( .A(n_15), .B(n_14), .C(n_10), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
OAI222xp33_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_1), .B1(n_11), .B2(n_13), .C1(n_8), .C2(n_9), .Y(n_18) );
endmodule