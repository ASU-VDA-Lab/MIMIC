module fake_netlist_5_1366_n_2035 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_451, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_483, n_155, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_507, n_119, n_497, n_275, n_252, n_26, n_295, n_133, n_330, n_506, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_492, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_470, n_325, n_449, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_457, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_145, n_48, n_50, n_337, n_430, n_313, n_88, n_479, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_309, n_30, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_441, n_450, n_312, n_476, n_429, n_345, n_210, n_494, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_480, n_237, n_425, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_409, n_500, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_391, n_434, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_52, n_278, n_110, n_2035);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_451;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_483;
input n_155;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_507;
input n_119;
input n_497;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_506;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_480;
input n_237;
input n_425;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_409;
input n_500;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_391;
input n_434;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_2035;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_877;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_1230;
wire n_668;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_920;
wire n_1289;
wire n_1517;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_1948;
wire n_1984;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_1218;
wire n_1931;
wire n_1070;
wire n_777;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1587;
wire n_1473;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_889;
wire n_973;
wire n_1700;
wire n_571;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_1819;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_832;
wire n_857;
wire n_1319;
wire n_561;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_677;
wire n_1333;
wire n_1121;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_514;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_1593;
wire n_1033;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_1609;
wire n_1989;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_662;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_1870;
wire n_512;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_1823;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_1805;
wire n_1816;
wire n_948;
wire n_1217;
wire n_628;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_1552;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_824;
wire n_1645;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_815;
wire n_1795;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1958;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_1519;
wire n_950;
wire n_1553;
wire n_1811;
wire n_1346;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_912;
wire n_968;
wire n_619;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_1432;
wire n_1357;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_1179;
wire n_621;
wire n_753;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_1560;
wire n_1605;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_1584;
wire n_665;
wire n_1835;
wire n_1726;
wire n_1440;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2003;
wire n_1457;
wire n_766;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_676;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_1999;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_1235;
wire n_980;
wire n_703;
wire n_698;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_1589;
wire n_517;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_542;
wire n_1546;
wire n_595;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_1937;
wire n_585;
wire n_1739;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_575;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2027;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;

INVx1_ASAP7_75t_L g508 ( 
.A(n_199),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_143),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_485),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_30),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_303),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_404),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_487),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_389),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_391),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_157),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_85),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_153),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_143),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_0),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_100),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_8),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_86),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_115),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_312),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_430),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_385),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_282),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_379),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_495),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_277),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_229),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_368),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_344),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_483),
.Y(n_536)
);

CKINVDCx14_ASAP7_75t_R g537 ( 
.A(n_347),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_109),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_361),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_428),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_4),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_261),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_90),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_65),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_463),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_294),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_3),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_17),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_279),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_462),
.Y(n_550)
);

BUFx10_ASAP7_75t_L g551 ( 
.A(n_99),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_26),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_238),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_213),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_194),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_30),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_240),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_263),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_441),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_269),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_307),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_459),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_465),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_166),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_319),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_186),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_79),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_301),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_187),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_346),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_349),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_222),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_413),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_100),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_275),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_371),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_109),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_357),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_305),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_309),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_504),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_494),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_442),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_115),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_406),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_110),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_252),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_322),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_19),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_401),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_200),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_276),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_245),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_278),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_153),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_215),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_458),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_266),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_183),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_281),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_270),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_370),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_130),
.Y(n_603)
);

CKINVDCx16_ASAP7_75t_R g604 ( 
.A(n_295),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_167),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_179),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_163),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_284),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_268),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_449),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_154),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_236),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_126),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_32),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_44),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_296),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_293),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_41),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_228),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_95),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_342),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_488),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_66),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_314),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_11),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_334),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_129),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_174),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_259),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_480),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_367),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_60),
.Y(n_632)
);

BUFx10_ASAP7_75t_L g633 ( 
.A(n_89),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_185),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_90),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_398),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_383),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_395),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_331),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_377),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_297),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_338),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_134),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_491),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_426),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_99),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_366),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_411),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_106),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_97),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_32),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_147),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_335),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_429),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_114),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_95),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_77),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_140),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_93),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_4),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_424),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_468),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_456),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_384),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_218),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_181),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_298),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_315),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_300),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_486),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_190),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_464),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_188),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_336),
.Y(n_674)
);

BUFx10_ASAP7_75t_L g675 ( 
.A(n_501),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_59),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_402),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_139),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_231),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_244),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_172),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_118),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_360),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_141),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_37),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_448),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_412),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_400),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_201),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_503),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_85),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_341),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_19),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_203),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_493),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_500),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_217),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_51),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_248),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_455),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_481),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_55),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_423),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_570),
.Y(n_704)
);

INVxp67_ASAP7_75t_SL g705 ( 
.A(n_529),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_606),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_523),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_606),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_549),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_545),
.Y(n_710)
);

INVxp33_ASAP7_75t_SL g711 ( 
.A(n_544),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_646),
.B(n_0),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_510),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_512),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_618),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_618),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_646),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_646),
.Y(n_718)
);

INVxp67_ASAP7_75t_SL g719 ( 
.A(n_534),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_646),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_508),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_517),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_562),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_525),
.Y(n_724)
);

CKINVDCx14_ASAP7_75t_R g725 ( 
.A(n_537),
.Y(n_725)
);

INVxp67_ASAP7_75t_SL g726 ( 
.A(n_570),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_545),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_547),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_567),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_577),
.Y(n_730)
);

INVxp67_ASAP7_75t_SL g731 ( 
.A(n_594),
.Y(n_731)
);

INVxp67_ASAP7_75t_SL g732 ( 
.A(n_594),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_513),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_509),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_557),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_613),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_688),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_620),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_627),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_634),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_649),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_511),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_514),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_650),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_651),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_652),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_657),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_590),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_659),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_516),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_578),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_660),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_682),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_527),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_549),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_688),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_518),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_566),
.B(n_1),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_684),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_685),
.Y(n_760)
);

INVxp67_ASAP7_75t_SL g761 ( 
.A(n_622),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_590),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_689),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_528),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_532),
.Y(n_765)
);

CKINVDCx14_ASAP7_75t_R g766 ( 
.A(n_537),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_691),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_702),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_549),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_535),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_526),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_530),
.Y(n_772)
);

CKINVDCx16_ASAP7_75t_R g773 ( 
.A(n_531),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_539),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_536),
.Y(n_775)
);

CKINVDCx20_ASAP7_75t_R g776 ( 
.A(n_596),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_509),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_569),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_683),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_546),
.Y(n_780)
);

INVxp33_ASAP7_75t_SL g781 ( 
.A(n_519),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_553),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_540),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_550),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_551),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_554),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_558),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_560),
.Y(n_788)
);

CKINVDCx16_ASAP7_75t_R g789 ( 
.A(n_604),
.Y(n_789)
);

INVxp67_ASAP7_75t_SL g790 ( 
.A(n_561),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_565),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_785),
.Y(n_792)
);

AND2x2_ASAP7_75t_R g793 ( 
.A(n_710),
.B(n_596),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_704),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_713),
.B(n_533),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_726),
.B(n_569),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_717),
.Y(n_797)
);

INVx5_ASAP7_75t_L g798 ( 
.A(n_709),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_709),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_711),
.A2(n_608),
.B1(n_598),
.B2(n_687),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_718),
.Y(n_801)
);

OA21x2_ASAP7_75t_L g802 ( 
.A1(n_771),
.A2(n_580),
.B(n_515),
.Y(n_802)
);

BUFx12f_ASAP7_75t_L g803 ( 
.A(n_714),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_720),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_704),
.B(n_614),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_772),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_733),
.B(n_542),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_734),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_709),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_709),
.Y(n_810)
);

OA21x2_ASAP7_75t_L g811 ( 
.A1(n_774),
.A2(n_782),
.B(n_780),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_731),
.B(n_607),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_755),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_743),
.B(n_515),
.Y(n_814)
);

INVx4_ASAP7_75t_L g815 ( 
.A(n_755),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_750),
.B(n_580),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_755),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_754),
.B(n_624),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_732),
.B(n_607),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_786),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_755),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_781),
.B(n_697),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_764),
.B(n_624),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_765),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_769),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_756),
.B(n_623),
.Y(n_826)
);

OA21x2_ASAP7_75t_L g827 ( 
.A1(n_787),
.A2(n_636),
.B(n_626),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_770),
.B(n_626),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_775),
.B(n_783),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_769),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_784),
.B(n_636),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_788),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_769),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_725),
.B(n_690),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_769),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_790),
.B(n_737),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_737),
.B(n_791),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_734),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_777),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_777),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_778),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_778),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_725),
.B(n_690),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_721),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_722),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_724),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_728),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_839),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_839),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_836),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_847),
.Y(n_851)
);

CKINVDCx6p67_ASAP7_75t_R g852 ( 
.A(n_803),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_847),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_839),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_817),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_836),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_796),
.B(n_705),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_839),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_847),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_805),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_814),
.B(n_766),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_839),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_840),
.Y(n_863)
);

AND3x2_ASAP7_75t_L g864 ( 
.A(n_822),
.B(n_712),
.C(n_697),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_840),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_840),
.Y(n_866)
);

OAI21xp33_ASAP7_75t_SL g867 ( 
.A1(n_796),
.A2(n_719),
.B(n_758),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_840),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_794),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_847),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_847),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_797),
.Y(n_872)
);

BUFx10_ASAP7_75t_L g873 ( 
.A(n_829),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_840),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_816),
.B(n_761),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_818),
.B(n_742),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_805),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_842),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_SL g879 ( 
.A1(n_800),
.A2(n_727),
.B1(n_735),
.B2(n_710),
.Y(n_879)
);

CKINVDCx6p67_ASAP7_75t_R g880 ( 
.A(n_803),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_842),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_823),
.B(n_773),
.Y(n_882)
);

INVx5_ASAP7_75t_L g883 ( 
.A(n_817),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_842),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_842),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_794),
.B(n_692),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_828),
.B(n_831),
.Y(n_887)
);

INVxp33_ASAP7_75t_SL g888 ( 
.A(n_824),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_842),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_812),
.B(n_706),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_838),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_838),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_841),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_834),
.B(n_843),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_812),
.B(n_708),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_801),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_819),
.A2(n_608),
.B1(n_598),
.B2(n_541),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_837),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_804),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_841),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_804),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_799),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_799),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_795),
.B(n_807),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_826),
.B(n_715),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_824),
.B(n_789),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_809),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_837),
.Y(n_908)
);

INVxp67_ASAP7_75t_SL g909 ( 
.A(n_825),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_811),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_810),
.Y(n_911)
);

BUFx6f_ASAP7_75t_SL g912 ( 
.A(n_837),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_826),
.B(n_757),
.Y(n_913)
);

AOI21x1_ASAP7_75t_L g914 ( 
.A1(n_802),
.A2(n_692),
.B(n_579),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_810),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_792),
.B(n_707),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_813),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_813),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_811),
.Y(n_919)
);

INVxp33_ASAP7_75t_SL g920 ( 
.A(n_792),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_821),
.Y(n_921)
);

INVx5_ASAP7_75t_L g922 ( 
.A(n_817),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_806),
.B(n_675),
.Y(n_923)
);

INVxp33_ASAP7_75t_L g924 ( 
.A(n_844),
.Y(n_924)
);

AOI21x1_ASAP7_75t_L g925 ( 
.A1(n_802),
.A2(n_581),
.B(n_576),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_899),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_860),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_899),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_901),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_904),
.B(n_723),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_872),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_898),
.B(n_845),
.Y(n_932)
);

XOR2xp5_ASAP7_75t_L g933 ( 
.A(n_888),
.B(n_751),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_872),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_910),
.B(n_802),
.Y(n_935)
);

INVxp67_ASAP7_75t_SL g936 ( 
.A(n_910),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_896),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_896),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_852),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_SL g940 ( 
.A(n_873),
.B(n_675),
.Y(n_940)
);

INVxp33_ASAP7_75t_L g941 ( 
.A(n_916),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_850),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_850),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_898),
.Y(n_944)
);

XNOR2xp5_ASAP7_75t_L g945 ( 
.A(n_879),
.B(n_779),
.Y(n_945)
);

NOR2xp67_ASAP7_75t_L g946 ( 
.A(n_856),
.B(n_821),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_856),
.Y(n_947)
);

XOR2xp5_ASAP7_75t_L g948 ( 
.A(n_888),
.B(n_727),
.Y(n_948)
);

OR2x6_ASAP7_75t_L g949 ( 
.A(n_879),
.B(n_716),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_908),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_919),
.A2(n_827),
.B(n_712),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_908),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_891),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_887),
.B(n_735),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_891),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_892),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_893),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_893),
.Y(n_958)
);

XOR2x2_ASAP7_75t_L g959 ( 
.A(n_897),
.B(n_793),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_900),
.Y(n_960)
);

NOR2xp67_ASAP7_75t_L g961 ( 
.A(n_919),
.B(n_833),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_902),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_902),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_903),
.Y(n_964)
);

INVxp33_ASAP7_75t_L g965 ( 
.A(n_897),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_852),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_907),
.Y(n_967)
);

INVx4_ASAP7_75t_L g968 ( 
.A(n_912),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_873),
.Y(n_969)
);

XNOR2xp5_ASAP7_75t_L g970 ( 
.A(n_906),
.B(n_748),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_860),
.B(n_748),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_877),
.B(n_762),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_911),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_894),
.B(n_820),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_876),
.B(n_762),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_911),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_915),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_915),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_875),
.B(n_776),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_877),
.Y(n_980)
);

OR2x2_ASAP7_75t_L g981 ( 
.A(n_913),
.B(n_693),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_917),
.Y(n_982)
);

INVxp33_ASAP7_75t_L g983 ( 
.A(n_890),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_917),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_918),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_873),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_918),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_880),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_882),
.B(n_776),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_924),
.B(n_832),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_873),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_857),
.B(n_895),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_SL g993 ( 
.A(n_920),
.B(n_615),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_921),
.Y(n_994)
);

XOR2xp5_ASAP7_75t_L g995 ( 
.A(n_920),
.B(n_568),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_921),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_895),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_905),
.Y(n_998)
);

AND2x6_ASAP7_75t_L g999 ( 
.A(n_857),
.B(n_549),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_886),
.B(n_869),
.Y(n_1000)
);

XOR2xp5_ASAP7_75t_L g1001 ( 
.A(n_861),
.B(n_571),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_909),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_886),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_848),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_886),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_886),
.B(n_846),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_855),
.Y(n_1007)
);

INVxp67_ASAP7_75t_L g1008 ( 
.A(n_923),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_851),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_851),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_848),
.Y(n_1011)
);

NAND2xp33_ASAP7_75t_R g1012 ( 
.A(n_864),
.B(n_827),
.Y(n_1012)
);

XOR2xp5_ASAP7_75t_L g1013 ( 
.A(n_880),
.B(n_572),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_849),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_853),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_853),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_859),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_859),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_870),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_867),
.B(n_573),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_870),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_871),
.B(n_811),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_871),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_849),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_912),
.B(n_520),
.Y(n_1025)
);

OR2x2_ASAP7_75t_SL g1026 ( 
.A(n_912),
.B(n_623),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_854),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_854),
.Y(n_1028)
);

INVxp33_ASAP7_75t_SL g1029 ( 
.A(n_858),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_858),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_862),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_863),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_865),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_865),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_866),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_866),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_868),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_868),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_874),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_855),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_874),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_974),
.B(n_878),
.Y(n_1042)
);

OAI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_965),
.A2(n_587),
.B1(n_592),
.B2(n_582),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_974),
.A2(n_600),
.B1(n_602),
.B2(n_597),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_992),
.B(n_575),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_941),
.B(n_930),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_955),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_1000),
.B(n_944),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_954),
.B(n_521),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_960),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_979),
.B(n_975),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_SL g1052 ( 
.A1(n_993),
.A2(n_633),
.B1(n_551),
.B2(n_563),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_944),
.Y(n_1053)
);

NAND2xp33_ASAP7_75t_L g1054 ( 
.A(n_1005),
.B(n_878),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_936),
.B(n_881),
.Y(n_1055)
);

BUFx12f_ASAP7_75t_L g1056 ( 
.A(n_968),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_990),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_1003),
.A2(n_884),
.B1(n_885),
.B2(n_881),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_1006),
.A2(n_885),
.B1(n_889),
.B2(n_884),
.Y(n_1059)
);

O2A1O1Ixp5_ASAP7_75t_L g1060 ( 
.A1(n_1020),
.A2(n_914),
.B(n_925),
.C(n_889),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_926),
.B(n_855),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_971),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_989),
.B(n_522),
.Y(n_1063)
);

NOR3xp33_ASAP7_75t_SL g1064 ( 
.A(n_969),
.B(n_538),
.C(n_524),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_928),
.Y(n_1065)
);

NOR2xp67_ASAP7_75t_L g1066 ( 
.A(n_942),
.B(n_925),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_929),
.B(n_609),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_944),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_935),
.A2(n_961),
.B(n_1022),
.Y(n_1069)
);

AND2x6_ASAP7_75t_SL g1070 ( 
.A(n_949),
.B(n_729),
.Y(n_1070)
);

NAND2x1_ASAP7_75t_L g1071 ( 
.A(n_1005),
.B(n_1007),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_1000),
.B(n_583),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_972),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_927),
.B(n_543),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_1005),
.Y(n_1075)
);

OAI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_940),
.A2(n_617),
.B1(n_621),
.B2(n_616),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1009),
.Y(n_1077)
);

AND2x4_ASAP7_75t_SL g1078 ( 
.A(n_968),
.B(n_633),
.Y(n_1078)
);

NAND2x1_ASAP7_75t_L g1079 ( 
.A(n_1007),
.B(n_833),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_931),
.B(n_637),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1010),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_1040),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_980),
.B(n_932),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_934),
.B(n_937),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_938),
.B(n_639),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_932),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_983),
.B(n_548),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_953),
.Y(n_1088)
);

OR2x6_ASAP7_75t_L g1089 ( 
.A(n_949),
.B(n_625),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_956),
.Y(n_1090)
);

BUFx8_ASAP7_75t_L g1091 ( 
.A(n_981),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_943),
.B(n_644),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1015),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_1040),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1016),
.Y(n_1095)
);

CKINVDCx11_ASAP7_75t_R g1096 ( 
.A(n_939),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_993),
.B(n_585),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_997),
.B(n_730),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1017),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1001),
.B(n_552),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_947),
.B(n_588),
.Y(n_1101)
);

NOR2xp67_ASAP7_75t_L g1102 ( 
.A(n_950),
.B(n_914),
.Y(n_1102)
);

NOR2x1p5_ASAP7_75t_L g1103 ( 
.A(n_986),
.B(n_555),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1002),
.B(n_645),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_995),
.B(n_991),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_951),
.A2(n_653),
.B(n_647),
.Y(n_1106)
);

NAND3xp33_ASAP7_75t_SL g1107 ( 
.A(n_1035),
.B(n_564),
.C(n_556),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_998),
.B(n_661),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_952),
.B(n_593),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1029),
.B(n_663),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_935),
.B(n_672),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_999),
.B(n_1018),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1019),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_1036),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_1038),
.B(n_736),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1021),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_999),
.B(n_677),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_999),
.B(n_808),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_999),
.B(n_808),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1023),
.B(n_961),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_957),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_958),
.B(n_601),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_962),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_949),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1025),
.B(n_738),
.Y(n_1125)
);

BUFx12f_ASAP7_75t_L g1126 ( 
.A(n_1026),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_963),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_1004),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_933),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_951),
.B(n_612),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_946),
.B(n_619),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1008),
.B(n_629),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_964),
.A2(n_563),
.B1(n_610),
.B2(n_559),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_946),
.B(n_1024),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1027),
.B(n_630),
.Y(n_1135)
);

INVxp33_ASAP7_75t_SL g1136 ( 
.A(n_948),
.Y(n_1136)
);

AO22x1_ASAP7_75t_L g1137 ( 
.A1(n_1008),
.A2(n_584),
.B1(n_586),
.B2(n_574),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_970),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1030),
.B(n_631),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_967),
.Y(n_1140)
);

NAND2x1p5_ASAP7_75t_L g1141 ( 
.A(n_1041),
.B(n_883),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_945),
.B(n_1013),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1039),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_1031),
.B(n_589),
.Y(n_1144)
);

NOR2xp67_ASAP7_75t_SL g1145 ( 
.A(n_1032),
.B(n_559),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1033),
.B(n_638),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1034),
.B(n_640),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_973),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_976),
.B(n_641),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_977),
.B(n_642),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_1037),
.B(n_591),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_978),
.B(n_648),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_982),
.B(n_654),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_984),
.B(n_985),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_987),
.B(n_994),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_996),
.B(n_662),
.Y(n_1156)
);

AND2x6_ASAP7_75t_SL g1157 ( 
.A(n_959),
.B(n_739),
.Y(n_1157)
);

NOR2x2_ASAP7_75t_L g1158 ( 
.A(n_1011),
.B(n_595),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1014),
.B(n_664),
.Y(n_1159)
);

NAND2x1p5_ASAP7_75t_L g1160 ( 
.A(n_1028),
.B(n_883),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1012),
.B(n_665),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_966),
.B(n_667),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_988),
.A2(n_669),
.B1(n_670),
.B2(n_668),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_974),
.B(n_674),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_974),
.B(n_679),
.Y(n_1165)
);

OR2x6_ASAP7_75t_L g1166 ( 
.A(n_968),
.B(n_740),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_981),
.B(n_741),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_974),
.B(n_680),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_955),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_941),
.B(n_599),
.Y(n_1170)
);

NOR2x2_ASAP7_75t_L g1171 ( 
.A(n_949),
.B(n_603),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_974),
.B(n_686),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_974),
.B(n_695),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_941),
.B(n_605),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_974),
.A2(n_699),
.B1(n_700),
.B2(n_696),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_974),
.B(n_701),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_974),
.B(n_703),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1035),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_941),
.B(n_611),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_926),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_974),
.B(n_825),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_974),
.B(n_835),
.Y(n_1182)
);

INVx5_ASAP7_75t_L g1183 ( 
.A(n_968),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_955),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_971),
.Y(n_1185)
);

OAI22x1_ASAP7_75t_SL g1186 ( 
.A1(n_939),
.A2(n_632),
.B1(n_635),
.B2(n_628),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_974),
.B(n_835),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_992),
.B(n_559),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_992),
.B(n_563),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1005),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_992),
.B(n_744),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_974),
.B(n_835),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_R g1193 ( 
.A(n_969),
.B(n_643),
.Y(n_1193)
);

OR2x2_ASAP7_75t_L g1194 ( 
.A(n_981),
.B(n_745),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_974),
.B(n_815),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_981),
.B(n_746),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_974),
.B(n_815),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_974),
.B(n_815),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_941),
.B(n_655),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_992),
.B(n_563),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_926),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_941),
.B(n_656),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_992),
.A2(n_610),
.B1(n_749),
.B2(n_747),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_992),
.B(n_752),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_974),
.B(n_610),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_941),
.B(n_658),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_974),
.A2(n_610),
.B1(n_671),
.B2(n_666),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_981),
.B(n_753),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_974),
.B(n_883),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_974),
.B(n_883),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_926),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_992),
.A2(n_760),
.B1(n_763),
.B2(n_759),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_992),
.B(n_817),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_974),
.B(n_883),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_941),
.B(n_673),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_926),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_951),
.A2(n_922),
.B(n_883),
.Y(n_1217)
);

AND2x6_ASAP7_75t_SL g1218 ( 
.A(n_989),
.B(n_767),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1086),
.B(n_768),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1065),
.Y(n_1220)
);

INVx5_ASAP7_75t_L g1221 ( 
.A(n_1056),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1051),
.B(n_676),
.Y(n_1222)
);

NAND2x1p5_ASAP7_75t_L g1223 ( 
.A(n_1053),
.B(n_922),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1088),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1057),
.B(n_678),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1164),
.B(n_681),
.Y(n_1226)
);

OAI221xp5_ASAP7_75t_L g1227 ( 
.A1(n_1049),
.A2(n_698),
.B1(n_694),
.B2(n_3),
.C(n_1),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1090),
.Y(n_1228)
);

NOR3xp33_ASAP7_75t_SL g1229 ( 
.A(n_1107),
.B(n_2),
.C(n_5),
.Y(n_1229)
);

NAND3xp33_ASAP7_75t_SL g1230 ( 
.A(n_1063),
.B(n_2),
.C(n_5),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1165),
.B(n_6),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1046),
.B(n_798),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1086),
.B(n_211),
.Y(n_1233)
);

AND2x6_ASAP7_75t_SL g1234 ( 
.A(n_1142),
.B(n_6),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1168),
.B(n_7),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1125),
.B(n_1191),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_1115),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1172),
.B(n_7),
.Y(n_1238)
);

INVxp67_ASAP7_75t_L g1239 ( 
.A(n_1115),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1180),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1173),
.B(n_8),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1094),
.Y(n_1242)
);

NOR2x1_ASAP7_75t_L g1243 ( 
.A(n_1053),
.B(n_817),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1114),
.Y(n_1244)
);

OR2x6_ASAP7_75t_L g1245 ( 
.A(n_1178),
.B(n_830),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1140),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1201),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1106),
.A2(n_830),
.B(n_922),
.C(n_11),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1176),
.B(n_9),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1183),
.B(n_212),
.Y(n_1250)
);

BUFx4f_ASAP7_75t_L g1251 ( 
.A(n_1126),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1211),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1170),
.B(n_9),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1148),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1075),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1047),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1096),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1050),
.Y(n_1258)
);

INVxp67_ASAP7_75t_SL g1259 ( 
.A(n_1075),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1204),
.B(n_1174),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1177),
.B(n_10),
.Y(n_1261)
);

INVx3_ASAP7_75t_L g1262 ( 
.A(n_1190),
.Y(n_1262)
);

AND3x1_ASAP7_75t_L g1263 ( 
.A(n_1100),
.B(n_10),
.C(n_12),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1179),
.B(n_12),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1190),
.Y(n_1265)
);

BUFx4f_ASAP7_75t_L g1266 ( 
.A(n_1166),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1199),
.B(n_13),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1183),
.B(n_214),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1062),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1042),
.B(n_13),
.Y(n_1270)
);

INVx5_ASAP7_75t_L g1271 ( 
.A(n_1166),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1044),
.A2(n_1043),
.B1(n_1207),
.B2(n_1216),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1202),
.B(n_1206),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1084),
.B(n_14),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1167),
.B(n_14),
.Y(n_1275)
);

AOI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1111),
.A2(n_1069),
.B(n_1066),
.Y(n_1276)
);

NOR3xp33_ASAP7_75t_SL g1277 ( 
.A(n_1163),
.B(n_15),
.C(n_16),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1077),
.Y(n_1278)
);

NOR3xp33_ASAP7_75t_SL g1279 ( 
.A(n_1076),
.B(n_15),
.C(n_16),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1073),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1136),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1215),
.B(n_1185),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1183),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_R g1284 ( 
.A(n_1138),
.B(n_216),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1194),
.B(n_17),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1195),
.B(n_1197),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1129),
.B(n_18),
.Y(n_1287)
);

INVx3_ASAP7_75t_SL g1288 ( 
.A(n_1158),
.Y(n_1288)
);

NAND2xp33_ASAP7_75t_SL g1289 ( 
.A(n_1064),
.B(n_830),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1198),
.B(n_18),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1169),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1091),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1082),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1184),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1091),
.Y(n_1295)
);

CKINVDCx11_ASAP7_75t_R g1296 ( 
.A(n_1070),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1068),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1128),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1081),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1093),
.Y(n_1300)
);

INVx3_ASAP7_75t_L g1301 ( 
.A(n_1082),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1048),
.A2(n_830),
.B1(n_922),
.B2(n_798),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1044),
.A2(n_830),
.B1(n_922),
.B2(n_798),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1095),
.B(n_20),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1161),
.B(n_798),
.Y(n_1305)
);

INVxp67_ASAP7_75t_L g1306 ( 
.A(n_1196),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1099),
.B(n_20),
.Y(n_1307)
);

NOR3xp33_ASAP7_75t_SL g1308 ( 
.A(n_1072),
.B(n_21),
.C(n_22),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1208),
.B(n_21),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1083),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1113),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1166),
.B(n_1098),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_1074),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1116),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1154),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_R g1316 ( 
.A(n_1105),
.B(n_219),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1128),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1087),
.B(n_22),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1162),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1193),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1155),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1055),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1207),
.B(n_1205),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1128),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1143),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1124),
.B(n_220),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1181),
.B(n_23),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1121),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1182),
.B(n_1187),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1089),
.B(n_1052),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1089),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1103),
.B(n_221),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1045),
.A2(n_224),
.B1(n_225),
.B2(n_223),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1218),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1143),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1123),
.Y(n_1336)
);

BUFx4f_ASAP7_75t_L g1337 ( 
.A(n_1143),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1157),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1127),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1078),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1061),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1171),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1067),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1192),
.B(n_23),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1108),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1110),
.B(n_24),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1079),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1175),
.B(n_25),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1104),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1212),
.B(n_25),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1132),
.B(n_1213),
.Y(n_1351)
);

AND2x6_ASAP7_75t_L g1352 ( 
.A(n_1209),
.B(n_226),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1080),
.B(n_26),
.Y(n_1353)
);

INVx8_ASAP7_75t_L g1354 ( 
.A(n_1109),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1071),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1144),
.B(n_27),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1134),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1085),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1137),
.B(n_27),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1160),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1092),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1122),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1130),
.A2(n_31),
.B1(n_28),
.B2(n_29),
.Y(n_1363)
);

CKINVDCx11_ASAP7_75t_R g1364 ( 
.A(n_1186),
.Y(n_1364)
);

NAND3xp33_ASAP7_75t_SL g1365 ( 
.A(n_1175),
.B(n_28),
.C(n_29),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1151),
.B(n_31),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1210),
.B(n_33),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1149),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1150),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1120),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1097),
.B(n_33),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1214),
.B(n_34),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1141),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1118),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1135),
.Y(n_1375)
);

OR2x2_ASAP7_75t_SL g1376 ( 
.A(n_1117),
.B(n_34),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1101),
.B(n_35),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1139),
.Y(n_1378)
);

INVxp67_ASAP7_75t_SL g1379 ( 
.A(n_1054),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1059),
.B(n_227),
.Y(n_1380)
);

AO22x1_ASAP7_75t_L g1381 ( 
.A1(n_1112),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1203),
.B(n_38),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1146),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1152),
.B(n_1153),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1147),
.Y(n_1385)
);

NOR3xp33_ASAP7_75t_SL g1386 ( 
.A(n_1156),
.B(n_39),
.C(n_40),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1131),
.B(n_230),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1119),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1159),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1058),
.A2(n_233),
.B1(n_234),
.B2(n_232),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1060),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1188),
.A2(n_237),
.B1(n_239),
.B2(n_235),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1189),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1200),
.B(n_39),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1102),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1102),
.B(n_241),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1066),
.B(n_1217),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1133),
.A2(n_243),
.B(n_242),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1145),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1096),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1236),
.B(n_40),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1276),
.A2(n_1391),
.B(n_1397),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1323),
.A2(n_247),
.B(n_246),
.Y(n_1403)
);

AOI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1305),
.A2(n_507),
.B(n_250),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1286),
.A2(n_251),
.B(n_249),
.Y(n_1405)
);

BUFx2_ASAP7_75t_SL g1406 ( 
.A(n_1221),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1273),
.B(n_41),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1260),
.B(n_42),
.Y(n_1408)
);

AO31x2_ASAP7_75t_L g1409 ( 
.A1(n_1248),
.A2(n_45),
.A3(n_43),
.B(n_44),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1345),
.B(n_43),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1347),
.A2(n_254),
.B(n_253),
.Y(n_1411)
);

AOI21x1_ASAP7_75t_SL g1412 ( 
.A1(n_1356),
.A2(n_45),
.B(n_46),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1243),
.A2(n_256),
.B(n_255),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1329),
.A2(n_258),
.B(n_257),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1328),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1242),
.A2(n_262),
.B(n_260),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1349),
.B(n_46),
.Y(n_1417)
);

INVxp67_ASAP7_75t_SL g1418 ( 
.A(n_1380),
.Y(n_1418)
);

AOI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1232),
.A2(n_506),
.B(n_264),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1313),
.B(n_47),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1244),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1312),
.B(n_47),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1315),
.B(n_48),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1380),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1424)
);

NOR3xp33_ASAP7_75t_L g1425 ( 
.A(n_1253),
.B(n_1264),
.C(n_1348),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1231),
.A2(n_1238),
.B(n_1235),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1241),
.A2(n_267),
.B(n_265),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1321),
.B(n_49),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1237),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1336),
.Y(n_1430)
);

AOI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1367),
.A2(n_272),
.B(n_271),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1222),
.B(n_50),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1220),
.Y(n_1433)
);

AND3x2_ASAP7_75t_L g1434 ( 
.A(n_1338),
.B(n_51),
.C(n_52),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1343),
.B(n_52),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1379),
.A2(n_274),
.B(n_273),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1358),
.B(n_53),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1322),
.A2(n_283),
.B(n_280),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1368),
.A2(n_286),
.B(n_285),
.Y(n_1439)
);

AND3x4_ASAP7_75t_L g1440 ( 
.A(n_1292),
.B(n_1257),
.C(n_1332),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1249),
.A2(n_288),
.B(n_287),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1239),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1221),
.Y(n_1443)
);

INVx6_ASAP7_75t_L g1444 ( 
.A(n_1221),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1361),
.B(n_54),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1375),
.A2(n_290),
.B(n_289),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1378),
.A2(n_292),
.B(n_291),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1269),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1293),
.A2(n_302),
.B(n_299),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1293),
.A2(n_306),
.B(n_304),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1280),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1370),
.A2(n_310),
.B(n_308),
.Y(n_1452)
);

AO31x2_ASAP7_75t_L g1453 ( 
.A1(n_1372),
.A2(n_58),
.A3(n_56),
.B(n_57),
.Y(n_1453)
);

AOI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1327),
.A2(n_313),
.B(n_311),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1309),
.B(n_57),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1301),
.A2(n_317),
.B(n_316),
.Y(n_1456)
);

OR2x6_ASAP7_75t_L g1457 ( 
.A(n_1312),
.B(n_318),
.Y(n_1457)
);

AO21x2_ASAP7_75t_L g1458 ( 
.A1(n_1290),
.A2(n_321),
.B(n_320),
.Y(n_1458)
);

O2A1O1Ixp5_ASAP7_75t_L g1459 ( 
.A1(n_1366),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1282),
.B(n_61),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1306),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1298),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1341),
.A2(n_324),
.B(n_323),
.Y(n_1463)
);

INVx4_ASAP7_75t_L g1464 ( 
.A(n_1283),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1357),
.A2(n_326),
.B(n_325),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1240),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1247),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1387),
.A2(n_1355),
.B(n_1374),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1362),
.B(n_62),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1261),
.A2(n_328),
.B(n_327),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1271),
.B(n_505),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1226),
.A2(n_330),
.B(n_329),
.Y(n_1472)
);

AO31x2_ASAP7_75t_L g1473 ( 
.A1(n_1344),
.A2(n_1270),
.A3(n_1390),
.B(n_1274),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1267),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1318),
.B(n_63),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1393),
.A2(n_333),
.B(n_332),
.Y(n_1476)
);

AO31x2_ASAP7_75t_L g1477 ( 
.A1(n_1346),
.A2(n_66),
.A3(n_64),
.B(n_65),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_SL g1478 ( 
.A(n_1271),
.B(n_67),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1272),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1283),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1383),
.B(n_68),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1225),
.A2(n_339),
.B(n_337),
.Y(n_1482)
);

OAI22x1_ASAP7_75t_L g1483 ( 
.A1(n_1330),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1271),
.B(n_340),
.Y(n_1484)
);

A2O1A1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1377),
.A2(n_1369),
.B(n_1351),
.C(n_1398),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1255),
.A2(n_345),
.B(n_343),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1319),
.B(n_70),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1385),
.B(n_1252),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1278),
.A2(n_1300),
.B1(n_1311),
.B2(n_1299),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1314),
.Y(n_1490)
);

OAI21xp33_ASAP7_75t_L g1491 ( 
.A1(n_1363),
.A2(n_72),
.B(n_73),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1339),
.B(n_74),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1340),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1262),
.A2(n_350),
.B(n_348),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1320),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1350),
.B(n_74),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1262),
.A2(n_352),
.B(n_351),
.Y(n_1497)
);

NOR2xp67_ASAP7_75t_L g1498 ( 
.A(n_1281),
.B(n_1389),
.Y(n_1498)
);

OAI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1351),
.A2(n_1228),
.B(n_1224),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1219),
.B(n_353),
.Y(n_1500)
);

XNOR2xp5_ASAP7_75t_L g1501 ( 
.A(n_1400),
.B(n_354),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1384),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1287),
.B(n_75),
.Y(n_1503)
);

AO21x1_ASAP7_75t_L g1504 ( 
.A1(n_1289),
.A2(n_76),
.B(n_78),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1265),
.A2(n_356),
.B(n_355),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1265),
.A2(n_359),
.B(n_358),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1283),
.Y(n_1507)
);

INVx6_ASAP7_75t_SL g1508 ( 
.A(n_1245),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1223),
.A2(n_363),
.B(n_362),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1246),
.Y(n_1510)
);

AOI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1396),
.A2(n_365),
.B(n_364),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1275),
.B(n_78),
.Y(n_1512)
);

INVx4_ASAP7_75t_L g1513 ( 
.A(n_1297),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1219),
.B(n_369),
.Y(n_1514)
);

A2O1A1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1384),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_1515)
);

NAND2x1_ASAP7_75t_L g1516 ( 
.A(n_1297),
.B(n_372),
.Y(n_1516)
);

OAI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1254),
.A2(n_374),
.B(n_373),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1360),
.A2(n_376),
.B(n_375),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1360),
.A2(n_380),
.B(n_378),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1256),
.A2(n_382),
.B(n_381),
.Y(n_1520)
);

A2O1A1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1227),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1304),
.B(n_82),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1307),
.B(n_1310),
.Y(n_1523)
);

AOI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1399),
.A2(n_387),
.B(n_386),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1285),
.B(n_83),
.Y(n_1525)
);

A2O1A1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1353),
.A2(n_86),
.B(n_83),
.C(n_84),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1382),
.B(n_84),
.Y(n_1527)
);

OA21x2_ASAP7_75t_L g1528 ( 
.A1(n_1258),
.A2(n_390),
.B(n_388),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1395),
.A2(n_393),
.B(n_392),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1359),
.B(n_87),
.Y(n_1530)
);

NOR2xp67_ASAP7_75t_SL g1531 ( 
.A(n_1297),
.B(n_87),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1395),
.A2(n_396),
.B(n_394),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1229),
.B(n_88),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1394),
.B(n_88),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_SL g1535 ( 
.A1(n_1333),
.A2(n_399),
.B(n_397),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1291),
.Y(n_1536)
);

OAI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1294),
.A2(n_405),
.B(n_403),
.Y(n_1537)
);

XNOR2xp5_ASAP7_75t_L g1538 ( 
.A(n_1342),
.B(n_407),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1373),
.A2(n_409),
.B(n_408),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1331),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1371),
.B(n_89),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1302),
.A2(n_414),
.B(n_410),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1245),
.Y(n_1543)
);

AOI221x1_ASAP7_75t_L g1544 ( 
.A1(n_1365),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.C(n_94),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1388),
.B(n_92),
.Y(n_1545)
);

AOI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1381),
.A2(n_416),
.B(n_415),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1303),
.A2(n_418),
.B(n_417),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1326),
.B(n_94),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1326),
.B(n_96),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1395),
.A2(n_420),
.B(n_419),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_1298),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1259),
.Y(n_1552)
);

BUFx10_ASAP7_75t_L g1553 ( 
.A(n_1332),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_SL g1554 ( 
.A1(n_1392),
.A2(n_422),
.B(n_421),
.Y(n_1554)
);

O2A1O1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1230),
.A2(n_1277),
.B(n_1279),
.C(n_1308),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1354),
.B(n_96),
.Y(n_1556)
);

INVxp67_ASAP7_75t_L g1557 ( 
.A(n_1263),
.Y(n_1557)
);

AOI21xp33_ASAP7_75t_L g1558 ( 
.A1(n_1354),
.A2(n_97),
.B(n_98),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1233),
.B(n_98),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1337),
.A2(n_427),
.B(n_425),
.Y(n_1560)
);

BUFx4_ASAP7_75t_SL g1561 ( 
.A(n_1295),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1425),
.B(n_1233),
.Y(n_1562)
);

OAI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1402),
.A2(n_1468),
.B(n_1414),
.Y(n_1563)
);

AOI21xp33_ASAP7_75t_L g1564 ( 
.A1(n_1426),
.A2(n_1266),
.B(n_1337),
.Y(n_1564)
);

OAI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1485),
.A2(n_1266),
.B(n_1386),
.Y(n_1565)
);

OR2x6_ASAP7_75t_L g1566 ( 
.A(n_1406),
.B(n_1250),
.Y(n_1566)
);

CKINVDCx20_ASAP7_75t_R g1567 ( 
.A(n_1421),
.Y(n_1567)
);

BUFx4f_ASAP7_75t_SL g1568 ( 
.A(n_1508),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1418),
.A2(n_1268),
.B(n_1250),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1542),
.A2(n_1352),
.B(n_1317),
.Y(n_1570)
);

OAI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1432),
.A2(n_1352),
.B(n_1268),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1523),
.A2(n_1352),
.B(n_1334),
.Y(n_1572)
);

AO31x2_ASAP7_75t_L g1573 ( 
.A1(n_1504),
.A2(n_1381),
.A3(n_1376),
.B(n_1335),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1415),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1407),
.B(n_1316),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1488),
.B(n_1288),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1408),
.B(n_1298),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1557),
.A2(n_1251),
.B1(n_1335),
.B2(n_1325),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1429),
.B(n_1317),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1491),
.A2(n_1296),
.B1(n_1364),
.B2(n_1325),
.Y(n_1580)
);

INVx5_ASAP7_75t_L g1581 ( 
.A(n_1480),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1480),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1495),
.Y(n_1583)
);

INVx4_ASAP7_75t_L g1584 ( 
.A(n_1480),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1496),
.B(n_1284),
.Y(n_1585)
);

AO31x2_ASAP7_75t_L g1586 ( 
.A1(n_1544),
.A2(n_1335),
.A3(n_1325),
.B(n_1324),
.Y(n_1586)
);

AOI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1479),
.A2(n_1234),
.B1(n_1324),
.B2(n_103),
.C(n_104),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1476),
.A2(n_1324),
.B(n_432),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1507),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1449),
.A2(n_433),
.B(n_431),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1527),
.B(n_101),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1450),
.A2(n_435),
.B(n_434),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1507),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1403),
.A2(n_437),
.B(n_436),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1430),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1493),
.B(n_438),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1530),
.B(n_101),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1541),
.B(n_102),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1464),
.B(n_1457),
.Y(n_1599)
);

AO21x1_ASAP7_75t_L g1600 ( 
.A1(n_1424),
.A2(n_102),
.B(n_103),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1461),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1448),
.Y(n_1602)
);

OA22x2_ASAP7_75t_L g1603 ( 
.A1(n_1434),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1482),
.A2(n_502),
.B(n_440),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1513),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1451),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1464),
.B(n_439),
.Y(n_1607)
);

OAI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1456),
.A2(n_444),
.B(n_443),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1499),
.B(n_105),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1423),
.B(n_107),
.Y(n_1610)
);

AOI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1546),
.A2(n_446),
.B(n_445),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1442),
.Y(n_1612)
);

A2O1A1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1555),
.A2(n_107),
.B(n_108),
.C(n_110),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1427),
.A2(n_499),
.B(n_447),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1422),
.B(n_450),
.Y(n_1615)
);

OAI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1486),
.A2(n_452),
.B(n_451),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1441),
.A2(n_1470),
.B(n_1517),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1443),
.B(n_453),
.Y(n_1618)
);

A2O1A1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1522),
.A2(n_108),
.B(n_111),
.C(n_112),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1520),
.A2(n_457),
.B(n_454),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1494),
.A2(n_498),
.B(n_497),
.Y(n_1621)
);

O2A1O1Ixp33_ASAP7_75t_SL g1622 ( 
.A1(n_1521),
.A2(n_111),
.B(n_112),
.C(n_113),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1512),
.B(n_113),
.Y(n_1623)
);

INVx3_ASAP7_75t_L g1624 ( 
.A(n_1513),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1537),
.A2(n_496),
.B(n_492),
.Y(n_1625)
);

OA21x2_ASAP7_75t_L g1626 ( 
.A1(n_1463),
.A2(n_490),
.B(n_489),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1540),
.Y(n_1627)
);

O2A1O1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1515),
.A2(n_114),
.B(n_116),
.C(n_117),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1428),
.B(n_116),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1435),
.B(n_117),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1487),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1444),
.Y(n_1632)
);

OAI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1497),
.A2(n_484),
.B(n_482),
.Y(n_1633)
);

AOI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1440),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1405),
.A2(n_479),
.B(n_478),
.Y(n_1635)
);

A2O1A1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1526),
.A2(n_119),
.B(n_120),
.C(n_121),
.Y(n_1636)
);

AO31x2_ASAP7_75t_L g1637 ( 
.A1(n_1438),
.A2(n_477),
.A3(n_476),
.B(n_475),
.Y(n_1637)
);

A2O1A1Ixp33_ASAP7_75t_L g1638 ( 
.A1(n_1472),
.A2(n_121),
.B(n_122),
.C(n_123),
.Y(n_1638)
);

AO21x2_ASAP7_75t_L g1639 ( 
.A1(n_1431),
.A2(n_474),
.B(n_473),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1552),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1452),
.A2(n_472),
.B(n_471),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1507),
.Y(n_1642)
);

INVxp67_ASAP7_75t_SL g1643 ( 
.A(n_1552),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_R g1644 ( 
.A1(n_1483),
.A2(n_1490),
.B1(n_1467),
.B2(n_1466),
.Y(n_1644)
);

A2O1A1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1534),
.A2(n_122),
.B(n_123),
.C(n_124),
.Y(n_1645)
);

OAI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1505),
.A2(n_470),
.B(n_469),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1465),
.A2(n_467),
.B(n_466),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1436),
.A2(n_461),
.B(n_460),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1525),
.B(n_124),
.Y(n_1649)
);

A2O1A1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1511),
.A2(n_125),
.B(n_126),
.C(n_127),
.Y(n_1650)
);

INVx3_ASAP7_75t_SL g1651 ( 
.A(n_1444),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1506),
.A2(n_125),
.B(n_127),
.Y(n_1652)
);

OAI21x1_ASAP7_75t_L g1653 ( 
.A1(n_1416),
.A2(n_128),
.B(n_129),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1437),
.B(n_128),
.Y(n_1654)
);

O2A1O1Ixp5_ASAP7_75t_SL g1655 ( 
.A1(n_1558),
.A2(n_210),
.B(n_131),
.C(n_132),
.Y(n_1655)
);

AO31x2_ASAP7_75t_L g1656 ( 
.A1(n_1489),
.A2(n_210),
.A3(n_131),
.B(n_132),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1498),
.B(n_130),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_1410),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1445),
.B(n_133),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1433),
.Y(n_1660)
);

O2A1O1Ixp33_ASAP7_75t_SL g1661 ( 
.A1(n_1516),
.A2(n_133),
.B(n_134),
.C(n_135),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1439),
.A2(n_1447),
.B(n_1446),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1528),
.A2(n_209),
.B(n_136),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1533),
.B(n_135),
.Y(n_1664)
);

AO21x2_ASAP7_75t_L g1665 ( 
.A1(n_1535),
.A2(n_136),
.B(n_137),
.Y(n_1665)
);

BUFx2_ASAP7_75t_L g1666 ( 
.A(n_1508),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1561),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1469),
.B(n_138),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_SL g1669 ( 
.A1(n_1503),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1528),
.A2(n_209),
.B(n_145),
.Y(n_1670)
);

INVx4_ASAP7_75t_L g1671 ( 
.A(n_1551),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1481),
.B(n_1401),
.Y(n_1672)
);

CKINVDCx20_ASAP7_75t_R g1673 ( 
.A(n_1501),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1536),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1543),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_1675)
);

INVx2_ASAP7_75t_SL g1676 ( 
.A(n_1553),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1548),
.B(n_146),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1560),
.A2(n_148),
.B(n_149),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1459),
.A2(n_150),
.B(n_151),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1559),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1529),
.A2(n_155),
.B(n_156),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_SL g1682 ( 
.A1(n_1471),
.A2(n_157),
.B(n_158),
.Y(n_1682)
);

AOI221xp5_ASAP7_75t_L g1683 ( 
.A1(n_1420),
.A2(n_1460),
.B1(n_1474),
.B2(n_1475),
.C(n_1502),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1510),
.B(n_158),
.Y(n_1684)
);

AO31x2_ASAP7_75t_L g1685 ( 
.A1(n_1536),
.A2(n_159),
.A3(n_160),
.B(n_161),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1411),
.A2(n_162),
.B(n_163),
.Y(n_1686)
);

NOR2x1_ASAP7_75t_L g1687 ( 
.A(n_1545),
.B(n_164),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1532),
.A2(n_208),
.B(n_165),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1492),
.Y(n_1689)
);

OAI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1549),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_1690)
);

INVx1_ASAP7_75t_SL g1691 ( 
.A(n_1583),
.Y(n_1691)
);

BUFx12f_ASAP7_75t_L g1692 ( 
.A(n_1667),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_SL g1693 ( 
.A1(n_1565),
.A2(n_1554),
.B1(n_1500),
.B2(n_1514),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_SL g1694 ( 
.A1(n_1634),
.A2(n_1556),
.B1(n_1538),
.B2(n_1457),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1617),
.A2(n_1478),
.B(n_1550),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_SL g1696 ( 
.A1(n_1562),
.A2(n_1500),
.B1(n_1514),
.B2(n_1455),
.Y(n_1696)
);

BUFx8_ASAP7_75t_L g1697 ( 
.A(n_1666),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1587),
.A2(n_1531),
.B1(n_1471),
.B2(n_1484),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1683),
.A2(n_1484),
.B1(n_1417),
.B2(n_1553),
.Y(n_1699)
);

OAI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1580),
.A2(n_1462),
.B1(n_1551),
.B2(n_1419),
.Y(n_1700)
);

INVx4_ASAP7_75t_L g1701 ( 
.A(n_1581),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1644),
.A2(n_1600),
.B1(n_1677),
.B2(n_1668),
.Y(n_1702)
);

CKINVDCx11_ASAP7_75t_R g1703 ( 
.A(n_1567),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1615),
.A2(n_1458),
.B1(n_1547),
.B2(n_1518),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1651),
.Y(n_1705)
);

INVx2_ASAP7_75t_SL g1706 ( 
.A(n_1632),
.Y(n_1706)
);

INVx5_ASAP7_75t_L g1707 ( 
.A(n_1566),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1585),
.A2(n_1462),
.B1(n_1551),
.B2(n_1404),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1609),
.A2(n_1519),
.B1(n_1539),
.B2(n_1413),
.Y(n_1709)
);

CKINVDCx16_ASAP7_75t_R g1710 ( 
.A(n_1673),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1575),
.A2(n_1454),
.B1(n_1524),
.B2(n_1412),
.Y(n_1711)
);

OAI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1576),
.A2(n_1473),
.B1(n_1409),
.B2(n_1477),
.Y(n_1712)
);

OAI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1603),
.A2(n_1409),
.B1(n_1473),
.B2(n_1477),
.Y(n_1713)
);

NAND2x1p5_ASAP7_75t_L g1714 ( 
.A(n_1581),
.B(n_1509),
.Y(n_1714)
);

BUFx10_ASAP7_75t_L g1715 ( 
.A(n_1596),
.Y(n_1715)
);

CKINVDCx11_ASAP7_75t_R g1716 ( 
.A(n_1631),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1658),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1627),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1690),
.A2(n_1680),
.B1(n_1687),
.B2(n_1678),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1640),
.Y(n_1720)
);

INVx3_ASAP7_75t_SL g1721 ( 
.A(n_1579),
.Y(n_1721)
);

BUFx2_ASAP7_75t_L g1722 ( 
.A(n_1627),
.Y(n_1722)
);

BUFx6f_ASAP7_75t_L g1723 ( 
.A(n_1582),
.Y(n_1723)
);

INVx5_ASAP7_75t_L g1724 ( 
.A(n_1566),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_SL g1725 ( 
.A1(n_1572),
.A2(n_1453),
.B1(n_168),
.B2(n_169),
.Y(n_1725)
);

CKINVDCx6p67_ASAP7_75t_R g1726 ( 
.A(n_1581),
.Y(n_1726)
);

BUFx4f_ASAP7_75t_SL g1727 ( 
.A(n_1582),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1664),
.A2(n_1453),
.B1(n_168),
.B2(n_169),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1672),
.A2(n_1453),
.B1(n_170),
.B2(n_171),
.Y(n_1729)
);

CKINVDCx20_ASAP7_75t_R g1730 ( 
.A(n_1568),
.Y(n_1730)
);

CKINVDCx20_ASAP7_75t_R g1731 ( 
.A(n_1666),
.Y(n_1731)
);

INVx5_ASAP7_75t_L g1732 ( 
.A(n_1589),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1689),
.A2(n_167),
.B1(n_170),
.B2(n_171),
.Y(n_1733)
);

INVx6_ASAP7_75t_L g1734 ( 
.A(n_1589),
.Y(n_1734)
);

OAI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1569),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_1735)
);

BUFx4f_ASAP7_75t_SL g1736 ( 
.A(n_1593),
.Y(n_1736)
);

INVx6_ASAP7_75t_L g1737 ( 
.A(n_1593),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1674),
.Y(n_1738)
);

INVx6_ASAP7_75t_L g1739 ( 
.A(n_1642),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1564),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_SL g1741 ( 
.A1(n_1604),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1669),
.A2(n_1614),
.B1(n_1594),
.B2(n_1679),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1577),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1642),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_SL g1745 ( 
.A1(n_1571),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_1745)
);

CKINVDCx6p67_ASAP7_75t_R g1746 ( 
.A(n_1584),
.Y(n_1746)
);

BUFx3_ASAP7_75t_L g1747 ( 
.A(n_1612),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1574),
.Y(n_1748)
);

INVx6_ASAP7_75t_L g1749 ( 
.A(n_1671),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1606),
.Y(n_1750)
);

CKINVDCx11_ASAP7_75t_R g1751 ( 
.A(n_1657),
.Y(n_1751)
);

BUFx8_ASAP7_75t_L g1752 ( 
.A(n_1597),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1681),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_1599),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1688),
.A2(n_184),
.B1(n_186),
.B2(n_188),
.Y(n_1755)
);

INVxp67_ASAP7_75t_SL g1756 ( 
.A(n_1643),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1595),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1660),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1665),
.A2(n_1591),
.B1(n_1620),
.B2(n_1625),
.Y(n_1759)
);

BUFx12f_ASAP7_75t_L g1760 ( 
.A(n_1676),
.Y(n_1760)
);

OAI22xp5_ASAP7_75t_SL g1761 ( 
.A1(n_1610),
.A2(n_208),
.B1(n_190),
.B2(n_191),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1601),
.B(n_207),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1684),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1685),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_1602),
.Y(n_1765)
);

BUFx2_ASAP7_75t_L g1766 ( 
.A(n_1599),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1629),
.B(n_207),
.Y(n_1767)
);

BUFx8_ASAP7_75t_L g1768 ( 
.A(n_1598),
.Y(n_1768)
);

CKINVDCx6p67_ASAP7_75t_R g1769 ( 
.A(n_1618),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1630),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1654),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_SL g1772 ( 
.A1(n_1659),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1578),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1613),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1605),
.Y(n_1775)
);

BUFx6f_ASAP7_75t_L g1776 ( 
.A(n_1624),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1718),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1748),
.Y(n_1778)
);

CKINVDCx20_ASAP7_75t_R g1779 ( 
.A(n_1703),
.Y(n_1779)
);

BUFx3_ASAP7_75t_L g1780 ( 
.A(n_1707),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1757),
.Y(n_1781)
);

CKINVDCx14_ASAP7_75t_R g1782 ( 
.A(n_1730),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1712),
.B(n_1656),
.Y(n_1783)
);

CKINVDCx6p67_ASAP7_75t_R g1784 ( 
.A(n_1692),
.Y(n_1784)
);

INVx2_ASAP7_75t_SL g1785 ( 
.A(n_1722),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1758),
.B(n_1623),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_L g1787 ( 
.A(n_1707),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1738),
.B(n_1563),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1764),
.B(n_1720),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1756),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1750),
.B(n_1649),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1763),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1714),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1713),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1711),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1707),
.B(n_1570),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1708),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1724),
.B(n_1588),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1747),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1695),
.Y(n_1800)
);

O2A1O1Ixp33_ASAP7_75t_L g1801 ( 
.A1(n_1774),
.A2(n_1636),
.B(n_1619),
.C(n_1645),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1724),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1717),
.B(n_1573),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1721),
.B(n_1586),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1724),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1766),
.B(n_1573),
.Y(n_1806)
);

AOI21x1_ASAP7_75t_L g1807 ( 
.A1(n_1735),
.A2(n_1611),
.B(n_1663),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1775),
.Y(n_1808)
);

INVx2_ASAP7_75t_SL g1809 ( 
.A(n_1754),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1709),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1691),
.B(n_1670),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1716),
.Y(n_1812)
);

OAI21x1_ASAP7_75t_L g1813 ( 
.A1(n_1704),
.A2(n_1662),
.B(n_1652),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1776),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1789),
.B(n_1725),
.Y(n_1815)
);

OR2x6_ASAP7_75t_L g1816 ( 
.A(n_1796),
.B(n_1682),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_1777),
.Y(n_1817)
);

BUFx2_ASAP7_75t_L g1818 ( 
.A(n_1796),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_1787),
.Y(n_1819)
);

BUFx2_ASAP7_75t_L g1820 ( 
.A(n_1796),
.Y(n_1820)
);

BUFx2_ASAP7_75t_L g1821 ( 
.A(n_1796),
.Y(n_1821)
);

BUFx2_ASAP7_75t_L g1822 ( 
.A(n_1802),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1789),
.B(n_1759),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1789),
.B(n_1702),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_1812),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1785),
.Y(n_1826)
);

AO21x2_ASAP7_75t_L g1827 ( 
.A1(n_1795),
.A2(n_1810),
.B(n_1813),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1783),
.B(n_1762),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1778),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1788),
.Y(n_1830)
);

BUFx2_ASAP7_75t_L g1831 ( 
.A(n_1802),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1781),
.B(n_1728),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1781),
.Y(n_1833)
);

AOI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1794),
.A2(n_1694),
.B1(n_1761),
.B2(n_1742),
.Y(n_1834)
);

AO21x2_ASAP7_75t_L g1835 ( 
.A1(n_1795),
.A2(n_1810),
.B(n_1800),
.Y(n_1835)
);

BUFx6f_ASAP7_75t_L g1836 ( 
.A(n_1787),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_R g1837 ( 
.A(n_1779),
.B(n_1705),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1829),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1818),
.B(n_1785),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1818),
.B(n_1799),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1833),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1820),
.B(n_1799),
.Y(n_1842)
);

AND2x4_ASAP7_75t_L g1843 ( 
.A(n_1820),
.B(n_1780),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1835),
.B(n_1783),
.Y(n_1844)
);

OAI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1834),
.A2(n_1794),
.B1(n_1800),
.B2(n_1811),
.Y(n_1845)
);

BUFx3_ASAP7_75t_L g1846 ( 
.A(n_1822),
.Y(n_1846)
);

HB1xp67_ASAP7_75t_L g1847 ( 
.A(n_1817),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1829),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1821),
.B(n_1804),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1829),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1835),
.B(n_1790),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1821),
.B(n_1804),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1835),
.B(n_1790),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1828),
.B(n_1824),
.Y(n_1854)
);

INVx1_ASAP7_75t_SL g1855 ( 
.A(n_1825),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1824),
.A2(n_1741),
.B1(n_1745),
.B2(n_1719),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1841),
.Y(n_1857)
);

BUFx2_ASAP7_75t_L g1858 ( 
.A(n_1846),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1838),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1838),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1848),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1849),
.B(n_1830),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1848),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1850),
.Y(n_1864)
);

INVx5_ASAP7_75t_L g1865 ( 
.A(n_1843),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1849),
.B(n_1830),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1857),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1858),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1865),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1865),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1860),
.Y(n_1871)
);

BUFx3_ASAP7_75t_L g1872 ( 
.A(n_1865),
.Y(n_1872)
);

AND2x4_ASAP7_75t_L g1873 ( 
.A(n_1868),
.B(n_1872),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1867),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1867),
.B(n_1854),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1871),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1869),
.B(n_1865),
.Y(n_1877)
);

NOR2xp67_ASAP7_75t_L g1878 ( 
.A(n_1870),
.B(n_1847),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1871),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1868),
.B(n_1828),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1868),
.B(n_1845),
.Y(n_1881)
);

AOI221x1_ASAP7_75t_SL g1882 ( 
.A1(n_1873),
.A2(n_1791),
.B1(n_1786),
.B2(n_1767),
.C(n_1675),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1874),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1873),
.A2(n_1834),
.B1(n_1816),
.B2(n_1815),
.Y(n_1884)
);

NAND2xp33_ASAP7_75t_SL g1885 ( 
.A(n_1881),
.B(n_1837),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1876),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1878),
.B(n_1877),
.Y(n_1887)
);

NAND2xp33_ASAP7_75t_SL g1888 ( 
.A(n_1880),
.B(n_1731),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1875),
.B(n_1855),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1879),
.B(n_1840),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1873),
.B(n_1840),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1873),
.B(n_1842),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1887),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1886),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1883),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1882),
.B(n_1852),
.Y(n_1896)
);

OAI21xp33_ASAP7_75t_L g1897 ( 
.A1(n_1884),
.A2(n_1856),
.B(n_1772),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1889),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1891),
.B(n_1784),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1890),
.Y(n_1900)
);

OAI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1896),
.A2(n_1892),
.B1(n_1893),
.B2(n_1898),
.Y(n_1901)
);

OAI322xp33_ASAP7_75t_L g1902 ( 
.A1(n_1894),
.A2(n_1844),
.A3(n_1853),
.B1(n_1851),
.B2(n_1733),
.C1(n_1743),
.C2(n_1812),
.Y(n_1902)
);

AOI32xp33_ASAP7_75t_L g1903 ( 
.A1(n_1897),
.A2(n_1885),
.A3(n_1888),
.B1(n_1815),
.B2(n_1843),
.Y(n_1903)
);

AOI21xp33_ASAP7_75t_L g1904 ( 
.A1(n_1899),
.A2(n_1811),
.B(n_1768),
.Y(n_1904)
);

INVx3_ASAP7_75t_L g1905 ( 
.A(n_1904),
.Y(n_1905)
);

AOI221xp5_ASAP7_75t_L g1906 ( 
.A1(n_1901),
.A2(n_1897),
.B1(n_1895),
.B2(n_1900),
.C(n_1801),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1902),
.Y(n_1907)
);

OAI31xp33_ASAP7_75t_L g1908 ( 
.A1(n_1903),
.A2(n_1782),
.A3(n_1650),
.B(n_1638),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1905),
.B(n_1784),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1907),
.Y(n_1910)
);

NAND4xp25_ASAP7_75t_L g1911 ( 
.A(n_1906),
.B(n_1698),
.C(n_1770),
.D(n_1771),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1908),
.B(n_1710),
.Y(n_1912)
);

NAND5xp2_ASAP7_75t_L g1913 ( 
.A(n_1906),
.B(n_1696),
.C(n_1699),
.D(n_1740),
.E(n_1628),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1910),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1912),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1911),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1909),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1913),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1910),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1910),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1910),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1910),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1912),
.Y(n_1923)
);

NOR2xp33_ASAP7_75t_L g1924 ( 
.A(n_1915),
.B(n_1923),
.Y(n_1924)
);

INVx2_ASAP7_75t_SL g1925 ( 
.A(n_1917),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1914),
.B(n_1862),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1919),
.Y(n_1927)
);

AO22x2_ASAP7_75t_L g1928 ( 
.A1(n_1920),
.A2(n_1706),
.B1(n_1861),
.B2(n_1860),
.Y(n_1928)
);

NOR3xp33_ASAP7_75t_L g1929 ( 
.A(n_1921),
.B(n_1751),
.C(n_1765),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1922),
.B(n_1697),
.Y(n_1930)
);

NOR2x1p5_ASAP7_75t_SL g1931 ( 
.A(n_1918),
.B(n_1861),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1916),
.B(n_1859),
.Y(n_1932)
);

NOR2x1_ASAP7_75t_L g1933 ( 
.A(n_1914),
.B(n_1607),
.Y(n_1933)
);

NOR3x1_ASAP7_75t_L g1934 ( 
.A(n_1915),
.B(n_1697),
.C(n_1822),
.Y(n_1934)
);

NOR3xp33_ASAP7_75t_L g1935 ( 
.A(n_1915),
.B(n_1607),
.C(n_1661),
.Y(n_1935)
);

NAND4xp25_ASAP7_75t_L g1936 ( 
.A(n_1924),
.B(n_1753),
.C(n_1755),
.D(n_1729),
.Y(n_1936)
);

OAI211xp5_ASAP7_75t_L g1937 ( 
.A1(n_1930),
.A2(n_1927),
.B(n_1925),
.C(n_1932),
.Y(n_1937)
);

NAND3xp33_ASAP7_75t_L g1938 ( 
.A(n_1929),
.B(n_1768),
.C(n_1752),
.Y(n_1938)
);

NOR3xp33_ASAP7_75t_L g1939 ( 
.A(n_1933),
.B(n_1635),
.C(n_1648),
.Y(n_1939)
);

NAND3xp33_ASAP7_75t_L g1940 ( 
.A(n_1926),
.B(n_1752),
.C(n_1655),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1934),
.Y(n_1941)
);

AOI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1935),
.A2(n_1760),
.B1(n_1773),
.B2(n_1746),
.Y(n_1942)
);

AOI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1928),
.A2(n_1843),
.B1(n_1727),
.B2(n_1736),
.Y(n_1943)
);

NOR3x1_ASAP7_75t_SL g1944 ( 
.A(n_1931),
.B(n_197),
.C(n_198),
.Y(n_1944)
);

OAI321xp33_ASAP7_75t_L g1945 ( 
.A1(n_1928),
.A2(n_1836),
.A3(n_1819),
.B1(n_1816),
.B2(n_1803),
.C(n_1844),
.Y(n_1945)
);

NOR2xp67_ASAP7_75t_SL g1946 ( 
.A(n_1925),
.B(n_1749),
.Y(n_1946)
);

OAI211xp5_ASAP7_75t_SL g1947 ( 
.A1(n_1924),
.A2(n_1647),
.B(n_1641),
.C(n_1693),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1944),
.Y(n_1948)
);

BUFx2_ASAP7_75t_L g1949 ( 
.A(n_1941),
.Y(n_1949)
);

NAND5xp2_ASAP7_75t_L g1950 ( 
.A(n_1937),
.B(n_1622),
.C(n_1823),
.D(n_1832),
.E(n_202),
.Y(n_1950)
);

NAND4xp25_ASAP7_75t_SL g1951 ( 
.A(n_1942),
.B(n_1655),
.C(n_1852),
.D(n_1839),
.Y(n_1951)
);

NOR5xp2_ASAP7_75t_L g1952 ( 
.A(n_1938),
.B(n_198),
.C(n_199),
.D(n_201),
.E(n_202),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1943),
.Y(n_1953)
);

OAI211xp5_ASAP7_75t_SL g1954 ( 
.A1(n_1946),
.A2(n_203),
.B(n_204),
.C(n_205),
.Y(n_1954)
);

OAI211xp5_ASAP7_75t_L g1955 ( 
.A1(n_1940),
.A2(n_1701),
.B(n_1732),
.C(n_205),
.Y(n_1955)
);

AOI221xp5_ASAP7_75t_L g1956 ( 
.A1(n_1945),
.A2(n_1846),
.B1(n_1831),
.B2(n_1744),
.C(n_1819),
.Y(n_1956)
);

OAI211xp5_ASAP7_75t_SL g1957 ( 
.A1(n_1939),
.A2(n_206),
.B(n_1700),
.C(n_1805),
.Y(n_1957)
);

NOR3xp33_ASAP7_75t_L g1958 ( 
.A(n_1936),
.B(n_1701),
.C(n_1805),
.Y(n_1958)
);

INVx5_ASAP7_75t_L g1959 ( 
.A(n_1949),
.Y(n_1959)
);

INVx2_ASAP7_75t_SL g1960 ( 
.A(n_1948),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1954),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1953),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1955),
.Y(n_1963)
);

NAND4xp75_ASAP7_75t_L g1964 ( 
.A(n_1956),
.B(n_1947),
.C(n_206),
.D(n_1839),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1958),
.B(n_1863),
.Y(n_1965)
);

NOR2x1_ASAP7_75t_L g1966 ( 
.A(n_1950),
.B(n_1723),
.Y(n_1966)
);

OAI21xp5_ASAP7_75t_SL g1967 ( 
.A1(n_1957),
.A2(n_1952),
.B(n_1951),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1949),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1948),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1948),
.B(n_1862),
.Y(n_1970)
);

HB1xp67_ASAP7_75t_L g1971 ( 
.A(n_1948),
.Y(n_1971)
);

NAND4xp75_ASAP7_75t_L g1972 ( 
.A(n_1948),
.B(n_1866),
.C(n_1726),
.D(n_1864),
.Y(n_1972)
);

INVx2_ASAP7_75t_SL g1973 ( 
.A(n_1959),
.Y(n_1973)
);

NOR3xp33_ASAP7_75t_L g1974 ( 
.A(n_1960),
.B(n_1805),
.C(n_1653),
.Y(n_1974)
);

AND2x4_ASAP7_75t_L g1975 ( 
.A(n_1970),
.B(n_1866),
.Y(n_1975)
);

NAND2xp33_ASAP7_75t_SL g1976 ( 
.A(n_1962),
.B(n_1723),
.Y(n_1976)
);

XNOR2xp5_ASAP7_75t_L g1977 ( 
.A(n_1971),
.B(n_1816),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1959),
.B(n_1842),
.Y(n_1978)
);

AND2x4_ASAP7_75t_SL g1979 ( 
.A(n_1969),
.B(n_1769),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1959),
.B(n_1831),
.Y(n_1980)
);

INVx1_ASAP7_75t_SL g1981 ( 
.A(n_1968),
.Y(n_1981)
);

NOR2xp67_ASAP7_75t_L g1982 ( 
.A(n_1963),
.B(n_1732),
.Y(n_1982)
);

AND2x4_ASAP7_75t_L g1983 ( 
.A(n_1966),
.B(n_1826),
.Y(n_1983)
);

INVxp67_ASAP7_75t_L g1984 ( 
.A(n_1961),
.Y(n_1984)
);

NOR3x1_ASAP7_75t_L g1985 ( 
.A(n_1967),
.B(n_1853),
.C(n_1851),
.Y(n_1985)
);

AND2x4_ASAP7_75t_L g1986 ( 
.A(n_1965),
.B(n_1819),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_L g1987 ( 
.A(n_1973),
.Y(n_1987)
);

NAND4xp75_ASAP7_75t_L g1988 ( 
.A(n_1982),
.B(n_1964),
.C(n_1972),
.D(n_1626),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1978),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1980),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1975),
.Y(n_1991)
);

NOR3xp33_ASAP7_75t_SL g1992 ( 
.A(n_1976),
.B(n_1749),
.C(n_1797),
.Y(n_1992)
);

OAI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1981),
.A2(n_1737),
.B1(n_1739),
.B2(n_1734),
.Y(n_1993)
);

BUFx2_ASAP7_75t_L g1994 ( 
.A(n_1983),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1977),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1979),
.Y(n_1996)
);

AOI22xp5_ASAP7_75t_L g1997 ( 
.A1(n_1987),
.A2(n_1984),
.B1(n_1986),
.B2(n_1974),
.Y(n_1997)
);

AOI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1994),
.A2(n_1985),
.B1(n_1734),
.B2(n_1737),
.Y(n_1998)
);

OAI22xp5_ASAP7_75t_SL g1999 ( 
.A1(n_1991),
.A2(n_1739),
.B1(n_1732),
.B2(n_1723),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1996),
.Y(n_2000)
);

OA22x2_ASAP7_75t_L g2001 ( 
.A1(n_1989),
.A2(n_1816),
.B1(n_1814),
.B2(n_1809),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1988),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1990),
.Y(n_2003)
);

OAI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1995),
.A2(n_1819),
.B1(n_1836),
.B2(n_1816),
.Y(n_2004)
);

AOI22xp33_ASAP7_75t_L g2005 ( 
.A1(n_1993),
.A2(n_1836),
.B1(n_1819),
.B2(n_1776),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_2000),
.Y(n_2006)
);

OAI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1998),
.A2(n_1992),
.B1(n_1819),
.B2(n_1836),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_2003),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_1999),
.Y(n_2009)
);

OAI22xp5_ASAP7_75t_SL g2010 ( 
.A1(n_2002),
.A2(n_1776),
.B1(n_1787),
.B2(n_1780),
.Y(n_2010)
);

OAI21xp33_ASAP7_75t_L g2011 ( 
.A1(n_1997),
.A2(n_1780),
.B(n_1836),
.Y(n_2011)
);

OA21x2_ASAP7_75t_L g2012 ( 
.A1(n_2005),
.A2(n_1686),
.B(n_1590),
.Y(n_2012)
);

AOI22xp5_ASAP7_75t_L g2013 ( 
.A1(n_2004),
.A2(n_1836),
.B1(n_1787),
.B2(n_1715),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_2008),
.Y(n_2014)
);

AOI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_2006),
.A2(n_2001),
.B1(n_1787),
.B2(n_1715),
.Y(n_2015)
);

AOI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_2011),
.A2(n_1809),
.B1(n_1827),
.B2(n_1639),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_2009),
.A2(n_1792),
.B(n_1808),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_2007),
.B(n_1637),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_2010),
.Y(n_2019)
);

AOI31xp33_ASAP7_75t_L g2020 ( 
.A1(n_2013),
.A2(n_1798),
.A3(n_1832),
.B(n_1793),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_2014),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_2015),
.B(n_2012),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_R g2023 ( 
.A(n_2019),
.B(n_1807),
.Y(n_2023)
);

XNOR2xp5_ASAP7_75t_L g2024 ( 
.A(n_2017),
.B(n_1823),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2018),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_2020),
.Y(n_2026)
);

AOI22xp5_ASAP7_75t_L g2027 ( 
.A1(n_2021),
.A2(n_2016),
.B1(n_1827),
.B2(n_1798),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_2026),
.B(n_1793),
.Y(n_2028)
);

AOI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_2022),
.A2(n_1626),
.B(n_1621),
.Y(n_2029)
);

OAI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_2028),
.A2(n_2025),
.B1(n_2027),
.B2(n_2024),
.Y(n_2030)
);

AOI31xp33_ASAP7_75t_L g2031 ( 
.A1(n_2029),
.A2(n_2023),
.A3(n_1798),
.B(n_1792),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_2030),
.A2(n_1616),
.B(n_1633),
.Y(n_2032)
);

AOI22xp33_ASAP7_75t_L g2033 ( 
.A1(n_2032),
.A2(n_2031),
.B1(n_1827),
.B2(n_1808),
.Y(n_2033)
);

AOI22xp5_ASAP7_75t_L g2034 ( 
.A1(n_2033),
.A2(n_1798),
.B1(n_1797),
.B2(n_1806),
.Y(n_2034)
);

AOI211xp5_ASAP7_75t_L g2035 ( 
.A1(n_2034),
.A2(n_1646),
.B(n_1592),
.C(n_1608),
.Y(n_2035)
);


endmodule