module fake_jpeg_15639_n_251 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_36),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_13),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_41),
.Y(n_62)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_27),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_18),
.B1(n_23),
.B2(n_28),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_51),
.B1(n_52),
.B2(n_42),
.Y(n_81)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_31),
.B(n_23),
.C(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_49),
.B(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_18),
.B1(n_31),
.B2(n_30),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_21),
.B1(n_17),
.B2(n_26),
.Y(n_52)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_63),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_21),
.B1(n_19),
.B2(n_29),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_42),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_19),
.B1(n_29),
.B2(n_15),
.Y(n_61)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_33),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_72),
.Y(n_110)
);

CKINVDCx6p67_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_68),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_81),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_56),
.B1(n_27),
.B2(n_25),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_38),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_75),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_64),
.B1(n_45),
.B2(n_54),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_74),
.A2(n_83),
.B1(n_78),
.B2(n_55),
.Y(n_100)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_41),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_47),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_42),
.B1(n_39),
.B2(n_15),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_79),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_39),
.B1(n_1),
.B2(n_2),
.Y(n_83)
);

CKINVDCx6p67_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_84),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_50),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_72),
.C(n_46),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_74),
.C(n_81),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_95),
.Y(n_119)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_99),
.Y(n_128)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_107),
.B1(n_85),
.B2(n_59),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_63),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_100),
.A2(n_59),
.B1(n_39),
.B2(n_25),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_49),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_25),
.B(n_2),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_33),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_106),
.Y(n_129)
);

CKINVDCx12_ASAP7_75t_R g106 ( 
.A(n_68),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_58),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_127),
.C(n_107),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_77),
.B1(n_87),
.B2(n_55),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_115),
.A2(n_117),
.B1(n_98),
.B2(n_92),
.Y(n_137)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_77),
.B1(n_87),
.B2(n_76),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_118),
.B(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_73),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_103),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_122),
.A2(n_103),
.B1(n_97),
.B2(n_106),
.Y(n_148)
);

A2O1A1O1Ixp25_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_104),
.B(n_93),
.C(n_110),
.D(n_89),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_131),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_85),
.C(n_84),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_101),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_97),
.B1(n_84),
.B2(n_69),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_92),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_109),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_90),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_125),
.B(n_115),
.Y(n_142)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_94),
.B(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_149),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_133),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_109),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_141),
.A2(n_12),
.B(n_4),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_148),
.B1(n_133),
.B2(n_129),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_103),
.C(n_86),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_154),
.C(n_128),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_112),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_147),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_112),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_25),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_117),
.Y(n_158)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_84),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_155),
.B(n_0),
.Y(n_167)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_158),
.B(n_177),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_166),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_3),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_162),
.C(n_164),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_123),
.C(n_120),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_131),
.B1(n_130),
.B2(n_116),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_167),
.B1(n_155),
.B2(n_135),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_151),
.B(n_114),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_13),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_152),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_2),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_176),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

BUFx12_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_145),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_181),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_182),
.B(n_183),
.Y(n_202)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_164),
.B(n_151),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_193),
.C(n_195),
.Y(n_199)
);

OA21x2_ASAP7_75t_SL g185 ( 
.A1(n_174),
.A2(n_150),
.B(n_162),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_185),
.A2(n_187),
.B1(n_192),
.B2(n_194),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_144),
.B1(n_138),
.B2(n_137),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_190),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_168),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_142),
.B1(n_135),
.B2(n_154),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_143),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_165),
.C(n_177),
.Y(n_203)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_201),
.Y(n_213)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_204),
.C(n_208),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_158),
.C(n_173),
.Y(n_204)
);

BUFx12_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_173),
.B1(n_160),
.B2(n_176),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_210),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_178),
.C(n_4),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g218 ( 
.A(n_209),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_178),
.B(n_5),
.C(n_6),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_191),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_216),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_193),
.C(n_180),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_215),
.B(n_217),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_180),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_200),
.C(n_207),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_3),
.C(n_5),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_219),
.B(n_6),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_3),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_220),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_206),
.C(n_212),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_222),
.B(n_229),
.Y(n_235)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_226),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_209),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_228),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_197),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_201),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_230),
.B(n_224),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_230),
.A2(n_202),
.B(n_221),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_233),
.A2(n_225),
.B(n_205),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_222),
.B(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_236),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_205),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_237),
.B(n_7),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_242),
.A3(n_233),
.B1(n_8),
.B2(n_9),
.C1(n_11),
.C2(n_12),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_231),
.B(n_7),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_7),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_240),
.A2(n_235),
.B(n_234),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_243),
.B(n_244),
.Y(n_247)
);

NAND4xp25_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_246),
.C(n_9),
.D(n_11),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_238),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g249 ( 
.A(n_248),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_249),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_247),
.Y(n_251)
);


endmodule