module fake_aes_6559_n_27 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_27);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVx1_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_10), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_5), .Y(n_16) );
AND2x4_ASAP7_75t_L g17 ( .A(n_9), .B(n_0), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
BUFx2_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
AOI22xp33_ASAP7_75t_SL g20 ( .A1(n_19), .A2(n_16), .B1(n_14), .B2(n_15), .Y(n_20) );
NAND3xp33_ASAP7_75t_SL g21 ( .A(n_20), .B(n_18), .C(n_0), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
NAND2x1p5_ASAP7_75t_SL g23 ( .A(n_22), .B(n_1), .Y(n_23) );
AOI22x1_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_2), .B1(n_3), .B2(n_6), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
NOR4xp25_ASAP7_75t_SL g26 ( .A(n_25), .B(n_7), .C(n_11), .D(n_12), .Y(n_26) );
INVx1_ASAP7_75t_SL g27 ( .A(n_26), .Y(n_27) );
endmodule