module real_aes_2674_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_791, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_791;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_756;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g213 ( .A(n_0), .B(n_135), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_1), .B(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_2), .B(n_141), .Y(n_499) );
AOI222xp33_ASAP7_75t_SL g102 ( .A1(n_3), .A2(n_103), .B1(n_108), .B2(n_454), .C1(n_459), .C2(n_465), .Y(n_102) );
XNOR2xp5_ASAP7_75t_L g109 ( .A(n_3), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_4), .B(n_131), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_5), .B(n_141), .Y(n_154) );
INVx1_ASAP7_75t_L g128 ( .A(n_6), .Y(n_128) );
NAND2xp33_ASAP7_75t_SL g205 ( .A(n_7), .B(n_139), .Y(n_205) );
INVx1_ASAP7_75t_L g186 ( .A(n_8), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_9), .A2(n_42), .B1(n_470), .B2(n_471), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_9), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_10), .Y(n_106) );
AND2x2_ASAP7_75t_L g152 ( .A(n_11), .B(n_145), .Y(n_152) );
AND2x2_ASAP7_75t_L g531 ( .A(n_12), .B(n_179), .Y(n_531) );
AND2x2_ASAP7_75t_L g539 ( .A(n_13), .B(n_202), .Y(n_539) );
INVx2_ASAP7_75t_L g146 ( .A(n_14), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_15), .B(n_131), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g445 ( .A(n_16), .Y(n_445) );
AOI221x1_ASAP7_75t_L g199 ( .A1(n_17), .A2(n_123), .B1(n_200), .B2(n_202), .C(n_204), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_18), .B(n_141), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_19), .B(n_141), .Y(n_512) );
INVx1_ASAP7_75t_L g449 ( .A(n_20), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_21), .A2(n_90), .B1(n_141), .B2(n_187), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_22), .A2(n_123), .B(n_156), .Y(n_155) );
AOI221xp5_ASAP7_75t_SL g166 ( .A1(n_23), .A2(n_37), .B1(n_123), .B2(n_141), .C(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_24), .B(n_135), .Y(n_157) );
AOI22xp5_ASAP7_75t_SL g439 ( .A1(n_25), .A2(n_78), .B1(n_440), .B2(n_441), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_25), .Y(n_441) );
OR2x2_ASAP7_75t_L g147 ( .A(n_26), .B(n_89), .Y(n_147) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_26), .A2(n_89), .B(n_146), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_27), .B(n_131), .Y(n_178) );
INVxp67_ASAP7_75t_L g198 ( .A(n_28), .Y(n_198) );
AND2x2_ASAP7_75t_L g229 ( .A(n_29), .B(n_144), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_30), .A2(n_123), .B(n_212), .Y(n_211) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_31), .A2(n_202), .B(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_32), .B(n_131), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_33), .A2(n_123), .B(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_34), .B(n_131), .Y(n_498) );
AND2x2_ASAP7_75t_L g124 ( .A(n_35), .B(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g139 ( .A(n_35), .B(n_128), .Y(n_139) );
INVx1_ASAP7_75t_L g194 ( .A(n_35), .Y(n_194) );
OR2x6_ASAP7_75t_L g447 ( .A(n_36), .B(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_38), .B(n_141), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_39), .A2(n_82), .B1(n_123), .B2(n_192), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_40), .B(n_131), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_41), .B(n_141), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_42), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_43), .B(n_135), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_44), .A2(n_123), .B(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g216 ( .A(n_45), .B(n_144), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_46), .B(n_135), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_47), .B(n_144), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_48), .B(n_141), .Y(n_487) );
INVx1_ASAP7_75t_L g127 ( .A(n_49), .Y(n_127) );
INVx1_ASAP7_75t_L g137 ( .A(n_49), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_50), .B(n_131), .Y(n_537) );
AND2x2_ASAP7_75t_L g503 ( .A(n_51), .B(n_144), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_52), .B(n_141), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_53), .B(n_135), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_54), .B(n_135), .Y(n_497) );
AND2x2_ASAP7_75t_L g148 ( .A(n_55), .B(n_144), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_56), .B(n_141), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_57), .B(n_131), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_58), .B(n_141), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_59), .A2(n_123), .B(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_60), .B(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_SL g181 ( .A(n_61), .B(n_145), .Y(n_181) );
AND2x2_ASAP7_75t_L g518 ( .A(n_62), .B(n_145), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_63), .A2(n_123), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_64), .B(n_131), .Y(n_158) );
AND2x2_ASAP7_75t_SL g266 ( .A(n_65), .B(n_179), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_66), .B(n_135), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_67), .B(n_135), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_68), .A2(n_93), .B1(n_123), .B2(n_192), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_69), .B(n_131), .Y(n_515) );
INVx1_ASAP7_75t_L g125 ( .A(n_70), .Y(n_125) );
INVx1_ASAP7_75t_L g133 ( .A(n_70), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_71), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_72), .B(n_135), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_73), .A2(n_123), .B(n_507), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_74), .A2(n_123), .B(n_566), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_75), .Y(n_787) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_76), .A2(n_123), .B(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g500 ( .A(n_77), .B(n_145), .Y(n_500) );
INVx1_ASAP7_75t_L g440 ( .A(n_78), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_79), .B(n_144), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_80), .B(n_141), .Y(n_140) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_81), .A2(n_84), .B1(n_141), .B2(n_187), .Y(n_264) );
INVx1_ASAP7_75t_L g450 ( .A(n_83), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_85), .B(n_135), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_86), .B(n_135), .Y(n_169) );
AND2x2_ASAP7_75t_L g569 ( .A(n_87), .B(n_179), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g122 ( .A1(n_88), .A2(n_123), .B(n_129), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_91), .B(n_131), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_92), .A2(n_123), .B(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_94), .B(n_131), .Y(n_567) );
INVxp67_ASAP7_75t_L g201 ( .A(n_95), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_96), .B(n_141), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_97), .B(n_131), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_98), .A2(n_123), .B(n_176), .Y(n_175) );
BUFx2_ASAP7_75t_L g517 ( .A(n_99), .Y(n_517) );
BUFx2_ASAP7_75t_L g107 ( .A(n_100), .Y(n_107) );
BUFx2_ASAP7_75t_SL g458 ( .A(n_100), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_101), .A2(n_467), .B1(n_468), .B2(n_469), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_101), .Y(n_467) );
CKINVDCx9p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
OR2x2_ASAP7_75t_SL g104 ( .A(n_105), .B(n_107), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_105), .A2(n_442), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g464 ( .A(n_105), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_107), .B(n_464), .Y(n_463) );
OAI21xp5_ASAP7_75t_SL g108 ( .A1(n_109), .A2(n_442), .B(n_451), .Y(n_108) );
AOI22x1_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_112), .B1(n_438), .B2(n_439), .Y(n_110) );
INVx4_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_112), .B(n_780), .Y(n_779) );
OAI22xp5_ASAP7_75t_SL g784 ( .A1(n_112), .A2(n_477), .B1(n_479), .B2(n_785), .Y(n_784) );
AND2x4_ASAP7_75t_L g112 ( .A(n_113), .B(n_377), .Y(n_112) );
NOR3xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_270), .C(n_321), .Y(n_113) );
OAI211xp5_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_160), .B(n_217), .C(n_248), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_149), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_119), .B(n_222), .Y(n_385) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g230 ( .A(n_120), .B(n_151), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_120), .B(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g247 ( .A(n_120), .B(n_237), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_120), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g284 ( .A(n_120), .B(n_260), .Y(n_284) );
INVx2_ASAP7_75t_L g310 ( .A(n_120), .Y(n_310) );
AND2x4_ASAP7_75t_L g319 ( .A(n_120), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g424 ( .A(n_120), .B(n_291), .Y(n_424) );
AO21x2_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_143), .B(n_148), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_140), .Y(n_121) );
AND2x6_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
BUFx3_ASAP7_75t_L g191 ( .A(n_124), .Y(n_191) );
AND2x6_ASAP7_75t_L g135 ( .A(n_125), .B(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g196 ( .A(n_125), .Y(n_196) );
AND2x4_ASAP7_75t_L g192 ( .A(n_126), .B(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AND2x4_ASAP7_75t_L g131 ( .A(n_127), .B(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g189 ( .A(n_127), .Y(n_189) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_128), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_134), .B(n_138), .Y(n_129) );
AND2x4_ASAP7_75t_L g142 ( .A(n_132), .B(n_136), .Y(n_142) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_135), .B(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_138), .A2(n_157), .B(n_158), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_138), .A2(n_168), .B(n_169), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_138), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_138), .A2(n_213), .B(n_214), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_138), .A2(n_226), .B(n_227), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_138), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_138), .A2(n_497), .B(n_498), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_138), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_138), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_138), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_138), .A2(n_536), .B(n_537), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_138), .A2(n_567), .B(n_568), .Y(n_566) );
INVx5_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g141 ( .A(n_139), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g206 ( .A(n_142), .Y(n_206) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_143), .A2(n_223), .B(n_229), .Y(n_222) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_143), .A2(n_223), .B(n_229), .Y(n_237) );
AOI21x1_ASAP7_75t_L g524 ( .A1(n_143), .A2(n_525), .B(n_531), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_144), .Y(n_143) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_144), .A2(n_166), .B(n_170), .Y(n_165) );
AO21x2_ASAP7_75t_L g545 ( .A1(n_144), .A2(n_546), .B(n_547), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_144), .A2(n_564), .B(n_565), .Y(n_563) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_SL g145 ( .A(n_146), .B(n_147), .Y(n_145) );
AND2x4_ASAP7_75t_L g159 ( .A(n_146), .B(n_147), .Y(n_159) );
AND2x2_ASAP7_75t_L g308 ( .A(n_149), .B(n_309), .Y(n_308) );
OAI32xp33_ASAP7_75t_L g391 ( .A1(n_149), .A2(n_313), .A3(n_317), .B1(n_324), .B2(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_149), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g245 ( .A(n_150), .B(n_246), .Y(n_245) );
NAND3xp33_ASAP7_75t_L g318 ( .A(n_150), .B(n_240), .C(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g344 ( .A(n_150), .B(n_247), .Y(n_344) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_151), .Y(n_234) );
INVx5_ASAP7_75t_L g269 ( .A(n_151), .Y(n_269) );
AND2x4_ASAP7_75t_L g325 ( .A(n_151), .B(n_237), .Y(n_325) );
OR2x2_ASAP7_75t_L g340 ( .A(n_151), .B(n_260), .Y(n_340) );
OR2x2_ASAP7_75t_L g366 ( .A(n_151), .B(n_222), .Y(n_366) );
AND2x2_ASAP7_75t_L g374 ( .A(n_151), .B(n_320), .Y(n_374) );
AND2x4_ASAP7_75t_SL g399 ( .A(n_151), .B(n_319), .Y(n_399) );
OR2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_159), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_159), .B(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_159), .B(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_159), .B(n_201), .Y(n_200) );
NOR3xp33_ASAP7_75t_L g204 ( .A(n_159), .B(n_205), .C(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_159), .A2(n_487), .B(n_488), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_159), .A2(n_505), .B(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_161), .B(n_319), .Y(n_395) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_171), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_162), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OR2x6_ASAP7_75t_SL g219 ( .A(n_163), .B(n_220), .Y(n_219) );
INVxp67_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g244 ( .A(n_164), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_164), .B(n_279), .Y(n_297) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_164), .Y(n_435) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g252 ( .A(n_165), .Y(n_252) );
AND2x2_ASAP7_75t_L g277 ( .A(n_165), .B(n_208), .Y(n_277) );
INVx2_ASAP7_75t_L g305 ( .A(n_165), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_165), .B(n_172), .Y(n_346) );
BUFx3_ASAP7_75t_L g370 ( .A(n_165), .Y(n_370) );
OR2x2_ASAP7_75t_L g382 ( .A(n_165), .B(n_172), .Y(n_382) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_165), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_171), .A2(n_413), .B1(n_416), .B2(n_417), .Y(n_412) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_182), .Y(n_171) );
INVx1_ASAP7_75t_L g240 ( .A(n_172), .Y(n_240) );
OR2x2_ASAP7_75t_L g251 ( .A(n_172), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g258 ( .A(n_172), .Y(n_258) );
AND2x4_ASAP7_75t_SL g275 ( .A(n_172), .B(n_183), .Y(n_275) );
AND2x4_ASAP7_75t_L g280 ( .A(n_172), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g289 ( .A(n_172), .Y(n_289) );
OR2x2_ASAP7_75t_L g295 ( .A(n_172), .B(n_183), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_172), .B(n_297), .Y(n_296) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_172), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_172), .B(n_277), .Y(n_411) );
OR2x2_ASAP7_75t_L g427 ( .A(n_172), .B(n_330), .Y(n_427) );
OR2x6_ASAP7_75t_L g172 ( .A(n_173), .B(n_181), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_179), .Y(n_173) );
INVx2_ASAP7_75t_SL g262 ( .A(n_179), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_179), .A2(n_512), .B(n_513), .Y(n_511) );
BUFx4f_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx3_ASAP7_75t_L g203 ( .A(n_180), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_182), .B(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g253 ( .A(n_182), .Y(n_253) );
AND2x2_ASAP7_75t_SL g360 ( .A(n_182), .B(n_244), .Y(n_360) );
AND2x4_ASAP7_75t_L g182 ( .A(n_183), .B(n_207), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_183), .B(n_208), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_183), .B(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_183), .B(n_252), .Y(n_256) );
INVx3_ASAP7_75t_L g281 ( .A(n_183), .Y(n_281) );
INVx1_ASAP7_75t_L g314 ( .A(n_183), .Y(n_314) );
AND2x2_ASAP7_75t_L g394 ( .A(n_183), .B(n_258), .Y(n_394) );
AND2x4_ASAP7_75t_L g183 ( .A(n_184), .B(n_199), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_187), .B1(n_192), .B2(n_197), .Y(n_184) );
AND2x4_ASAP7_75t_L g187 ( .A(n_188), .B(n_191), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
NOR2x1p5_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx3_ASAP7_75t_L g493 ( .A(n_202), .Y(n_493) );
INVx4_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AOI21x1_ASAP7_75t_L g209 ( .A1(n_203), .A2(n_210), .B(n_216), .Y(n_209) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_203), .A2(n_533), .B(n_539), .Y(n_532) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_208), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g279 ( .A(n_208), .Y(n_279) );
AND2x2_ASAP7_75t_L g304 ( .A(n_208), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g330 ( .A(n_208), .B(n_252), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_208), .B(n_281), .Y(n_347) );
INVx1_ASAP7_75t_L g353 ( .A(n_208), .Y(n_353) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_215), .Y(n_210) );
AOI222xp33_ASAP7_75t_SL g217 ( .A1(n_218), .A2(n_221), .B1(n_231), .B2(n_238), .C1(n_241), .C2(n_245), .Y(n_217) );
CKINVDCx16_ASAP7_75t_R g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_230), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_222), .B(n_291), .Y(n_342) );
AND2x4_ASAP7_75t_L g358 ( .A(n_222), .B(n_269), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_228), .Y(n_223) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_233), .B(n_235), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g283 ( .A(n_234), .B(n_284), .Y(n_283) );
AOI222xp33_ASAP7_75t_L g248 ( .A1(n_235), .A2(n_249), .B1(n_254), .B2(n_259), .C1(n_267), .C2(n_791), .Y(n_248) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g387 ( .A(n_236), .B(n_291), .Y(n_387) );
OR2x2_ASAP7_75t_L g430 ( .A(n_236), .B(n_336), .Y(n_430) );
AND2x2_ASAP7_75t_L g259 ( .A(n_237), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g320 ( .A(n_237), .Y(n_320) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_237), .Y(n_335) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_238), .A2(n_349), .B(n_354), .C(n_355), .Y(n_348) );
INVx1_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g376 ( .A(n_240), .Y(n_376) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g306 ( .A(n_245), .Y(n_306) );
AND2x2_ASAP7_75t_L g290 ( .A(n_246), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g299 ( .A(n_246), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OAI31xp33_ASAP7_75t_L g341 ( .A1(n_249), .A2(n_267), .A3(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g343 ( .A1(n_250), .A2(n_300), .B(n_344), .C(n_345), .Y(n_343) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_253), .Y(n_250) );
OR2x2_ASAP7_75t_L g332 ( .A(n_251), .B(n_281), .Y(n_332) );
INVx2_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
BUFx2_ASAP7_75t_L g300 ( .A(n_260), .Y(n_300) );
AND2x2_ASAP7_75t_L g309 ( .A(n_260), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_261), .Y(n_291) );
AOI21x1_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_263), .B(n_266), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_269), .B(n_326), .Y(n_418) );
OAI211xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_282), .B(n_285), .C(n_307), .Y(n_270) );
INVxp33_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_273), .B(n_278), .Y(n_272) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g311 ( .A(n_275), .B(n_304), .Y(n_311) );
OR2x2_ASAP7_75t_L g287 ( .A(n_276), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g317 ( .A(n_276), .B(n_291), .Y(n_317) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g393 ( .A(n_277), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g416 ( .A(n_278), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_280), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_280), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g428 ( .A(n_280), .B(n_304), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_280), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g371 ( .A(n_281), .B(n_353), .Y(n_371) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
AOI322xp5_ASAP7_75t_L g425 ( .A1(n_284), .A2(n_304), .A3(n_358), .B1(n_383), .B2(n_426), .C1(n_428), .C2(n_429), .Y(n_425) );
AOI211xp5_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_290), .B(n_292), .C(n_301), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_288), .B(n_316), .Y(n_338) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g303 ( .A(n_289), .B(n_304), .Y(n_303) );
NOR2x1p5_ASAP7_75t_L g369 ( .A(n_289), .B(n_370), .Y(n_369) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_289), .Y(n_402) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_290), .A2(n_308), .B(n_311), .C(n_312), .Y(n_307) );
AND2x4_ASAP7_75t_L g326 ( .A(n_291), .B(n_310), .Y(n_326) );
INVx2_ASAP7_75t_L g336 ( .A(n_291), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_291), .B(n_325), .Y(n_356) );
AND2x2_ASAP7_75t_L g398 ( .A(n_291), .B(n_399), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_291), .B(n_415), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_291), .B(n_319), .Y(n_437) );
AOI21xp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_296), .B(n_298), .Y(n_292) );
AND2x2_ASAP7_75t_L g388 ( .A(n_294), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g316 ( .A(n_297), .Y(n_316) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_306), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_309), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g403 ( .A(n_309), .Y(n_403) );
O2A1O1Ixp33_ASAP7_75t_SL g312 ( .A1(n_313), .A2(n_315), .B(n_317), .C(n_318), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_316), .Y(n_400) );
INVx3_ASAP7_75t_SL g415 ( .A(n_319), .Y(n_415) );
NAND5xp2_ASAP7_75t_L g321 ( .A(n_322), .B(n_341), .C(n_348), .D(n_361), .E(n_372), .Y(n_321) );
AOI222xp33_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_327), .B1(n_331), .B2(n_333), .C1(n_337), .C2(n_339), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_324), .A2(n_405), .B1(n_409), .B2(n_410), .Y(n_404) );
INVx2_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g354 ( .A(n_325), .B(n_326), .Y(n_354) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_335), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_336), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g373 ( .A(n_336), .B(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g384 ( .A(n_336), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g414 ( .A(n_340), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g362 ( .A(n_347), .Y(n_362) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVxp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AOI21xp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B(n_359), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_358), .A2(n_362), .B1(n_363), .B2(n_367), .Y(n_361) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_358), .Y(n_409) );
INVx2_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g375 ( .A(n_360), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g380 ( .A(n_362), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVx1_ASAP7_75t_SL g408 ( .A(n_371), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
NOR3xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_396), .C(n_419), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_379), .B(n_395), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_383), .B1(n_386), .B2(n_388), .C(n_391), .Y(n_379) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g420 ( .A(n_382), .B(n_408), .Y(n_420) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
OAI321xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_400), .A3(n_401), .B1(n_403), .B2(n_404), .C(n_412), .Y(n_396) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_410), .A2(n_432), .B1(n_436), .B2(n_437), .Y(n_431) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI211xp5_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_421), .B(n_425), .C(n_431), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVxp33_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx2_ASAP7_75t_L g453 ( .A(n_444), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
OR2x6_ASAP7_75t_SL g477 ( .A(n_445), .B(n_446), .Y(n_477) );
AND2x6_ASAP7_75t_SL g782 ( .A(n_445), .B(n_447), .Y(n_782) );
OR2x2_ASAP7_75t_L g789 ( .A(n_445), .B(n_447), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g461 ( .A(n_453), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
CKINVDCx11_ASAP7_75t_R g456 ( .A(n_457), .Y(n_456) );
CKINVDCx8_ASAP7_75t_R g457 ( .A(n_458), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVxp67_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_472), .B(n_783), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_466), .A2(n_784), .B(n_786), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OAI21x1_ASAP7_75t_SL g473 ( .A1(n_474), .A2(n_478), .B(n_779), .Y(n_473) );
BUFx4f_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_476), .Y(n_475) );
CKINVDCx11_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
INVx4_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND3x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_657), .C(n_753), .Y(n_479) );
NOR3xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_599), .C(n_626), .Y(n_480) );
OAI211xp5_ASAP7_75t_SL g481 ( .A1(n_482), .A2(n_519), .B(n_548), .C(n_572), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_501), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g549 ( .A1(n_483), .A2(n_550), .B(n_554), .C(n_560), .Y(n_549) );
OR2x2_ASAP7_75t_L g672 ( .A(n_483), .B(n_609), .Y(n_672) );
INVx2_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g639 ( .A(n_484), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_484), .B(n_610), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_484), .B(n_755), .Y(n_770) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_492), .Y(n_484) );
AND2x2_ASAP7_75t_L g556 ( .A(n_485), .B(n_502), .Y(n_556) );
INVx1_ASAP7_75t_L g576 ( .A(n_485), .Y(n_576) );
OR2x2_ASAP7_75t_L g591 ( .A(n_485), .B(n_510), .Y(n_591) );
INVx2_ASAP7_75t_L g597 ( .A(n_485), .Y(n_597) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_485), .Y(n_652) );
INVx1_ASAP7_75t_L g729 ( .A(n_485), .Y(n_729) );
NOR2x1_ASAP7_75t_SL g578 ( .A(n_492), .B(n_510), .Y(n_578) );
AND2x2_ASAP7_75t_L g608 ( .A(n_492), .B(n_597), .Y(n_608) );
AO21x1_ASAP7_75t_SL g492 ( .A1(n_493), .A2(n_494), .B(n_500), .Y(n_492) );
AO21x2_ASAP7_75t_L g559 ( .A1(n_493), .A2(n_494), .B(n_500), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_499), .Y(n_494) );
OR2x2_ASAP7_75t_L g602 ( .A(n_501), .B(n_603), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_501), .B(n_709), .Y(n_708) );
INVx3_ASAP7_75t_L g730 ( .A(n_501), .Y(n_730) );
NAND2x1_ASAP7_75t_L g501 ( .A(n_502), .B(n_510), .Y(n_501) );
OR2x2_ASAP7_75t_SL g590 ( .A(n_502), .B(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g594 ( .A(n_502), .Y(n_594) );
INVx4_ASAP7_75t_L g610 ( .A(n_502), .Y(n_610) );
OR2x2_ASAP7_75t_L g625 ( .A(n_502), .B(n_558), .Y(n_625) );
AND2x2_ASAP7_75t_L g664 ( .A(n_502), .B(n_578), .Y(n_664) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_502), .Y(n_676) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
AND2x2_ASAP7_75t_L g557 ( .A(n_510), .B(n_558), .Y(n_557) );
OR2x2_ASAP7_75t_L g609 ( .A(n_510), .B(n_610), .Y(n_609) );
BUFx2_ASAP7_75t_L g624 ( .A(n_510), .Y(n_624) );
AND2x2_ASAP7_75t_L g640 ( .A(n_510), .B(n_610), .Y(n_640) );
AND2x2_ASAP7_75t_L g653 ( .A(n_510), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g685 ( .A(n_510), .B(n_597), .Y(n_685) );
INVx2_ASAP7_75t_SL g755 ( .A(n_510), .Y(n_755) );
OR2x6_ASAP7_75t_L g510 ( .A(n_511), .B(n_518), .Y(n_510) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NOR2xp67_ASAP7_75t_L g520 ( .A(n_521), .B(n_540), .Y(n_520) );
OAI211xp5_ASAP7_75t_L g626 ( .A1(n_521), .A2(n_627), .B(n_631), .C(n_647), .Y(n_626) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g722 ( .A(n_522), .B(n_561), .Y(n_722) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_532), .Y(n_522) );
INVx2_ASAP7_75t_L g571 ( .A(n_523), .Y(n_571) );
AND2x4_ASAP7_75t_SL g582 ( .A(n_523), .B(n_562), .Y(n_582) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_523), .Y(n_586) );
AND2x2_ASAP7_75t_L g644 ( .A(n_523), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g718 ( .A(n_523), .Y(n_718) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_524), .Y(n_620) );
AND2x2_ASAP7_75t_L g663 ( .A(n_524), .B(n_532), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_530), .Y(n_525) );
INVx2_ASAP7_75t_L g553 ( .A(n_532), .Y(n_553) );
AND2x2_ASAP7_75t_L g613 ( .A(n_532), .B(n_562), .Y(n_613) );
INVx2_ASAP7_75t_L g645 ( .A(n_532), .Y(n_645) );
OR2x2_ASAP7_75t_L g668 ( .A(n_532), .B(n_543), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_538), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_540), .B(n_585), .Y(n_692) );
AND2x2_ASAP7_75t_L g726 ( .A(n_540), .B(n_662), .Y(n_726) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OAI31xp33_ASAP7_75t_SL g647 ( .A1(n_541), .A2(n_628), .A3(n_648), .B(n_655), .Y(n_647) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_542), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx3_ASAP7_75t_L g581 ( .A(n_543), .Y(n_581) );
AND2x2_ASAP7_75t_L g598 ( .A(n_543), .B(n_561), .Y(n_598) );
AND2x4_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
AND2x4_ASAP7_75t_L g588 ( .A(n_544), .B(n_545), .Y(n_588) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g733 ( .A(n_551), .Y(n_733) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NOR2x1_ASAP7_75t_L g615 ( .A(n_553), .B(n_562), .Y(n_615) );
AND2x2_ASAP7_75t_L g656 ( .A(n_553), .B(n_571), .Y(n_656) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
AND2x2_ASAP7_75t_L g636 ( .A(n_557), .B(n_594), .Y(n_636) );
AND2x2_ASAP7_75t_L g595 ( .A(n_558), .B(n_596), .Y(n_595) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_558), .Y(n_604) );
INVx2_ASAP7_75t_L g654 ( .A(n_558), .Y(n_654) );
AND2x2_ASAP7_75t_L g744 ( .A(n_558), .B(n_729), .Y(n_744) );
INVx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g750 ( .A(n_560), .Y(n_750) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_561), .B(n_570), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_561), .B(n_620), .Y(n_689) );
AND2x2_ASAP7_75t_L g737 ( .A(n_561), .B(n_663), .Y(n_737) );
INVx4_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g646 ( .A(n_562), .B(n_618), .Y(n_646) );
AND2x2_ASAP7_75t_L g655 ( .A(n_562), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g667 ( .A(n_562), .Y(n_667) );
BUFx2_ASAP7_75t_L g683 ( .A(n_562), .Y(n_683) );
AND2x4_ASAP7_75t_L g717 ( .A(n_562), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g762 ( .A(n_562), .B(n_663), .Y(n_762) );
OR2x6_ASAP7_75t_L g562 ( .A(n_563), .B(n_569), .Y(n_562) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
AOI222xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_579), .B1(n_583), .B2(n_589), .C1(n_592), .C2(n_598), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_574), .A2(n_638), .B1(n_641), .B2(n_646), .Y(n_637) );
OR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
AND2x2_ASAP7_75t_L g621 ( .A(n_575), .B(n_622), .Y(n_621) );
AND2x4_ASAP7_75t_SL g635 ( .A(n_575), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_575), .B(n_640), .Y(n_773) );
INVx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g734 ( .A(n_576), .B(n_640), .Y(n_734) );
OR2x2_ASAP7_75t_L g711 ( .A(n_577), .B(n_593), .Y(n_711) );
OR2x2_ASAP7_75t_L g719 ( .A(n_577), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g703 ( .A(n_578), .B(n_596), .Y(n_703) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
OR2x2_ASAP7_75t_L g611 ( .A(n_581), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g761 ( .A(n_581), .B(n_762), .Y(n_761) );
AND2x2_ASAP7_75t_L g712 ( .A(n_582), .B(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_582), .B(n_741), .Y(n_740) );
INVx2_ASAP7_75t_SL g747 ( .A(n_582), .Y(n_747) );
INVxp67_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
INVx2_ASAP7_75t_L g732 ( .A(n_585), .Y(n_732) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g634 ( .A(n_586), .B(n_613), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_587), .B(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g633 ( .A(n_587), .Y(n_633) );
NOR2x1_ASAP7_75t_L g642 ( .A(n_587), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g736 ( .A(n_587), .B(n_608), .Y(n_736) );
INVx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g670 ( .A(n_588), .B(n_656), .Y(n_670) );
AND2x2_ASAP7_75t_L g713 ( .A(n_588), .B(n_645), .Y(n_713) );
AND2x4_ASAP7_75t_L g628 ( .A(n_589), .B(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g769 ( .A(n_591), .B(n_625), .Y(n_769) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_593), .B(n_608), .Y(n_752) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_594), .B(n_608), .Y(n_674) );
A2O1A1Ixp33_ASAP7_75t_L g735 ( .A1(n_594), .A2(n_635), .B(n_736), .C(n_737), .Y(n_735) );
AND2x2_ASAP7_75t_L g766 ( .A(n_594), .B(n_744), .Y(n_766) );
INVx1_ASAP7_75t_L g677 ( .A(n_595), .Y(n_677) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_598), .B(n_662), .Y(n_661) );
OAI21xp33_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_611), .B(n_614), .Y(n_599) );
NOR2x1_ASAP7_75t_L g600 ( .A(n_601), .B(n_605), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_602), .A2(n_755), .B1(n_756), .B2(n_758), .Y(n_754) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g630 ( .A(n_604), .Y(n_630) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NOR2xp67_ASAP7_75t_L g651 ( .A(n_610), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g702 ( .A(n_610), .Y(n_702) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI21xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_616), .B(n_621), .Y(n_614) );
INVx1_ASAP7_75t_L g693 ( .A(n_615), .Y(n_693) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx2_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_635), .B(n_637), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
OR2x2_ASAP7_75t_L g678 ( .A(n_633), .B(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g715 ( .A(n_633), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_633), .B(n_663), .Y(n_751) );
INVx1_ASAP7_75t_L g771 ( .A(n_634), .Y(n_771) );
AOI221xp5_ASAP7_75t_L g738 ( .A1(n_636), .A2(n_739), .B1(n_742), .B2(n_745), .C(n_748), .Y(n_738) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI321xp33_ASAP7_75t_L g759 ( .A1(n_641), .A2(n_676), .A3(n_760), .B1(n_763), .B2(n_765), .C(n_767), .Y(n_759) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g700 ( .A(n_645), .Y(n_700) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g694 ( .A(n_650), .Y(n_694) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g720 ( .A(n_651), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_653), .A2(n_681), .B1(n_685), .B2(n_686), .C(n_691), .Y(n_680) );
INVxp67_ASAP7_75t_L g709 ( .A(n_654), .Y(n_709) );
INVx1_ASAP7_75t_L g679 ( .A(n_656), .Y(n_679) );
NOR2xp67_ASAP7_75t_L g657 ( .A(n_658), .B(n_704), .Y(n_657) );
NAND3xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_680), .C(n_695), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_664), .B1(n_665), .B2(n_671), .C(n_673), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g778 ( .A(n_663), .Y(n_778) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_666), .B(n_669), .Y(n_665) );
OR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g758 ( .A(n_667), .B(n_713), .Y(n_758) );
INVx2_ASAP7_75t_SL g690 ( .A(n_668), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_669), .A2(n_674), .B1(n_675), .B2(n_678), .Y(n_673) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_677), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_678), .B(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g684 ( .A(n_679), .Y(n_684) );
AOI222xp33_ASAP7_75t_L g723 ( .A1(n_681), .A2(n_724), .B1(n_726), .B2(n_727), .C1(n_731), .C2(n_734), .Y(n_723) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_682), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g757 ( .A(n_682), .B(n_736), .Y(n_757) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_690), .B(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_690), .B(n_750), .Y(n_749) );
AOI21xp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B(n_694), .Y(n_691) );
NAND2xp33_ASAP7_75t_SL g695 ( .A(n_696), .B(n_701), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
BUFx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_701), .B(n_776), .Y(n_775) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
NAND4xp25_ASAP7_75t_SL g704 ( .A(n_705), .B(n_723), .C(n_735), .D(n_738), .Y(n_704) );
O2A1O1Ixp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_710), .B(n_712), .C(n_714), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_711), .A2(n_715), .B1(n_719), .B2(n_721), .Y(n_714) );
INVx1_ASAP7_75t_L g741 ( .A(n_713), .Y(n_741) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_730), .Y(n_727) );
BUFx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_730), .B(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVxp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVxp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_747), .A2(n_769), .B1(n_770), .B2(n_771), .Y(n_768) );
AOI21xp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_751), .B(n_752), .Y(n_748) );
NOR4xp25_ASAP7_75t_L g753 ( .A(n_754), .B(n_759), .C(n_772), .D(n_774), .Y(n_753) );
INVxp67_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx3_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
CKINVDCx11_ASAP7_75t_R g785 ( .A(n_782), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
BUFx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
endmodule