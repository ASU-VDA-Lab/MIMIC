module real_jpeg_26408_n_6 (n_5, n_4, n_39, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_39;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_1),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_2),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_3),
.B(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

OR2x2_ASAP7_75t_SL g29 ( 
.A(n_3),
.B(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_3),
.B(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_3),
.B(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_4),
.A2(n_15),
.B(n_20),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_5),
.B(n_9),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_9),
.Y(n_11)
);

AOI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_13),
.B(n_21),
.C(n_31),
.Y(n_6)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_L g21 ( 
.A1(n_10),
.A2(n_15),
.B1(n_22),
.B2(n_27),
.Y(n_21)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_18),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_11),
.A2(n_18),
.B1(n_23),
.B2(n_24),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_12),
.B(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_17),
.Y(n_16)
);

OAI322xp33_ASAP7_75t_L g31 ( 
.A1(n_17),
.A2(n_19),
.A3(n_26),
.B1(n_30),
.B2(n_32),
.C1(n_33),
.C2(n_39),
.Y(n_31)
);

AOI211xp5_ASAP7_75t_SL g33 ( 
.A1(n_18),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);


endmodule