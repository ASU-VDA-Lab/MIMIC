module fake_jpeg_17034_n_243 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_243);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_243;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_32),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_32),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_0),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_16),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_42),
.B(n_22),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_20),
.B1(n_26),
.B2(n_22),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_50),
.B1(n_17),
.B2(n_21),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_23),
.B1(n_31),
.B2(n_20),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_16),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_26),
.Y(n_52)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_31),
.B1(n_20),
.B2(n_26),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_58),
.B1(n_35),
.B2(n_21),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_33),
.B(n_21),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_31),
.B1(n_16),
.B2(n_17),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_25),
.Y(n_62)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_63),
.B(n_67),
.Y(n_116)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_25),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_69),
.A2(n_82),
.B1(n_85),
.B2(n_47),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_34),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_30),
.C(n_27),
.Y(n_118)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_19),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_72),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_87),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_77),
.B1(n_41),
.B2(n_37),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_50),
.Y(n_76)
);

NOR2xp67_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_83),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_35),
.B1(n_38),
.B2(n_34),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_78),
.A2(n_27),
.B1(n_18),
.B2(n_2),
.Y(n_120)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_45),
.B(n_24),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_28),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_94),
.B1(n_19),
.B2(n_24),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_47),
.A2(n_17),
.B1(n_22),
.B2(n_19),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_89),
.A2(n_24),
.B1(n_28),
.B2(n_38),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_35),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_92),
.Y(n_113)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_41),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g135 ( 
.A(n_97),
.B(n_99),
.C(n_103),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_39),
.B1(n_41),
.B2(n_37),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_102),
.A2(n_107),
.B1(n_108),
.B2(n_85),
.Y(n_145)
);

AOI32xp33_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_37),
.A3(n_39),
.B1(n_41),
.B2(n_38),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_106),
.B(n_93),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_37),
.B1(n_28),
.B2(n_30),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_32),
.B1(n_30),
.B2(n_27),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_79),
.A2(n_30),
.B1(n_27),
.B2(n_18),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_92),
.B(n_61),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_118),
.B(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_89),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_121),
.A2(n_125),
.B1(n_136),
.B2(n_145),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_122),
.B(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_128),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_65),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_80),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_61),
.Y(n_128)
);

XOR2x1_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_94),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_116),
.B(n_112),
.Y(n_148)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_132),
.B(n_137),
.Y(n_150)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_81),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_141),
.Y(n_156)
);

AOI22x1_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_93),
.B1(n_94),
.B2(n_65),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_65),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_99),
.Y(n_157)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_140),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_64),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_100),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_110),
.Y(n_168)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_144),
.B(n_108),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_144),
.A2(n_97),
.B1(n_98),
.B2(n_118),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_147),
.A2(n_136),
.B1(n_138),
.B2(n_145),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_122),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_112),
.B(n_100),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_131),
.B(n_123),
.Y(n_177)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_112),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_87),
.Y(n_159)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_114),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_166),
.Y(n_183)
);

AO221x1_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_66),
.B1(n_71),
.B2(n_119),
.C(n_110),
.Y(n_162)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_139),
.B(n_119),
.Y(n_166)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_184),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_171),
.Y(n_200)
);

NOR3xp33_ASAP7_75t_SL g171 ( 
.A(n_150),
.B(n_129),
.C(n_135),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_146),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_161),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_163),
.A2(n_131),
.B1(n_135),
.B2(n_132),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_176),
.A2(n_158),
.B1(n_163),
.B2(n_148),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_177),
.A2(n_179),
.B(n_160),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_143),
.B(n_137),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_156),
.B(n_84),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_74),
.Y(n_182)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_74),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_154),
.C(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_188),
.A2(n_0),
.B(n_1),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_190),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_159),
.C(n_158),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_193),
.C(n_201),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_155),
.C(n_157),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_165),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_174),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_153),
.B1(n_167),
.B2(n_164),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_198),
.B1(n_60),
.B2(n_91),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_173),
.A2(n_183),
.B1(n_178),
.B2(n_175),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_166),
.C(n_161),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_202),
.B(n_208),
.Y(n_222)
);

AOI321xp33_ASAP7_75t_L g204 ( 
.A1(n_189),
.A2(n_171),
.A3(n_176),
.B1(n_169),
.B2(n_179),
.C(n_178),
.Y(n_204)
);

AOI321xp33_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_206),
.A3(n_213),
.B1(n_203),
.B2(n_6),
.C(n_7),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_201),
.A2(n_183),
.B1(n_177),
.B2(n_167),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_207),
.B1(n_211),
.B2(n_212),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_200),
.A2(n_164),
.B1(n_146),
.B2(n_162),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_15),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_192),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_214),
.C(n_210),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_191),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_193),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_60),
.C(n_15),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_219),
.C(n_220),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_223),
.B(n_8),
.Y(n_229)
);

INVxp33_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_204),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_209),
.C(n_205),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_190),
.C(n_199),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_0),
.C(n_1),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_3),
.C(n_6),
.Y(n_227)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_218),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_227),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_7),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_9),
.Y(n_231)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_217),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_231),
.B(n_232),
.Y(n_237)
);

NOR2xp67_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_215),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_225),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_235),
.A2(n_236),
.B(n_10),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_9),
.C(n_10),
.Y(n_236)
);

AOI321xp33_ASAP7_75t_L g238 ( 
.A1(n_237),
.A2(n_231),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_238),
.A2(n_239),
.B(n_14),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_241),
.B(n_11),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_238),
.B(n_11),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_12),
.Y(n_243)
);


endmodule