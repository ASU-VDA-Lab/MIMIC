module real_aes_119_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_0), .B(n_504), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_1), .A2(n_506), .B(n_507), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_2), .B(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_3), .B(n_182), .Y(n_540) );
INVx1_ASAP7_75t_L g137 ( .A(n_4), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_5), .B(n_146), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_6), .B(n_182), .Y(n_528) );
INVx1_ASAP7_75t_L g192 ( .A(n_7), .Y(n_192) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_8), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_9), .Y(n_208) );
NAND2xp33_ASAP7_75t_L g561 ( .A(n_10), .B(n_179), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_11), .A2(n_494), .B1(n_821), .B2(n_822), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_11), .Y(n_821) );
INVx2_ASAP7_75t_L g145 ( .A(n_12), .Y(n_145) );
AOI221x1_ASAP7_75t_L g585 ( .A1(n_13), .A2(n_26), .B1(n_504), .B2(n_506), .C(n_586), .Y(n_585) );
AND3x1_ASAP7_75t_L g108 ( .A(n_14), .B(n_40), .C(n_109), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_14), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_15), .B(n_504), .Y(n_557) );
INVx1_ASAP7_75t_L g180 ( .A(n_16), .Y(n_180) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_17), .A2(n_168), .B(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_18), .B(n_222), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_19), .B(n_182), .Y(n_517) );
AO21x1_ASAP7_75t_L g535 ( .A1(n_20), .A2(n_504), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g106 ( .A(n_21), .Y(n_106) );
AOI221xp5_ASAP7_75t_L g114 ( .A1(n_22), .A2(n_115), .B1(n_795), .B2(n_796), .C(n_800), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g795 ( .A(n_22), .Y(n_795) );
INVx1_ASAP7_75t_L g177 ( .A(n_23), .Y(n_177) );
INVx1_ASAP7_75t_SL g252 ( .A(n_24), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_25), .B(n_157), .Y(n_156) );
AOI33xp33_ASAP7_75t_L g229 ( .A1(n_27), .A2(n_54), .A3(n_134), .B1(n_152), .B2(n_230), .B3(n_231), .Y(n_229) );
NAND2x1_ASAP7_75t_L g578 ( .A(n_28), .B(n_182), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_29), .Y(n_801) );
NAND2x1_ASAP7_75t_L g527 ( .A(n_30), .B(n_179), .Y(n_527) );
INVx1_ASAP7_75t_L g201 ( .A(n_31), .Y(n_201) );
OA21x2_ASAP7_75t_L g144 ( .A1(n_32), .A2(n_86), .B(n_145), .Y(n_144) );
OR2x2_ASAP7_75t_L g147 ( .A(n_32), .B(n_86), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_33), .B(n_190), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_34), .B(n_179), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_35), .B(n_182), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_36), .B(n_179), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_37), .Y(n_807) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_38), .A2(n_506), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g140 ( .A(n_39), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g151 ( .A(n_39), .Y(n_151) );
AND2x2_ASAP7_75t_L g166 ( .A(n_39), .B(n_137), .Y(n_166) );
OR2x6_ASAP7_75t_L g121 ( .A(n_40), .B(n_105), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_41), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_42), .B(n_504), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_43), .B(n_190), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_44), .A2(n_131), .B1(n_143), .B2(n_146), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_45), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_46), .B(n_157), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_47), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_48), .B(n_179), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_49), .B(n_168), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_50), .B(n_157), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_51), .A2(n_506), .B(n_526), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_52), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_53), .B(n_179), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_55), .B(n_157), .Y(n_220) );
INVx1_ASAP7_75t_L g135 ( .A(n_56), .Y(n_135) );
INVx1_ASAP7_75t_L g159 ( .A(n_56), .Y(n_159) );
AND2x2_ASAP7_75t_L g221 ( .A(n_57), .B(n_222), .Y(n_221) );
AOI221xp5_ASAP7_75t_L g189 ( .A1(n_58), .A2(n_75), .B1(n_149), .B2(n_190), .C(n_191), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_59), .B(n_190), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_60), .B(n_182), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_61), .B(n_143), .Y(n_210) );
AOI21xp5_ASAP7_75t_SL g240 ( .A1(n_62), .A2(n_149), .B(n_241), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_63), .A2(n_506), .B(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_64), .A2(n_100), .B1(n_112), .B2(n_823), .Y(n_99) );
INVx1_ASAP7_75t_L g173 ( .A(n_65), .Y(n_173) );
AO21x1_ASAP7_75t_L g537 ( .A1(n_66), .A2(n_506), .B(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_67), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g219 ( .A(n_68), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_69), .B(n_504), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_70), .A2(n_149), .B(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g551 ( .A(n_71), .B(n_223), .Y(n_551) );
INVx1_ASAP7_75t_L g141 ( .A(n_72), .Y(n_141) );
INVx1_ASAP7_75t_L g161 ( .A(n_72), .Y(n_161) );
AND2x2_ASAP7_75t_L g530 ( .A(n_73), .B(n_197), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_74), .B(n_190), .Y(n_232) );
AND2x2_ASAP7_75t_L g254 ( .A(n_76), .B(n_197), .Y(n_254) );
INVx1_ASAP7_75t_L g174 ( .A(n_77), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_78), .A2(n_149), .B(n_251), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g148 ( .A1(n_79), .A2(n_149), .B(n_155), .C(n_167), .Y(n_148) );
INVx1_ASAP7_75t_L g107 ( .A(n_80), .Y(n_107) );
AND2x2_ASAP7_75t_L g501 ( .A(n_81), .B(n_197), .Y(n_501) );
AND2x2_ASAP7_75t_SL g238 ( .A(n_82), .B(n_197), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_83), .B(n_504), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_84), .A2(n_149), .B1(n_227), .B2(n_228), .Y(n_226) );
AND2x2_ASAP7_75t_L g536 ( .A(n_85), .B(n_146), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_87), .B(n_179), .Y(n_518) );
AND2x2_ASAP7_75t_L g581 ( .A(n_88), .B(n_197), .Y(n_581) );
INVx1_ASAP7_75t_L g242 ( .A(n_89), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_90), .B(n_182), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_91), .A2(n_506), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_92), .B(n_179), .Y(n_587) );
AND2x2_ASAP7_75t_L g233 ( .A(n_93), .B(n_197), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_94), .B(n_182), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_95), .A2(n_199), .B(n_200), .C(n_202), .Y(n_198) );
BUFx2_ASAP7_75t_SL g817 ( .A(n_96), .Y(n_817) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_97), .A2(n_506), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_98), .B(n_157), .Y(n_243) );
BUFx4f_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_102), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_SL g103 ( .A(n_104), .B(n_108), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AO21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_813), .B(n_818), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g113 ( .A(n_114), .B(n_805), .Y(n_113) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_122), .B1(n_494), .B2(n_793), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_117), .A2(n_122), .B1(n_494), .B2(n_798), .Y(n_797) );
CKINVDCx11_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
OR2x6_ASAP7_75t_SL g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AND2x6_ASAP7_75t_SL g794 ( .A(n_119), .B(n_121), .Y(n_794) );
OR2x2_ASAP7_75t_L g804 ( .A(n_119), .B(n_121), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_119), .B(n_120), .Y(n_812) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_428), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_351), .Y(n_123) );
NAND3xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_298), .C(n_331), .Y(n_124) );
AOI211xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_255), .B(n_264), .C(n_288), .Y(n_125) );
OAI21xp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_184), .B(n_234), .Y(n_126) );
OR2x2_ASAP7_75t_L g308 ( .A(n_127), .B(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g463 ( .A(n_127), .B(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AOI22xp33_ASAP7_75t_SL g353 ( .A1(n_128), .A2(n_354), .B1(n_358), .B2(n_360), .Y(n_353) );
AND2x2_ASAP7_75t_L g390 ( .A(n_128), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_169), .Y(n_128) );
INVx1_ASAP7_75t_L g287 ( .A(n_129), .Y(n_287) );
AND2x4_ASAP7_75t_L g304 ( .A(n_129), .B(n_285), .Y(n_304) );
INVx2_ASAP7_75t_L g326 ( .A(n_129), .Y(n_326) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_129), .Y(n_409) );
AND2x2_ASAP7_75t_L g480 ( .A(n_129), .B(n_237), .Y(n_480) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_148), .Y(n_129) );
NOR3xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_138), .C(n_142), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g190 ( .A(n_133), .B(n_139), .Y(n_190) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
OR2x6_ASAP7_75t_L g164 ( .A(n_134), .B(n_153), .Y(n_164) );
INVxp33_ASAP7_75t_L g230 ( .A(n_134), .Y(n_230) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g154 ( .A(n_135), .B(n_137), .Y(n_154) );
AND2x4_ASAP7_75t_L g182 ( .A(n_135), .B(n_160), .Y(n_182) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x6_ASAP7_75t_L g506 ( .A(n_140), .B(n_154), .Y(n_506) );
INVx2_ASAP7_75t_L g153 ( .A(n_141), .Y(n_153) );
AND2x6_ASAP7_75t_L g179 ( .A(n_141), .B(n_158), .Y(n_179) );
INVx4_ASAP7_75t_L g197 ( .A(n_143), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_143), .B(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx4f_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
AND2x4_ASAP7_75t_L g146 ( .A(n_145), .B(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_SL g223 ( .A(n_145), .B(n_147), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_146), .B(n_165), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_146), .A2(n_240), .B(n_244), .Y(n_239) );
INVx1_ASAP7_75t_SL g513 ( .A(n_146), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_146), .B(n_542), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_146), .A2(n_557), .B(n_558), .Y(n_556) );
INVxp67_ASAP7_75t_L g209 ( .A(n_149), .Y(n_209) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_154), .Y(n_149) );
NOR2x1p5_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
INVx1_ASAP7_75t_L g231 ( .A(n_152), .Y(n_231) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_162), .B(n_165), .Y(n_155) );
INVx1_ASAP7_75t_L g175 ( .A(n_157), .Y(n_175) );
AND2x4_ASAP7_75t_L g504 ( .A(n_157), .B(n_166), .Y(n_504) );
AND2x4_ASAP7_75t_L g157 ( .A(n_158), .B(n_160), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_164), .A2(n_173), .B1(n_174), .B2(n_175), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_SL g191 ( .A1(n_164), .A2(n_165), .B(n_192), .C(n_193), .Y(n_191) );
INVxp67_ASAP7_75t_L g199 ( .A(n_164), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_164), .A2(n_165), .B(n_219), .C(n_220), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_164), .A2(n_165), .B(n_242), .C(n_243), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_SL g251 ( .A1(n_164), .A2(n_165), .B(n_252), .C(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g227 ( .A(n_165), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_165), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_165), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_165), .A2(n_527), .B(n_528), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_165), .A2(n_539), .B(n_540), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_165), .A2(n_548), .B(n_549), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_165), .A2(n_560), .B(n_561), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_165), .A2(n_578), .B(n_579), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_165), .A2(n_587), .B(n_588), .Y(n_586) );
INVx5_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_166), .Y(n_202) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_167), .A2(n_225), .B(n_233), .Y(n_224) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_167), .A2(n_225), .B(n_233), .Y(n_269) );
INVx2_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_168), .A2(n_189), .B(n_194), .Y(n_188) );
AND2x2_ASAP7_75t_L g245 ( .A(n_169), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g274 ( .A(n_169), .Y(n_274) );
INVx3_ASAP7_75t_L g285 ( .A(n_169), .Y(n_285) );
AND2x4_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_176), .B(n_183), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_175), .B(n_201), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B1(n_180), .B2(n_181), .Y(n_176) );
INVxp67_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVxp67_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_184), .A2(n_475), .B1(n_477), .B2(n_479), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_184), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_212), .Y(n_185) );
INVx3_ASAP7_75t_L g258 ( .A(n_186), .Y(n_258) );
AND2x2_ASAP7_75t_L g266 ( .A(n_186), .B(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_186), .Y(n_296) );
NAND2x1_ASAP7_75t_SL g490 ( .A(n_186), .B(n_257), .Y(n_490) );
AND2x4_ASAP7_75t_L g186 ( .A(n_187), .B(n_195), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g263 ( .A(n_188), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_188), .B(n_269), .Y(n_281) );
AND2x2_ASAP7_75t_L g294 ( .A(n_188), .B(n_195), .Y(n_294) );
AND2x4_ASAP7_75t_L g301 ( .A(n_188), .B(n_302), .Y(n_301) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_188), .Y(n_350) );
INVxp67_ASAP7_75t_L g357 ( .A(n_188), .Y(n_357) );
INVx1_ASAP7_75t_L g362 ( .A(n_188), .Y(n_362) );
INVx1_ASAP7_75t_L g211 ( .A(n_190), .Y(n_211) );
INVx1_ASAP7_75t_L g261 ( .A(n_195), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_195), .B(n_271), .Y(n_280) );
INVx2_ASAP7_75t_L g348 ( .A(n_195), .Y(n_348) );
INVx1_ASAP7_75t_L g387 ( .A(n_195), .Y(n_387) );
OR2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_205), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B1(n_203), .B2(n_204), .Y(n_196) );
INVx3_ASAP7_75t_L g204 ( .A(n_197), .Y(n_204) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_204), .A2(n_215), .B(n_221), .Y(n_214) );
AO21x2_ASAP7_75t_L g271 ( .A1(n_204), .A2(n_215), .B(n_221), .Y(n_271) );
AO21x2_ASAP7_75t_L g544 ( .A1(n_204), .A2(n_545), .B(n_551), .Y(n_544) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_204), .A2(n_545), .B(n_551), .Y(n_566) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_204), .A2(n_575), .B(n_581), .Y(n_574) );
AO21x2_ASAP7_75t_L g599 ( .A1(n_204), .A2(n_575), .B(n_581), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_209), .B1(n_210), .B2(n_211), .Y(n_205) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g317 ( .A(n_212), .B(n_294), .Y(n_317) );
AND2x2_ASAP7_75t_L g385 ( .A(n_212), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g399 ( .A(n_212), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_212), .B(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_224), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NOR2x1_ASAP7_75t_L g262 ( .A(n_214), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g355 ( .A(n_214), .B(n_348), .Y(n_355) );
AND2x2_ASAP7_75t_L g446 ( .A(n_214), .B(n_268), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_222), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_222), .A2(n_503), .B(n_505), .Y(n_502) );
OA21x2_ASAP7_75t_L g584 ( .A1(n_222), .A2(n_585), .B(n_589), .Y(n_584) );
OA21x2_ASAP7_75t_L g629 ( .A1(n_222), .A2(n_585), .B(n_589), .Y(n_629) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g257 ( .A(n_224), .Y(n_257) );
INVx2_ASAP7_75t_L g302 ( .A(n_224), .Y(n_302) );
AND2x2_ASAP7_75t_L g347 ( .A(n_224), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_226), .B(n_232), .Y(n_225) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_245), .Y(n_235) );
AND2x2_ASAP7_75t_L g389 ( .A(n_236), .B(n_390), .Y(n_389) );
OR2x6_ASAP7_75t_L g448 ( .A(n_236), .B(n_449), .Y(n_448) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx4_ASAP7_75t_L g278 ( .A(n_237), .Y(n_278) );
AND2x4_ASAP7_75t_L g286 ( .A(n_237), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g321 ( .A(n_237), .B(n_246), .Y(n_321) );
INVx2_ASAP7_75t_L g370 ( .A(n_237), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_237), .B(n_344), .Y(n_419) );
AND2x2_ASAP7_75t_L g456 ( .A(n_237), .B(n_274), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_237), .B(n_339), .Y(n_464) );
OR2x6_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AND2x2_ASAP7_75t_L g297 ( .A(n_245), .B(n_286), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_245), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_SL g436 ( .A(n_245), .B(n_324), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_245), .B(n_337), .Y(n_458) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_246), .Y(n_276) );
AND2x2_ASAP7_75t_L g284 ( .A(n_246), .B(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_246), .Y(n_307) );
INVx2_ASAP7_75t_L g310 ( .A(n_246), .Y(n_310) );
INVx1_ASAP7_75t_L g343 ( .A(n_246), .Y(n_343) );
INVx1_ASAP7_75t_L g391 ( .A(n_246), .Y(n_391) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B(n_254), .Y(n_246) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_247), .A2(n_524), .B(n_530), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
NAND2xp33_ASAP7_75t_L g255 ( .A(n_256), .B(n_259), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_257), .B(n_260), .Y(n_333) );
OR2x2_ASAP7_75t_L g405 ( .A(n_257), .B(n_406), .Y(n_405) );
AND4x1_ASAP7_75t_SL g451 ( .A(n_257), .B(n_433), .C(n_452), .D(n_453), .Y(n_451) );
OR2x2_ASAP7_75t_L g475 ( .A(n_258), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
AND2x2_ASAP7_75t_L g312 ( .A(n_261), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_261), .B(n_270), .Y(n_462) );
AND2x2_ASAP7_75t_L g487 ( .A(n_262), .B(n_347), .Y(n_487) );
OAI32xp33_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_272), .A3(n_277), .B1(n_279), .B2(n_282), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g360 ( .A(n_267), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g460 ( .A(n_267), .B(n_414), .Y(n_460) );
AND2x4_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
AND2x2_ASAP7_75t_L g356 ( .A(n_268), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g442 ( .A(n_268), .Y(n_442) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_269), .B(n_271), .Y(n_476) );
INVx3_ASAP7_75t_L g293 ( .A(n_270), .Y(n_293) );
NAND2x1p5_ASAP7_75t_L g471 ( .A(n_270), .B(n_398), .Y(n_471) );
INVx3_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_271), .Y(n_330) );
AND2x2_ASAP7_75t_L g349 ( .A(n_271), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g483 ( .A(n_273), .Y(n_483) );
NAND2x1_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g323 ( .A(n_274), .Y(n_323) );
NOR2x1_ASAP7_75t_L g424 ( .A(n_274), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_277), .B(n_383), .Y(n_382) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g315 ( .A(n_278), .B(n_283), .Y(n_315) );
AND2x4_ASAP7_75t_L g337 ( .A(n_278), .B(n_287), .Y(n_337) );
AND2x4_ASAP7_75t_SL g408 ( .A(n_278), .B(n_409), .Y(n_408) );
NOR2x1_ASAP7_75t_L g434 ( .A(n_278), .B(n_359), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_279), .A2(n_402), .B1(n_405), .B2(n_407), .Y(n_401) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx2_ASAP7_75t_SL g421 ( .A(n_280), .Y(n_421) );
INVx2_ASAP7_75t_L g313 ( .A(n_281), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_284), .B(n_290), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_284), .A2(n_420), .B1(n_423), .B2(n_426), .Y(n_422) );
INVx1_ASAP7_75t_L g344 ( .A(n_285), .Y(n_344) );
AND2x2_ASAP7_75t_L g367 ( .A(n_285), .B(n_326), .Y(n_367) );
INVx2_ASAP7_75t_L g290 ( .A(n_286), .Y(n_290) );
OAI21xp5_ASAP7_75t_SL g288 ( .A1(n_289), .A2(n_291), .B(n_295), .Y(n_288) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_292), .A2(n_364), .B1(n_368), .B2(n_369), .Y(n_363) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_293), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_293), .B(n_361), .Y(n_377) );
INVx1_ASAP7_75t_L g381 ( .A(n_293), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
NOR3xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_314), .C(n_318), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_303), .B1(n_308), .B2(n_311), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g328 ( .A(n_301), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g368 ( .A(n_301), .B(n_355), .Y(n_368) );
AND2x2_ASAP7_75t_L g420 ( .A(n_301), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g437 ( .A(n_301), .B(n_387), .Y(n_437) );
AND2x2_ASAP7_75t_L g492 ( .A(n_301), .B(n_386), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx4_ASAP7_75t_L g359 ( .A(n_304), .Y(n_359) );
AND2x2_ASAP7_75t_L g369 ( .A(n_304), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_L g374 ( .A(n_307), .Y(n_374) );
AND2x2_ASAP7_75t_L g383 ( .A(n_307), .B(n_367), .Y(n_383) );
INVx1_ASAP7_75t_L g418 ( .A(n_309), .Y(n_418) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g339 ( .A(n_310), .Y(n_339) );
INVxp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_312), .B(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_313), .B(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_322), .B(n_327), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_320), .B(n_359), .Y(n_468) );
INVx2_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AOI21xp33_ASAP7_75t_SL g331 ( .A1(n_323), .A2(n_332), .B(n_334), .Y(n_331) );
AND2x2_ASAP7_75t_L g478 ( .A(n_323), .B(n_337), .Y(n_478) );
AND2x4_ASAP7_75t_L g341 ( .A(n_324), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_SL g375 ( .A(n_324), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_324), .B(n_391), .Y(n_457) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI21xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_340), .B(n_345), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_337), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_337), .B(n_342), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_338), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g400 ( .A(n_338), .Y(n_400) );
INVx1_ASAP7_75t_L g404 ( .A(n_338), .Y(n_404) );
AND2x2_ASAP7_75t_L g488 ( .A(n_338), .B(n_456), .Y(n_488) );
AND2x2_ASAP7_75t_L g491 ( .A(n_338), .B(n_408), .Y(n_491) );
INVx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_SL g342 ( .A(n_343), .B(n_344), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_343), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g470 ( .A(n_347), .Y(n_470) );
AND2x2_ASAP7_75t_L g361 ( .A(n_348), .B(n_362), .Y(n_361) );
NAND4xp75_ASAP7_75t_L g351 ( .A(n_352), .B(n_371), .C(n_392), .D(n_410), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_363), .Y(n_352) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g441 ( .A(n_355), .B(n_442), .Y(n_441) );
NAND2x1p5_ASAP7_75t_L g427 ( .A(n_356), .B(n_421), .Y(n_427) );
NAND2xp5_ASAP7_75t_R g443 ( .A(n_359), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g493 ( .A(n_359), .Y(n_493) );
INVx2_ASAP7_75t_L g406 ( .A(n_361), .Y(n_406) );
BUFx3_ASAP7_75t_L g398 ( .A(n_362), .Y(n_398) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g449 ( .A(n_367), .Y(n_449) );
AND2x2_ASAP7_75t_L g403 ( .A(n_369), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g425 ( .A(n_370), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_376), .B(n_378), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_374), .B(n_408), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_375), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_377), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_382), .B1(n_384), .B2(n_388), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
OA21x2_ASAP7_75t_L g393 ( .A1(n_386), .A2(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g414 ( .A(n_386), .Y(n_414) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g445 ( .A(n_387), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g453 ( .A(n_387), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_388), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g423 ( .A(n_391), .B(n_424), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_399), .B(n_401), .Y(n_392) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g440 ( .A(n_397), .B(n_441), .Y(n_440) );
INVx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_404), .Y(n_452) );
INVx2_ASAP7_75t_SL g444 ( .A(n_408), .Y(n_444) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_422), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_415), .B1(n_417), .B2(n_420), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g473 ( .A(n_417), .Y(n_473) );
NOR2x1_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_465), .Y(n_428) );
NAND3xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_438), .C(n_450), .Y(n_429) );
NOR2x1_ASAP7_75t_L g430 ( .A(n_431), .B(n_435), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
AOI22xp33_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_443), .B1(n_445), .B2(n_447), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NOR3xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .C(n_461), .Y(n_450) );
AOI21xp33_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_458), .B(n_459), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_484), .Y(n_465) );
NOR3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_474), .C(n_481), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B1(n_472), .B2(n_473), .Y(n_467) );
OR2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
NOR3xp33_ASAP7_75t_L g481 ( .A(n_475), .B(n_480), .C(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AOI222xp33_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_488), .B1(n_489), .B2(n_491), .C1(n_492), .C2(n_493), .Y(n_484) );
INVx1_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g822 ( .A(n_494), .Y(n_822) );
AND2x4_ASAP7_75t_L g494 ( .A(n_495), .B(n_678), .Y(n_494) );
NOR3xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_633), .C(n_662), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_497), .B(n_606), .Y(n_496) );
AOI221xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_531), .B1(n_552), .B2(n_563), .C(n_567), .Y(n_497) );
INVx3_ASAP7_75t_SL g723 ( .A(n_498), .Y(n_723) );
AND2x2_ASAP7_75t_SL g498 ( .A(n_499), .B(n_510), .Y(n_498) );
NAND2x1p5_ASAP7_75t_L g569 ( .A(n_499), .B(n_522), .Y(n_569) );
INVx4_ASAP7_75t_L g604 ( .A(n_499), .Y(n_604) );
AND2x2_ASAP7_75t_L g626 ( .A(n_499), .B(n_523), .Y(n_626) );
AND2x2_ASAP7_75t_L g632 ( .A(n_499), .B(n_571), .Y(n_632) );
INVx5_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g601 ( .A(n_500), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_500), .B(n_522), .Y(n_677) );
AND2x2_ASAP7_75t_L g682 ( .A(n_500), .B(n_523), .Y(n_682) );
AND2x2_ASAP7_75t_L g694 ( .A(n_500), .B(n_555), .Y(n_694) );
NOR2x1_ASAP7_75t_SL g733 ( .A(n_500), .B(n_571), .Y(n_733) );
OR2x6_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
INVx2_ASAP7_75t_L g562 ( .A(n_510), .Y(n_562) );
AND2x2_ASAP7_75t_L g666 ( .A(n_510), .B(n_615), .Y(n_666) );
AND2x2_ASAP7_75t_L g763 ( .A(n_510), .B(n_694), .Y(n_763) );
AND2x4_ASAP7_75t_L g510 ( .A(n_511), .B(n_522), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g595 ( .A(n_512), .Y(n_595) );
INVx2_ASAP7_75t_L g617 ( .A(n_512), .Y(n_617) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_520), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_513), .B(n_521), .Y(n_520) );
AO21x2_ASAP7_75t_L g571 ( .A1(n_513), .A2(n_514), .B(n_520), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_519), .Y(n_514) );
AND2x2_ASAP7_75t_L g592 ( .A(n_522), .B(n_554), .Y(n_592) );
INVx2_ASAP7_75t_L g596 ( .A(n_522), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_522), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g695 ( .A(n_522), .B(n_660), .Y(n_695) );
OR2x2_ASAP7_75t_L g742 ( .A(n_522), .B(n_555), .Y(n_742) );
INVx4_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_523), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_529), .Y(n_524) );
AND2x2_ASAP7_75t_L g739 ( .A(n_531), .B(n_620), .Y(n_739) );
AND2x2_ASAP7_75t_L g789 ( .A(n_531), .B(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
OR2x2_ASAP7_75t_L g665 ( .A(n_532), .B(n_609), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_543), .Y(n_532) );
AND2x2_ASAP7_75t_L g598 ( .A(n_533), .B(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g628 ( .A(n_533), .B(n_629), .Y(n_628) );
AND2x4_ASAP7_75t_L g649 ( .A(n_533), .B(n_629), .Y(n_649) );
AND2x4_ASAP7_75t_L g684 ( .A(n_533), .B(n_672), .Y(n_684) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g565 ( .A(n_534), .Y(n_565) );
OAI21x1_ASAP7_75t_SL g534 ( .A1(n_535), .A2(n_537), .B(n_541), .Y(n_534) );
INVx1_ASAP7_75t_L g542 ( .A(n_536), .Y(n_542) );
AND2x2_ASAP7_75t_L g611 ( .A(n_543), .B(n_564), .Y(n_611) );
AND2x2_ASAP7_75t_L g697 ( .A(n_543), .B(n_629), .Y(n_697) );
AND2x2_ASAP7_75t_L g708 ( .A(n_543), .B(n_573), .Y(n_708) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g572 ( .A(n_544), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g639 ( .A(n_544), .B(n_574), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_546), .B(n_550), .Y(n_545) );
INVx2_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_562), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_554), .B(n_604), .Y(n_661) );
AND2x2_ASAP7_75t_L g705 ( .A(n_554), .B(n_571), .Y(n_705) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_555), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g615 ( .A(n_555), .Y(n_615) );
BUFx3_ASAP7_75t_L g624 ( .A(n_555), .Y(n_624) );
AND2x2_ASAP7_75t_L g647 ( .A(n_555), .B(n_617), .Y(n_647) );
OAI322xp33_ASAP7_75t_L g567 ( .A1(n_562), .A2(n_568), .A3(n_572), .B1(n_582), .B2(n_590), .C1(n_597), .C2(n_602), .Y(n_567) );
INVx1_ASAP7_75t_L g728 ( .A(n_562), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_563), .B(n_603), .Y(n_602) );
AND2x4_ASAP7_75t_L g641 ( .A(n_563), .B(n_583), .Y(n_641) );
INVx2_ASAP7_75t_L g686 ( .A(n_563), .Y(n_686) );
AND2x2_ASAP7_75t_L g702 ( .A(n_563), .B(n_644), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_563), .B(n_720), .Y(n_750) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
AND2x2_ASAP7_75t_SL g653 ( .A(n_564), .B(n_629), .Y(n_653) );
OR2x2_ASAP7_75t_L g674 ( .A(n_564), .B(n_591), .Y(n_674) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
BUFx2_ASAP7_75t_L g646 ( .A(n_565), .Y(n_646) );
INVx2_ASAP7_75t_L g591 ( .A(n_566), .Y(n_591) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_566), .Y(n_593) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx2_ASAP7_75t_L g636 ( .A(n_569), .Y(n_636) );
INVxp67_ASAP7_75t_SL g656 ( .A(n_570), .Y(n_656) );
INVx1_ASAP7_75t_L g754 ( .A(n_570), .Y(n_754) );
INVxp67_ASAP7_75t_SL g769 ( .A(n_570), .Y(n_769) );
NAND2x1_ASAP7_75t_L g779 ( .A(n_572), .B(n_583), .Y(n_779) );
INVx1_ASAP7_75t_L g786 ( .A(n_572), .Y(n_786) );
BUFx2_ASAP7_75t_L g620 ( .A(n_573), .Y(n_620) );
AND2x2_ASAP7_75t_L g696 ( .A(n_573), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
BUFx3_ASAP7_75t_L g605 ( .A(n_574), .Y(n_605) );
INVxp67_ASAP7_75t_L g609 ( .A(n_574), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_580), .Y(n_575) );
NAND3xp33_ASAP7_75t_L g597 ( .A(n_582), .B(n_598), .C(n_600), .Y(n_597) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_SL g618 ( .A(n_583), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_583), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g770 ( .A(n_583), .B(n_719), .Y(n_770) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g672 ( .A(n_584), .Y(n_672) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_584), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B1(n_593), .B2(n_594), .Y(n_590) );
AND2x4_ASAP7_75t_SL g719 ( .A(n_591), .B(n_599), .Y(n_719) );
AND2x2_ASAP7_75t_L g732 ( .A(n_592), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_593), .Y(n_734) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx2_ASAP7_75t_L g691 ( .A(n_595), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_595), .B(n_604), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_596), .B(n_614), .Y(n_613) );
AND3x2_ASAP7_75t_L g631 ( .A(n_596), .B(n_624), .C(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g655 ( .A(n_596), .Y(n_655) );
AND2x2_ASAP7_75t_L g768 ( .A(n_596), .B(n_769), .Y(n_768) );
BUFx2_ASAP7_75t_L g644 ( .A(n_599), .Y(n_644) );
INVx1_ASAP7_75t_L g722 ( .A(n_599), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_600), .B(n_623), .Y(n_761) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_601), .B(n_705), .Y(n_710) );
AND2x4_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
AND2x2_ASAP7_75t_L g701 ( .A(n_604), .B(n_647), .Y(n_701) );
INVx1_ASAP7_75t_SL g652 ( .A(n_605), .Y(n_652) );
AND2x2_ASAP7_75t_L g760 ( .A(n_605), .B(n_672), .Y(n_760) );
AND2x2_ASAP7_75t_L g781 ( .A(n_605), .B(n_653), .Y(n_781) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_612), .B1(n_618), .B2(n_621), .C(n_627), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g773 ( .A(n_609), .Y(n_773) );
AOI21xp33_ASAP7_75t_SL g627 ( .A1(n_610), .A2(n_628), .B(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g619 ( .A(n_611), .B(n_620), .Y(n_619) );
AOI222xp33_ASAP7_75t_L g642 ( .A1(n_611), .A2(n_643), .B1(n_645), .B2(n_650), .C1(n_654), .C2(n_657), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_611), .B(n_760), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_612), .A2(n_641), .B1(n_664), .B2(n_666), .Y(n_663) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g648 ( .A(n_615), .Y(n_648) );
AND2x2_ASAP7_75t_L g767 ( .A(n_615), .B(n_733), .Y(n_767) );
OAI32xp33_ASAP7_75t_L g771 ( .A1(n_615), .A2(n_640), .A3(n_692), .B1(n_700), .B2(n_772), .Y(n_771) );
AND2x2_ASAP7_75t_L g776 ( .A(n_615), .B(n_626), .Y(n_776) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g660 ( .A(n_617), .Y(n_660) );
OAI21xp5_ASAP7_75t_SL g667 ( .A1(n_618), .A2(n_668), .B(n_675), .Y(n_667) );
INVx1_ASAP7_75t_L g731 ( .A(n_620), .Y(n_731) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
AND2x2_ASAP7_75t_L g635 ( .A(n_623), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g643 ( .A(n_626), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g716 ( .A(n_626), .B(n_647), .Y(n_716) );
INVx1_ASAP7_75t_SL g787 ( .A(n_628), .Y(n_787) );
AND2x2_ASAP7_75t_L g721 ( .A(n_629), .B(n_722), .Y(n_721) );
OAI222xp33_ASAP7_75t_L g774 ( .A1(n_630), .A2(n_683), .B1(n_762), .B2(n_775), .C1(n_777), .C2(n_779), .Y(n_774) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x4_ASAP7_75t_L g747 ( .A(n_632), .B(n_748), .Y(n_747) );
OAI21xp33_ASAP7_75t_SL g633 ( .A1(n_634), .A2(n_637), .B(n_642), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_636), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g715 ( .A(n_638), .Y(n_715) );
INVx1_ASAP7_75t_L g683 ( .A(n_639), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_639), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g737 ( .A(n_644), .Y(n_737) );
AO22x1_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B1(n_648), .B2(n_649), .Y(n_645) );
OAI322xp33_ASAP7_75t_L g757 ( .A1(n_646), .A2(n_707), .A3(n_710), .B1(n_758), .B2(n_759), .C1(n_761), .C2(n_762), .Y(n_757) );
AND2x2_ASAP7_75t_SL g681 ( .A(n_647), .B(n_682), .Y(n_681) );
OR2x2_ASAP7_75t_L g676 ( .A(n_648), .B(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g736 ( .A(n_649), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g778 ( .A(n_649), .B(n_708), .Y(n_778) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g758 ( .A(n_652), .Y(n_758) );
INVx1_ASAP7_75t_SL g687 ( .A(n_653), .Y(n_687) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
OR2x2_ASAP7_75t_L g689 ( .A(n_661), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g727 ( .A(n_661), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_667), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_673), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g700 ( .A(n_671), .B(n_686), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_671), .B(n_708), .Y(n_707) );
BUFx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g730 ( .A(n_674), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NOR2x1_ASAP7_75t_L g678 ( .A(n_679), .B(n_743), .Y(n_678) );
NAND4xp25_ASAP7_75t_L g679 ( .A(n_680), .B(n_698), .C(n_711), .D(n_724), .Y(n_679) );
AOI322xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_683), .A3(n_684), .B1(n_685), .B2(n_688), .C1(n_693), .C2(n_696), .Y(n_680) );
AOI211xp5_ASAP7_75t_L g780 ( .A1(n_681), .A2(n_781), .B(n_782), .C(n_785), .Y(n_780) );
AND2x2_ASAP7_75t_L g792 ( .A(n_682), .B(n_769), .Y(n_792) );
INVx1_ASAP7_75t_L g714 ( .A(n_684), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_684), .B(n_719), .Y(n_756) );
NAND2xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_692), .B(n_705), .Y(n_772) );
AND2x4_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
AOI222xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .B1(n_702), .B2(n_703), .C1(n_706), .C2(n_709), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_701), .A2(n_712), .B1(n_715), .B2(n_716), .C(n_717), .Y(n_711) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AOI21xp33_ASAP7_75t_SL g717 ( .A1(n_718), .A2(n_720), .B(n_723), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_729), .B1(n_732), .B2(n_734), .C(n_735), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_727), .B(n_728), .Y(n_726) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g784 ( .A(n_733), .Y(n_784) );
AOI21xp33_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_738), .B(n_740), .Y(n_735) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
INVx2_ASAP7_75t_L g748 ( .A(n_742), .Y(n_748) );
OR2x2_ASAP7_75t_L g783 ( .A(n_742), .B(n_784), .Y(n_783) );
NAND3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_764), .C(n_780), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_757), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_749), .B(n_751), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_755), .Y(n_751) );
INVx1_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
AOI221xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_770), .B1(n_771), .B2(n_773), .C(n_774), .Y(n_764) );
INVxp67_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NOR2x1_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_779), .B(n_783), .Y(n_782) );
O2A1O1Ixp33_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_787), .B(n_788), .C(n_791), .Y(n_785) );
INVxp67_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
CKINVDCx11_ASAP7_75t_R g793 ( .A(n_794), .Y(n_793) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_794), .Y(n_799) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx3_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
INVx2_ASAP7_75t_SL g802 ( .A(n_803), .Y(n_802) );
INVx3_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVxp67_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_806), .A2(n_811), .B(n_820), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
BUFx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
BUFx3_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_SL g813 ( .A(n_814), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_815), .B(n_819), .Y(n_818) );
CKINVDCx11_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
CKINVDCx8_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
INVx3_ASAP7_75t_SL g823 ( .A(n_824), .Y(n_823) );
endmodule