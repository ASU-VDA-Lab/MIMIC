module fake_jpeg_28524_n_100 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_100);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_100;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_45),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_3),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_4),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_4),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_5),
.Y(n_57)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_17),
.B(n_31),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp67_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_39),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_52),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_33),
.B1(n_42),
.B2(n_35),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_58),
.B1(n_11),
.B2(n_12),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_5),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_42),
.B1(n_35),
.B2(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_6),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_6),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_72),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_59),
.B(n_7),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_74),
.B1(n_13),
.B2(n_14),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_84),
.Y(n_91)
);

CKINVDCx10_ASAP7_75t_R g81 ( 
.A(n_69),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_16),
.B(n_18),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_70),
.C(n_62),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_87),
.B(n_81),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_70),
.C(n_22),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_90),
.B1(n_82),
.B2(n_77),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_93),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_91),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_88),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_75),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_76),
.B(n_86),
.Y(n_98)
);

AOI31xp33_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_83),
.A3(n_29),
.B(n_32),
.Y(n_99)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_99),
.Y(n_100)
);


endmodule