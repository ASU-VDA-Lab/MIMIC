module fake_jpeg_12600_n_153 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_21),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_44),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_18),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_9),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_66),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_70),
.B1(n_71),
.B2(n_53),
.Y(n_81)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_66),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_56),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_28),
.B1(n_43),
.B2(n_42),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_47),
.Y(n_75)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_85),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_82),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_51),
.B1(n_75),
.B2(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_87),
.Y(n_98)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_61),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_7),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_89),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_63),
.B(n_48),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_101),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_46),
.B1(n_64),
.B2(n_50),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_93),
.A2(n_97),
.B1(n_20),
.B2(n_24),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_89),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_96),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_55),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_64),
.B1(n_51),
.B2(n_75),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_100),
.B1(n_106),
.B2(n_29),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_60),
.B1(n_59),
.B2(n_68),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_58),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_16),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_105),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_7),
.B(n_8),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_27),
.B1(n_40),
.B2(n_38),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_10),
.B(n_11),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_19),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_119),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_12),
.C(n_13),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_25),
.C(n_33),
.Y(n_134)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_124),
.Y(n_130)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_126),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_101),
.B1(n_30),
.B2(n_31),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_37),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_136),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_35),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_131),
.A2(n_125),
.B(n_118),
.C(n_120),
.D(n_117),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_140),
.B(n_141),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_122),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_144),
.C(n_135),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_126),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_142),
.C(n_127),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_149),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_147),
.A2(n_138),
.B(n_137),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

OAI321xp33_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_145),
.A3(n_130),
.B1(n_133),
.B2(n_127),
.C(n_141),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_132),
.Y(n_153)
);


endmodule