module fake_netlist_6_2160_n_4257 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_442, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_443, n_246, n_38, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_417, n_14, n_446, n_89, n_374, n_366, n_407, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_433, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_54, n_328, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4257);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_89;
input n_374;
input n_366;
input n_407;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_433;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4257;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_801;
wire n_3766;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3783;
wire n_700;
wire n_3773;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_3844;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4168;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_2324;
wire n_1854;
wire n_1575;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_4134;
wire n_3465;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_471;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4087;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_461;
wire n_1371;
wire n_1285;
wire n_873;
wire n_2886;
wire n_2974;
wire n_3946;
wire n_1985;
wire n_4213;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_852;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_836;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_3979;
wire n_616;
wire n_658;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_2212;
wire n_3929;
wire n_758;
wire n_516;
wire n_3494;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_491;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_4187;
wire n_940;
wire n_770;
wire n_567;
wire n_1971;
wire n_1781;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_538;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_494;
wire n_539;
wire n_493;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_454;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2551;
wire n_2364;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_659;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_913;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4071;
wire n_4255;
wire n_3506;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_473;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_3943;
wire n_564;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_451;
wire n_824;
wire n_686;
wire n_4102;
wire n_757;
wire n_594;
wire n_2113;
wire n_1641;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_577;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_619;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_572;
wire n_813;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_606;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_3910;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4009;
wire n_2633;
wire n_483;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_630;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_792;
wire n_2522;
wire n_476;
wire n_3949;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_982;
wire n_2674;
wire n_2832;
wire n_4226;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_932;
wire n_2831;
wire n_2998;
wire n_3446;
wire n_4158;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_905;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_2692;
wire n_993;
wire n_3842;
wire n_689;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_966;
wire n_3888;
wire n_2908;
wire n_3168;
wire n_764;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4161;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3055;
wire n_3092;
wire n_3492;
wire n_3966;
wire n_3895;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_1014;
wire n_3734;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_882;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_586;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_2711;
wire n_3490;
wire n_4199;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_702;
wire n_2749;
wire n_2008;
wire n_3346;
wire n_2192;
wire n_3298;
wire n_2345;
wire n_2254;
wire n_3281;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_4072;
wire n_3940;
wire n_4220;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_690;
wire n_2347;
wire n_1886;
wire n_2092;
wire n_3917;
wire n_1654;
wire n_816;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3428;
wire n_3153;
wire n_3410;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2519;
wire n_2319;
wire n_4043;
wire n_825;
wire n_728;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_515;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_696;
wire n_1515;
wire n_961;
wire n_3510;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_593;
wire n_4169;
wire n_514;
wire n_4055;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_3271;
wire n_950;
wire n_4248;
wire n_2812;
wire n_484;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_590;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_462;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_2431;
wire n_3073;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3780;
wire n_3696;
wire n_4082;
wire n_1634;
wire n_2078;
wire n_3252;
wire n_2932;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_3253;
wire n_3337;
wire n_3431;
wire n_3209;
wire n_3450;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_4002;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_449;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_495;
wire n_815;
wire n_3953;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_4191;
wire n_1364;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_963;
wire n_639;
wire n_2767;
wire n_794;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_872;
wire n_1139;
wire n_1714;
wire n_3922;
wire n_3179;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_542;
wire n_847;
wire n_851;
wire n_644;
wire n_682;
wire n_2537;
wire n_2897;
wire n_3970;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_3171;
wire n_791;
wire n_1913;
wire n_4216;
wire n_3608;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_4162;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3975;
wire n_3782;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_765;
wire n_987;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_705;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_3887;
wire n_1022;
wire n_614;
wire n_529;
wire n_2307;
wire n_2069;
wire n_3704;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_4096;
wire n_1431;
wire n_4123;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_1809;
wire n_3119;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_3731;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_4218;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_478;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_3693;
wire n_3788;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_777;
wire n_1299;
wire n_2896;
wire n_526;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3325;
wire n_3203;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_4175;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_3893;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_1507;
wire n_2482;
wire n_552;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_745;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1774;
wire n_623;
wire n_1048;
wire n_1398;
wire n_1201;
wire n_884;
wire n_2682;
wire n_2354;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_3393;
wire n_527;
wire n_683;
wire n_811;
wire n_474;
wire n_1207;
wire n_2442;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3451;
wire n_3480;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_2545;
wire n_3577;
wire n_3540;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_589;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2581;
wire n_1363;
wire n_2294;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3591;
wire n_767;
wire n_3641;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_477;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1564;
wire n_1736;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_505;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_3909;
wire n_3944;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2301;
wire n_2209;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_511;
wire n_2990;
wire n_3847;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2552;
wire n_2410;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3323;
wire n_3364;
wire n_4020;
wire n_4176;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_453;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_1745;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_497;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1892;
wire n_1459;
wire n_1614;
wire n_3188;
wire n_3742;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4034;
wire n_1617;
wire n_4056;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_463;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_4206;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_3862;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_4132;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1832;
wire n_1645;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_3016;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2993;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_1129;
wire n_4030;
wire n_4126;
wire n_3870;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_664;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_587;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_607;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3194;
wire n_3113;
wire n_3250;
wire n_1934;
wire n_3276;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_617;
wire n_3886;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3926;
wire n_3797;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_4234;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_517;
wire n_4211;
wire n_4182;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_621;
wire n_1037;
wire n_1397;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_3592;
wire n_468;
wire n_2755;
wire n_3141;
wire n_923;
wire n_504;
wire n_1409;
wire n_4230;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_466;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_4155;
wire n_2740;
wire n_746;
wire n_4238;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_3042;
wire n_1356;
wire n_1589;
wire n_3213;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4109;
wire n_4192;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_4038;
wire n_3957;
wire n_2790;
wire n_4131;
wire n_2808;
wire n_2037;
wire n_4195;
wire n_4159;
wire n_3710;
wire n_3784;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_1870;
wire n_2964;
wire n_4174;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_662;
wire n_3475;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_450;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2699;
wire n_2272;
wire n_2046;
wire n_2200;
wire n_3029;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_456;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_482;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3439;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_4135;
wire n_2871;
wire n_4209;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_3858;
wire n_4183;
wire n_1489;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_543;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_4040;
wire n_804;
wire n_464;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_799;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1475;
wire n_1229;
wire n_2759;
wire n_3457;
wire n_2945;
wire n_3061;
wire n_3517;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3469;
wire n_3932;
wire n_2266;
wire n_2960;
wire n_3958;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_3156;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_502;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1794;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1650;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_834;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_743;
wire n_766;
wire n_3124;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2888;
wire n_2885;
wire n_2715;
wire n_2793;
wire n_1804;
wire n_2923;
wire n_3711;
wire n_3776;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_3308;
wire n_1113;
wire n_2833;
wire n_1600;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_841;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_4203;
wire n_3808;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1882;
wire n_2951;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_3726;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_591;
wire n_3758;
wire n_1879;
wire n_853;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_680;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_1976;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_2969;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_535;
wire n_691;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_1598;
wire n_3493;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_3898;
wire n_2284;
wire n_3739;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_1303;
wire n_761;
wire n_2769;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_4106;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4027;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_647;
wire n_4160;
wire n_4231;
wire n_844;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2255;
wire n_2112;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_3486;
wire n_4086;
wire n_908;
wire n_752;
wire n_2649;
wire n_2721;
wire n_944;
wire n_3556;
wire n_2034;
wire n_576;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_2444;
wire n_839;
wire n_2743;
wire n_3962;
wire n_708;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_4166;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_498;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3256;
wire n_1276;
wire n_3868;
wire n_3802;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4142;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_492;
wire n_3680;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_719;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_455;
wire n_2666;
wire n_4105;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_4244;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_829;
wire n_1156;
wire n_1362;
wire n_3123;
wire n_2600;
wire n_984;
wire n_3380;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_570;
wire n_859;
wire n_2033;
wire n_3086;
wire n_735;
wire n_4104;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_3285;
wire n_519;
wire n_4208;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_2723;
wire n_2440;
wire n_2233;
wire n_481;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_3989;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_1606;
wire n_810;
wire n_4108;
wire n_1133;
wire n_635;
wire n_1194;
wire n_3374;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_4051;
wire n_1051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_3383;
wire n_3709;
wire n_753;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_467;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_4148;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_4057;
wire n_2968;
wire n_4201;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_3903;
wire n_730;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_3896;
wire n_2774;
wire n_3815;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_640;
wire n_4129;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3584;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_457;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_531;
wire n_827;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g449 ( 
.A(n_11),
.Y(n_449)
);

BUFx10_ASAP7_75t_L g450 ( 
.A(n_432),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_288),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_336),
.Y(n_452)
);

BUFx4f_ASAP7_75t_SL g453 ( 
.A(n_439),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_266),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_345),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_13),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_25),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_115),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_354),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_12),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_56),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_160),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_316),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_75),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_54),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_69),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_253),
.Y(n_467)
);

BUFx10_ASAP7_75t_L g468 ( 
.A(n_100),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_36),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_344),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_434),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_114),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_349),
.Y(n_473)
);

INVxp33_ASAP7_75t_SL g474 ( 
.A(n_26),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_318),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_421),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_447),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_193),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_288),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_247),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_262),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_48),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_168),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_374),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_378),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_226),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_325),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_245),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_384),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_282),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_90),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_333),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_149),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_153),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_208),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_224),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_257),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_150),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_320),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_357),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_339),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_58),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_8),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_406),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_91),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_25),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_110),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_255),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_418),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_131),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_422),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_286),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_152),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_135),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_196),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_362),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_297),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_7),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_309),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_376),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_228),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_6),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_215),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_87),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_278),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_303),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_315),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_245),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_59),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_122),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_381),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_431),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_402),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_275),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_82),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_389),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_115),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_277),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_401),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_253),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_394),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_42),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_442),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_133),
.Y(n_544)
);

BUFx8_ASAP7_75t_SL g545 ( 
.A(n_226),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_183),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_107),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_90),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_155),
.Y(n_549)
);

CKINVDCx14_ASAP7_75t_R g550 ( 
.A(n_207),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_98),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_420),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_342),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_264),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_188),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_48),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_332),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_192),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_319),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_300),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_57),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_33),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_31),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_266),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_237),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_437),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_220),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_416),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_204),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_386),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_399),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_16),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_427),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_400),
.Y(n_574)
);

BUFx10_ASAP7_75t_L g575 ( 
.A(n_145),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_368),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_142),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_444),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_268),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_105),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_286),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_236),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_367),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_255),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_408),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_162),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_69),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_139),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_59),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_34),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_260),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_158),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_172),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_30),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_238),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_155),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_75),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_37),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_359),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_211),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_379),
.Y(n_601)
);

CKINVDCx16_ASAP7_75t_R g602 ( 
.A(n_312),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_438),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_230),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_63),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_429),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_88),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_314),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_14),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_250),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_163),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_154),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_97),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_177),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_348),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_403),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_329),
.Y(n_617)
);

CKINVDCx14_ASAP7_75t_R g618 ( 
.A(n_328),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_102),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_387),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_391),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_285),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_148),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_113),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_216),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_100),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_299),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_166),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_297),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_151),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_3),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_419),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_436),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_26),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_272),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_8),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_16),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_161),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_270),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_396),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_18),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_143),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_57),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_148),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_53),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_301),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_293),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_390),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_78),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_187),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_352),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_172),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_294),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_364),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_66),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_168),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_110),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_88),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_313),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_248),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_292),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_22),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_247),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_121),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_232),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_106),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_181),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_212),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_241),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_265),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_94),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_12),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_14),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_191),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_281),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_76),
.Y(n_676)
);

CKINVDCx16_ASAP7_75t_R g677 ( 
.A(n_118),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_111),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_198),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_20),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_250),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_127),
.Y(n_682)
);

CKINVDCx14_ASAP7_75t_R g683 ( 
.A(n_36),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_341),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_353),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_279),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_363),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_276),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_424),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_0),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_440),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_263),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_105),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_217),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_146),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_181),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_67),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_358),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_182),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_365),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_289),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_448),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_183),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_40),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_251),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_53),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_215),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_317),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_292),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_201),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_55),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_132),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_257),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_79),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_96),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_195),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_142),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_289),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_267),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_392),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_412),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_405),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_383),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_294),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_430),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_191),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_256),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_240),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_360),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_194),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_277),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_274),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_129),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_121),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_244),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_199),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_118),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_150),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_371),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_125),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_103),
.Y(n_741)
);

BUFx10_ASAP7_75t_L g742 ( 
.A(n_111),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_23),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_269),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_213),
.Y(n_745)
);

CKINVDCx14_ASAP7_75t_R g746 ( 
.A(n_311),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_43),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_157),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_441),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_205),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_260),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_116),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_38),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_251),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_423),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_216),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_303),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_236),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_66),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_410),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_2),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_323),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_220),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_194),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_92),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_351),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_87),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_138),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_230),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_166),
.Y(n_770)
);

CKINVDCx16_ASAP7_75t_R g771 ( 
.A(n_164),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_263),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_164),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_256),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_123),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_304),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_330),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_249),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_76),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_527),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_456),
.Y(n_781)
);

NOR2xp67_ASAP7_75t_L g782 ( 
.A(n_631),
.B(n_0),
.Y(n_782)
);

BUFx5_ASAP7_75t_L g783 ( 
.A(n_459),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_545),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_456),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_527),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_545),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_631),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_452),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_456),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_456),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_456),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_456),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_498),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_498),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_498),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_536),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_722),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_498),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_498),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_498),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_523),
.Y(n_802)
);

BUFx2_ASAP7_75t_SL g803 ( 
.A(n_471),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_455),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_473),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_523),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_523),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_475),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_476),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_523),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_484),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_499),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_557),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_504),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_523),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_523),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_597),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_597),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_597),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_509),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_511),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_516),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_535),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_597),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_597),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_621),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_597),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_676),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_676),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_722),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_519),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_676),
.Y(n_832)
);

NOR2xp67_ASAP7_75t_L g833 ( 
.A(n_703),
.B(n_1),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_676),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_676),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_676),
.Y(n_836)
);

BUFx8_ASAP7_75t_SL g837 ( 
.A(n_535),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_747),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_532),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_747),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_554),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_747),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_648),
.Y(n_843)
);

INVx1_ASAP7_75t_SL g844 ( 
.A(n_554),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_747),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_689),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_533),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_539),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_541),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_543),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_747),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_747),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_449),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_553),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_568),
.Y(n_855)
);

INVxp33_ASAP7_75t_SL g856 ( 
.A(n_703),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_570),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_449),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_449),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_464),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_738),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_571),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_464),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_464),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_480),
.Y(n_865)
);

INVxp67_ASAP7_75t_SL g866 ( 
.A(n_760),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_762),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_480),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_480),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_512),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_574),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_576),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_512),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_512),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_521),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_521),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_601),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_521),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_549),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_606),
.Y(n_880)
);

INVxp67_ASAP7_75t_SL g881 ( 
.A(n_760),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_608),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_549),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_549),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_615),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_616),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_588),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_588),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_588),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_624),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_722),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_624),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_658),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_624),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_647),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_647),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_738),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_647),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_649),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_658),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_617),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_649),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_620),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_649),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_632),
.Y(n_905)
);

INVxp33_ASAP7_75t_L g906 ( 
.A(n_775),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_777),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_753),
.Y(n_908)
);

INVx1_ASAP7_75t_SL g909 ( 
.A(n_753),
.Y(n_909)
);

CKINVDCx16_ASAP7_75t_R g910 ( 
.A(n_503),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_777),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_656),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_656),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_656),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_659),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_618),
.Y(n_916)
);

INVx1_ASAP7_75t_SL g917 ( 
.A(n_466),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_740),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_684),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_775),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_685),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_740),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_777),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_740),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_748),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_496),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_687),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_691),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_748),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_698),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_702),
.Y(n_931)
);

XOR2xp5_ASAP7_75t_L g932 ( 
.A(n_577),
.B(n_1),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_720),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_721),
.Y(n_934)
);

INVx1_ASAP7_75t_SL g935 ( 
.A(n_534),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_748),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_725),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_757),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_757),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_757),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_618),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_746),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_774),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_774),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_774),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_503),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_488),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_566),
.B(n_654),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_488),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_729),
.Y(n_950)
);

NOR2xp67_ASAP7_75t_L g951 ( 
.A(n_465),
.B(n_2),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_739),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_488),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_562),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_562),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_749),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_477),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_562),
.Y(n_958)
);

INVxp33_ASAP7_75t_L g959 ( 
.A(n_458),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_527),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_527),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_572),
.Y(n_962)
);

CKINVDCx14_ASAP7_75t_R g963 ( 
.A(n_550),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_755),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_477),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_550),
.Y(n_966)
);

CKINVDCx16_ASAP7_75t_R g967 ( 
.A(n_677),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_572),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_683),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_683),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_477),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_572),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_494),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_607),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_607),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_451),
.Y(n_976)
);

INVxp67_ASAP7_75t_SL g977 ( 
.A(n_566),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_454),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_607),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_531),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_642),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_457),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_461),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_467),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_642),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_472),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_642),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_673),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_673),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_540),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_478),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_481),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_673),
.Y(n_993)
);

INVxp33_ASAP7_75t_SL g994 ( 
.A(n_482),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_450),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_486),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_677),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_704),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_531),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_704),
.Y(n_1000)
);

CKINVDCx16_ASAP7_75t_R g1001 ( 
.A(n_771),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_704),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_494),
.Y(n_1003)
);

INVxp67_ASAP7_75t_L g1004 ( 
.A(n_458),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_490),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_462),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_491),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_493),
.Y(n_1008)
);

NOR2xp67_ASAP7_75t_L g1009 ( 
.A(n_465),
.B(n_3),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_495),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_462),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_469),
.Y(n_1012)
);

CKINVDCx20_ASAP7_75t_R g1013 ( 
.A(n_746),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_487),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_469),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_497),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_531),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_502),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_479),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_479),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_483),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_483),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_527),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_559),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_487),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_505),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_514),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_514),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_515),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_515),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_506),
.Y(n_1031)
);

CKINVDCx14_ASAP7_75t_R g1032 ( 
.A(n_468),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_450),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_508),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_510),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_518),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_513),
.Y(n_1037)
);

INVx1_ASAP7_75t_SL g1038 ( 
.A(n_595),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_518),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_517),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_652),
.Y(n_1041)
);

CKINVDCx16_ASAP7_75t_R g1042 ( 
.A(n_771),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_501),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_525),
.Y(n_1044)
);

INVxp67_ASAP7_75t_SL g1045 ( 
.A(n_654),
.Y(n_1045)
);

BUFx8_ASAP7_75t_SL g1046 ( 
.A(n_577),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_522),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_526),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_528),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_522),
.Y(n_1050)
);

INVxp67_ASAP7_75t_SL g1051 ( 
.A(n_459),
.Y(n_1051)
);

INVxp67_ASAP7_75t_SL g1052 ( 
.A(n_463),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_529),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_524),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_524),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_547),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_501),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_547),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_602),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_530),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_548),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_548),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_555),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_527),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_555),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_450),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_559),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_559),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_556),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_537),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_538),
.Y(n_1071)
);

INVxp67_ASAP7_75t_L g1072 ( 
.A(n_556),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_560),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_578),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_560),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_668),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_544),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_567),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_567),
.Y(n_1079)
);

INVxp33_ASAP7_75t_L g1080 ( 
.A(n_580),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_450),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_580),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_582),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_582),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_551),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_558),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_561),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_563),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_587),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_587),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_463),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_564),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_592),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_578),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_565),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_592),
.Y(n_1096)
);

CKINVDCx20_ASAP7_75t_R g1097 ( 
.A(n_602),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_569),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_579),
.Y(n_1099)
);

INVxp67_ASAP7_75t_SL g1100 ( 
.A(n_470),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_581),
.Y(n_1101)
);

INVxp67_ASAP7_75t_L g1102 ( 
.A(n_594),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_594),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_600),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_600),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_625),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_625),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_630),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_584),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_586),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_630),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_634),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_634),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_635),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_589),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_635),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_636),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_590),
.Y(n_1118)
);

INVxp67_ASAP7_75t_SL g1119 ( 
.A(n_470),
.Y(n_1119)
);

CKINVDCx16_ASAP7_75t_R g1120 ( 
.A(n_468),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_593),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_636),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_641),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_596),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_641),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_598),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_643),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_643),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_646),
.Y(n_1129)
);

BUFx2_ASAP7_75t_SL g1130 ( 
.A(n_471),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_604),
.Y(n_1131)
);

INVx2_ASAP7_75t_SL g1132 ( 
.A(n_468),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_552),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_453),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_605),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_609),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_610),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_453),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_646),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_612),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_613),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_653),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_614),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_789),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_947),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_947),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_804),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_815),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_797),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_805),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_813),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_949),
.Y(n_1152)
);

INVxp67_ASAP7_75t_SL g1153 ( 
.A(n_923),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_949),
.Y(n_1154)
);

INVxp67_ASAP7_75t_L g1155 ( 
.A(n_946),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_953),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_808),
.Y(n_1157)
);

INVxp67_ASAP7_75t_L g1158 ( 
.A(n_997),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_826),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_809),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_953),
.Y(n_1161)
);

CKINVDCx20_ASAP7_75t_R g1162 ( 
.A(n_843),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_954),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_954),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_811),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_812),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_955),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_948),
.B(n_489),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_814),
.Y(n_1169)
);

CKINVDCx20_ASAP7_75t_R g1170 ( 
.A(n_846),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_955),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_958),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_820),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_821),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_958),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_962),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_962),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_867),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_968),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_968),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_972),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_822),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_972),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_831),
.Y(n_1184)
);

CKINVDCx20_ASAP7_75t_R g1185 ( 
.A(n_916),
.Y(n_1185)
);

INVxp33_ASAP7_75t_SL g1186 ( 
.A(n_966),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_839),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_941),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_974),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_974),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_847),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_975),
.Y(n_1192)
);

INVxp67_ASAP7_75t_L g1193 ( 
.A(n_1126),
.Y(n_1193)
);

INVxp67_ASAP7_75t_L g1194 ( 
.A(n_1131),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_975),
.Y(n_1195)
);

CKINVDCx14_ASAP7_75t_R g1196 ( 
.A(n_1032),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_848),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_979),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_849),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_R g1200 ( 
.A(n_963),
.B(n_622),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_994),
.B(n_489),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_976),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_850),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_815),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_854),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_979),
.Y(n_1206)
);

INVxp67_ASAP7_75t_SL g1207 ( 
.A(n_923),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_981),
.Y(n_1208)
);

XOR2xp5_ASAP7_75t_L g1209 ( 
.A(n_932),
.B(n_638),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_855),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_985),
.Y(n_1211)
);

CKINVDCx16_ASAP7_75t_R g1212 ( 
.A(n_910),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_981),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_825),
.Y(n_1214)
);

CKINVDCx16_ASAP7_75t_R g1215 ( 
.A(n_910),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_857),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_862),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_871),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_872),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_942),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_877),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_880),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_977),
.B(n_492),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_823),
.B(n_460),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_987),
.Y(n_1225)
);

INVx1_ASAP7_75t_SL g1226 ( 
.A(n_917),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_781),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_1013),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_781),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_882),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_1134),
.Y(n_1231)
);

INVxp67_ASAP7_75t_SL g1232 ( 
.A(n_923),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_987),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_988),
.Y(n_1234)
);

INVxp67_ASAP7_75t_L g1235 ( 
.A(n_985),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_988),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_989),
.Y(n_1237)
);

INVxp67_ASAP7_75t_L g1238 ( 
.A(n_1132),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_885),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_1132),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_886),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_866),
.B(n_492),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_901),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_989),
.Y(n_1244)
);

CKINVDCx16_ASAP7_75t_R g1245 ( 
.A(n_967),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_903),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_978),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_993),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_1138),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_993),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_905),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1051),
.B(n_1052),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_998),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_998),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1014),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_1025),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_915),
.Y(n_1257)
);

INVxp33_ASAP7_75t_SL g1258 ( 
.A(n_969),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1000),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1000),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_919),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_921),
.B(n_471),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_927),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1002),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_928),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_930),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_1043),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_1057),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_1059),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_931),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_933),
.B(n_578),
.Y(n_1271)
);

INVxp67_ASAP7_75t_SL g1272 ( 
.A(n_798),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_934),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_937),
.B(n_603),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1002),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_785),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_825),
.Y(n_1277)
);

INVxp67_ASAP7_75t_L g1278 ( 
.A(n_837),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_982),
.Y(n_1279)
);

CKINVDCx20_ASAP7_75t_R g1280 ( 
.A(n_1097),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_798),
.B(n_830),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_785),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_950),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_790),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_881),
.B(n_520),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_790),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_967),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_791),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_830),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_893),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_791),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_952),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_792),
.Y(n_1293)
);

INVxp67_ASAP7_75t_SL g1294 ( 
.A(n_891),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_956),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1045),
.B(n_520),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_792),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_793),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_964),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_793),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1046),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_983),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_794),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_794),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_795),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_984),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_986),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_991),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_1001),
.Y(n_1309)
);

CKINVDCx16_ASAP7_75t_R g1310 ( 
.A(n_1001),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_992),
.B(n_573),
.Y(n_1311)
);

CKINVDCx16_ASAP7_75t_R g1312 ( 
.A(n_1042),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1042),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_996),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_795),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1005),
.Y(n_1316)
);

INVxp67_ASAP7_75t_SL g1317 ( 
.A(n_891),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_926),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_796),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1007),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1008),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1010),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_796),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_799),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1016),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_893),
.Y(n_1326)
);

INVxp33_ASAP7_75t_L g1327 ( 
.A(n_788),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_799),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1018),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_935),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_842),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_907),
.Y(n_1332)
);

INVxp33_ASAP7_75t_SL g1333 ( 
.A(n_970),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1026),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_1031),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_800),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1034),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_800),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_801),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_801),
.Y(n_1340)
);

INVxp67_ASAP7_75t_SL g1341 ( 
.A(n_907),
.Y(n_1341)
);

CKINVDCx16_ASAP7_75t_R g1342 ( 
.A(n_1120),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_802),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_802),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_990),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_SL g1346 ( 
.A(n_995),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1035),
.Y(n_1347)
);

INVxp67_ASAP7_75t_L g1348 ( 
.A(n_908),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1037),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_806),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1040),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1044),
.Y(n_1352)
);

INVxp33_ASAP7_75t_SL g1353 ( 
.A(n_784),
.Y(n_1353)
);

INVxp67_ASAP7_75t_SL g1354 ( 
.A(n_911),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_807),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_807),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_810),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_810),
.Y(n_1358)
);

CKINVDCx16_ASAP7_75t_R g1359 ( 
.A(n_1120),
.Y(n_1359)
);

CKINVDCx16_ASAP7_75t_R g1360 ( 
.A(n_1038),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_908),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_803),
.B(n_603),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_1041),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_816),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_1076),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_816),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1048),
.B(n_573),
.Y(n_1367)
);

CKINVDCx16_ASAP7_75t_R g1368 ( 
.A(n_995),
.Y(n_1368)
);

NAND2xp33_ASAP7_75t_R g1369 ( 
.A(n_1049),
.B(n_474),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1053),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_817),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1060),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_817),
.Y(n_1373)
);

INVxp67_ASAP7_75t_L g1374 ( 
.A(n_841),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1070),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_1071),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_818),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_786),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_818),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_819),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_819),
.Y(n_1381)
);

CKINVDCx16_ASAP7_75t_R g1382 ( 
.A(n_1033),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_1077),
.Y(n_1383)
);

CKINVDCx20_ASAP7_75t_R g1384 ( 
.A(n_1085),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1086),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1087),
.B(n_1088),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1092),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_786),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1095),
.Y(n_1389)
);

INVxp67_ASAP7_75t_SL g1390 ( 
.A(n_911),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_824),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_R g1392 ( 
.A(n_1098),
.B(n_623),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_1099),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1101),
.Y(n_1394)
);

INVxp67_ASAP7_75t_SL g1395 ( 
.A(n_973),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_824),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1109),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_786),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_827),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_827),
.Y(n_1400)
);

INVxp33_ASAP7_75t_SL g1401 ( 
.A(n_787),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1110),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1115),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_828),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1118),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1121),
.B(n_485),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_828),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1124),
.Y(n_1408)
);

CKINVDCx16_ASAP7_75t_R g1409 ( 
.A(n_1033),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_829),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1135),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_832),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1136),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1137),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_1140),
.Y(n_1415)
);

INVxp33_ASAP7_75t_SL g1416 ( 
.A(n_1141),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_832),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1143),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1066),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_834),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_834),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_1066),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_835),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_835),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_836),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_803),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_836),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1130),
.B(n_485),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1081),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1130),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_838),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_844),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_1081),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1091),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_856),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_900),
.B(n_460),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_838),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_840),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_840),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_845),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_909),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_851),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_851),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_920),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_852),
.Y(n_1445)
);

INVxp67_ASAP7_75t_SL g1446 ( 
.A(n_1003),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1398),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1281),
.B(n_1100),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1398),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1145),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1153),
.B(n_1119),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1146),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1207),
.B(n_852),
.Y(n_1453)
);

INVx4_ASAP7_75t_L g1454 ( 
.A(n_1398),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1148),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1398),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1168),
.B(n_1201),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1152),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1154),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1289),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1289),
.Y(n_1461)
);

AND2x2_ASAP7_75t_SL g1462 ( 
.A(n_1311),
.B(n_603),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1432),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1232),
.B(n_783),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1156),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1161),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1398),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1367),
.B(n_1262),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1281),
.B(n_1091),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1378),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1252),
.B(n_853),
.Y(n_1471)
);

CKINVDCx16_ASAP7_75t_R g1472 ( 
.A(n_1360),
.Y(n_1472)
);

CKINVDCx6p67_ASAP7_75t_R g1473 ( 
.A(n_1342),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1223),
.A2(n_833),
.B1(n_782),
.B2(n_861),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1276),
.A2(n_965),
.B(n_957),
.Y(n_1475)
);

INVx4_ASAP7_75t_L g1476 ( 
.A(n_1378),
.Y(n_1476)
);

OA22x2_ASAP7_75t_SL g1477 ( 
.A1(n_1395),
.A2(n_661),
.B1(n_671),
.B2(n_653),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1296),
.A2(n_951),
.B1(n_1009),
.B2(n_897),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1163),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1374),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1148),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1426),
.B(n_906),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1204),
.Y(n_1483)
);

AND2x2_ASAP7_75t_SL g1484 ( 
.A(n_1242),
.B(n_723),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1252),
.B(n_853),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1272),
.B(n_783),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1164),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1204),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1214),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1167),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1378),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1294),
.B(n_783),
.Y(n_1492)
);

AOI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1369),
.A2(n_920),
.B1(n_627),
.B2(n_628),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1214),
.Y(n_1494)
);

OA21x2_ASAP7_75t_L g1495 ( 
.A1(n_1282),
.A2(n_965),
.B(n_957),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1277),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1388),
.Y(n_1497)
);

BUFx6f_ASAP7_75t_L g1498 ( 
.A(n_1388),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1285),
.A2(n_629),
.B1(n_637),
.B2(n_626),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1171),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1172),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1317),
.B(n_783),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1175),
.Y(n_1503)
);

INVx5_ASAP7_75t_L g1504 ( 
.A(n_1388),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1277),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1331),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1193),
.A2(n_644),
.B1(n_645),
.B2(n_639),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_SL g1508 ( 
.A1(n_1209),
.A2(n_932),
.B1(n_697),
.B2(n_638),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1176),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1194),
.A2(n_655),
.B1(n_657),
.B2(n_650),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1341),
.B(n_783),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1252),
.B(n_858),
.Y(n_1512)
);

INVx6_ASAP7_75t_L g1513 ( 
.A(n_1434),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1331),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1441),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1354),
.B(n_783),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1177),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1441),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1284),
.Y(n_1519)
);

INVx6_ASAP7_75t_L g1520 ( 
.A(n_1434),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1386),
.A2(n_662),
.B1(n_663),
.B2(n_660),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1426),
.B(n_959),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1179),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1226),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1430),
.B(n_1080),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1318),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_SL g1527 ( 
.A1(n_1196),
.A2(n_697),
.B1(n_681),
.B2(n_696),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1390),
.B(n_783),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1180),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1271),
.B(n_783),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1181),
.B(n_858),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1286),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1288),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1183),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1189),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1291),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1293),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1190),
.B(n_860),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1192),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_1330),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_SL g1541 ( 
.A1(n_1209),
.A2(n_718),
.B1(n_770),
.B2(n_674),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1227),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1298),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_L g1544 ( 
.A(n_1300),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1195),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1303),
.A2(n_980),
.B(n_971),
.Y(n_1546)
);

BUFx8_ASAP7_75t_SL g1547 ( 
.A(n_1301),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1430),
.B(n_1004),
.Y(n_1548)
);

INVx5_ASAP7_75t_L g1549 ( 
.A(n_1332),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1274),
.B(n_783),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_1304),
.Y(n_1551)
);

INVx6_ASAP7_75t_L g1552 ( 
.A(n_1332),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1227),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1305),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1198),
.Y(n_1555)
);

BUFx12f_ASAP7_75t_L g1556 ( 
.A(n_1301),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1315),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1319),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1323),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1206),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1208),
.B(n_859),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1324),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1406),
.B(n_1428),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_SL g1564 ( 
.A1(n_1287),
.A2(n_507),
.B1(n_611),
.B2(n_542),
.Y(n_1564)
);

CKINVDCx6p67_ASAP7_75t_R g1565 ( 
.A(n_1359),
.Y(n_1565)
);

XOR2xp5_ASAP7_75t_L g1566 ( 
.A(n_1309),
.B(n_665),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1213),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1328),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1336),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1225),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1446),
.B(n_842),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1238),
.B(n_1072),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1345),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1233),
.B(n_860),
.Y(n_1574)
);

OA21x2_ASAP7_75t_L g1575 ( 
.A1(n_1338),
.A2(n_980),
.B(n_971),
.Y(n_1575)
);

NOR2x1_ASAP7_75t_L g1576 ( 
.A(n_1362),
.B(n_500),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1234),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1236),
.Y(n_1578)
);

BUFx3_ASAP7_75t_L g1579 ( 
.A(n_1237),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1339),
.B(n_999),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1229),
.A2(n_1017),
.B(n_999),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1244),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1340),
.B(n_1017),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1248),
.B(n_864),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1250),
.B(n_859),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1363),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1365),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1253),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1343),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1344),
.B(n_1024),
.Y(n_1590)
);

OA21x2_ASAP7_75t_L g1591 ( 
.A1(n_1350),
.A2(n_1067),
.B(n_1024),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1355),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1392),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1254),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1259),
.Y(n_1595)
);

BUFx6f_ASAP7_75t_L g1596 ( 
.A(n_1356),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1357),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1358),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1229),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_L g1600 ( 
.A(n_1364),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1211),
.A2(n_667),
.B1(n_669),
.B2(n_664),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1444),
.Y(n_1602)
);

BUFx6f_ASAP7_75t_L g1603 ( 
.A(n_1366),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1235),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1371),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1260),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1264),
.B(n_863),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1185),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1275),
.B(n_863),
.Y(n_1609)
);

BUFx3_ASAP7_75t_L g1610 ( 
.A(n_1419),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1373),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1377),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1379),
.B(n_869),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1380),
.B(n_1068),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1381),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1391),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1240),
.B(n_468),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1224),
.B(n_1436),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1396),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1224),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1399),
.B(n_869),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1445),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1400),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1404),
.B(n_1068),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1313),
.A2(n_507),
.B1(n_611),
.B2(n_542),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_SL g1626 ( 
.A1(n_1255),
.A2(n_666),
.B1(n_715),
.B2(n_619),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1407),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1410),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1412),
.Y(n_1629)
);

NOR2x1_ASAP7_75t_L g1630 ( 
.A(n_1422),
.B(n_500),
.Y(n_1630)
);

AND2x2_ASAP7_75t_SL g1631 ( 
.A(n_1212),
.B(n_723),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1155),
.A2(n_672),
.B1(n_675),
.B2(n_670),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1444),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1436),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1256),
.A2(n_666),
.B1(n_715),
.B2(n_619),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1188),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1290),
.Y(n_1637)
);

AND2x2_ASAP7_75t_SL g1638 ( 
.A(n_1215),
.B(n_723),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1417),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1420),
.B(n_873),
.Y(n_1640)
);

BUFx6f_ASAP7_75t_L g1641 ( 
.A(n_1421),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1423),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1424),
.Y(n_1643)
);

INVx3_ASAP7_75t_L g1644 ( 
.A(n_1445),
.Y(n_1644)
);

OA21x2_ASAP7_75t_L g1645 ( 
.A1(n_1425),
.A2(n_1094),
.B(n_1074),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1158),
.A2(n_679),
.B1(n_680),
.B2(n_678),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1326),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1427),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1431),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1437),
.Y(n_1650)
);

OAI22x1_ASAP7_75t_R g1651 ( 
.A1(n_1267),
.A2(n_686),
.B1(n_688),
.B2(n_682),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1438),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_L g1653 ( 
.A(n_1439),
.Y(n_1653)
);

AND2x6_ASAP7_75t_L g1654 ( 
.A(n_1440),
.B(n_552),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1348),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1442),
.B(n_873),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1443),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1416),
.A2(n_694),
.B1(n_699),
.B2(n_693),
.Y(n_1658)
);

OAI21x1_ASAP7_75t_L g1659 ( 
.A1(n_1297),
.A2(n_890),
.B(n_888),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1361),
.A2(n_705),
.B1(n_707),
.B2(n_701),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1297),
.Y(n_1661)
);

BUFx6f_ASAP7_75t_L g1662 ( 
.A(n_1144),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1202),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1368),
.B(n_864),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1247),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1346),
.Y(n_1666)
);

INVx6_ASAP7_75t_L g1667 ( 
.A(n_1382),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1279),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1307),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1316),
.B(n_888),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1325),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1372),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1402),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1346),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1409),
.B(n_865),
.Y(n_1675)
);

INVx5_ASAP7_75t_L g1676 ( 
.A(n_1245),
.Y(n_1676)
);

AND2x6_ASAP7_75t_L g1677 ( 
.A(n_1346),
.B(n_552),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1144),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1147),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1416),
.B(n_1102),
.Y(n_1680)
);

AND2x6_ASAP7_75t_L g1681 ( 
.A(n_1200),
.B(n_552),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1147),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_1150),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1150),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1220),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1157),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1157),
.Y(n_1687)
);

INVx4_ASAP7_75t_L g1688 ( 
.A(n_1160),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1186),
.A2(n_894),
.B(n_890),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1327),
.B(n_1006),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1160),
.B(n_786),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1165),
.B(n_546),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1165),
.B(n_786),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1429),
.B(n_894),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1166),
.B(n_460),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1166),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1169),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1169),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1310),
.B(n_865),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1173),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1312),
.B(n_868),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1173),
.B(n_960),
.Y(n_1702)
);

BUFx2_ASAP7_75t_L g1703 ( 
.A(n_1435),
.Y(n_1703)
);

OAI21x1_ASAP7_75t_L g1704 ( 
.A1(n_1186),
.A2(n_585),
.B(n_583),
.Y(n_1704)
);

AOI22x1_ASAP7_75t_SL g1705 ( 
.A1(n_1435),
.A2(n_710),
.B1(n_712),
.B2(n_709),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1174),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1174),
.B(n_960),
.Y(n_1707)
);

OA21x2_ASAP7_75t_L g1708 ( 
.A1(n_1182),
.A2(n_870),
.B(n_868),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1182),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1184),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1258),
.A2(n_713),
.B1(n_716),
.B2(n_714),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1184),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1187),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1187),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1191),
.Y(n_1715)
);

INVx3_ASAP7_75t_L g1716 ( 
.A(n_1191),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1197),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1197),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1433),
.B(n_870),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1199),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1199),
.Y(n_1721)
);

INVx6_ASAP7_75t_L g1722 ( 
.A(n_1258),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1302),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1203),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1203),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1205),
.B(n_874),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1205),
.Y(n_1727)
);

NAND3xp33_ASAP7_75t_L g1728 ( 
.A(n_1302),
.B(n_726),
.C(n_724),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1210),
.A2(n_728),
.B1(n_731),
.B2(n_727),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1210),
.B(n_874),
.Y(n_1730)
);

INVx3_ASAP7_75t_L g1731 ( 
.A(n_1216),
.Y(n_1731)
);

BUFx8_ASAP7_75t_L g1732 ( 
.A(n_1353),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1216),
.B(n_960),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1468),
.B(n_1217),
.Y(n_1734)
);

OR2x6_ASAP7_75t_L g1735 ( 
.A(n_1667),
.B(n_1524),
.Y(n_1735)
);

INVxp33_ASAP7_75t_L g1736 ( 
.A(n_1480),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1457),
.B(n_1306),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1462),
.A2(n_1218),
.B1(n_1219),
.B2(n_1217),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1563),
.B(n_1306),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1620),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1522),
.B(n_1308),
.Y(n_1741)
);

OAI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1474),
.A2(n_1314),
.B1(n_1320),
.B2(n_1308),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1484),
.A2(n_1462),
.B1(n_1708),
.B2(n_1485),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1618),
.B(n_1314),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1514),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1484),
.A2(n_585),
.B1(n_599),
.B2(n_583),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1450),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1450),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1508),
.A2(n_1269),
.B1(n_1280),
.B2(n_1268),
.Y(n_1749)
);

OAI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1620),
.A2(n_1321),
.B1(n_1322),
.B2(n_1320),
.Y(n_1750)
);

OR2x6_ASAP7_75t_L g1751 ( 
.A(n_1667),
.B(n_1278),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1451),
.A2(n_1634),
.B1(n_1708),
.B2(n_1448),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1452),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1460),
.B(n_1006),
.Y(n_1754)
);

AND2x2_ASAP7_75t_SL g1755 ( 
.A(n_1631),
.B(n_661),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1618),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1708),
.A2(n_599),
.B1(n_640),
.B2(n_633),
.Y(n_1757)
);

BUFx10_ASAP7_75t_L g1758 ( 
.A(n_1680),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1460),
.B(n_1011),
.Y(n_1759)
);

AO22x2_ASAP7_75t_L g1760 ( 
.A1(n_1478),
.A2(n_743),
.B1(n_768),
.B2(n_764),
.Y(n_1760)
);

OAI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1634),
.A2(n_1322),
.B1(n_1329),
.B2(n_1321),
.Y(n_1761)
);

OAI22xp33_ASAP7_75t_SL g1762 ( 
.A1(n_1530),
.A2(n_633),
.B1(n_651),
.B2(n_640),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1525),
.B(n_1329),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1664),
.B(n_1334),
.Y(n_1764)
);

INVx3_ASAP7_75t_L g1765 ( 
.A(n_1561),
.Y(n_1765)
);

OAI22xp33_ASAP7_75t_SL g1766 ( 
.A1(n_1550),
.A2(n_651),
.B1(n_708),
.B2(n_700),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_1461),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1514),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1514),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1455),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_SL g1771 ( 
.A1(n_1541),
.A2(n_1151),
.B1(n_1159),
.B2(n_1149),
.Y(n_1771)
);

OAI22xp33_ASAP7_75t_SL g1772 ( 
.A1(n_1452),
.A2(n_1459),
.B1(n_1500),
.B2(n_1458),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1527),
.A2(n_1170),
.B1(n_1178),
.B2(n_1162),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_SL g1774 ( 
.A1(n_1626),
.A2(n_1228),
.B1(n_1249),
.B2(n_1231),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1548),
.B(n_1334),
.Y(n_1775)
);

OR2x6_ASAP7_75t_L g1776 ( 
.A(n_1667),
.B(n_591),
.Y(n_1776)
);

OAI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1493),
.A2(n_1337),
.B1(n_1347),
.B2(n_1335),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_SL g1778 ( 
.A1(n_1635),
.A2(n_1376),
.B1(n_1383),
.B2(n_1370),
.Y(n_1778)
);

AO22x2_ASAP7_75t_L g1779 ( 
.A1(n_1705),
.A2(n_743),
.B1(n_764),
.B2(n_591),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1471),
.A2(n_700),
.B1(n_766),
.B2(n_708),
.Y(n_1780)
);

AO22x2_ASAP7_75t_L g1781 ( 
.A1(n_1705),
.A2(n_743),
.B1(n_764),
.B2(n_591),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1458),
.Y(n_1782)
);

AOI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1471),
.A2(n_766),
.B1(n_768),
.B2(n_1335),
.Y(n_1783)
);

OAI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1690),
.A2(n_1347),
.B1(n_1349),
.B2(n_1337),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1664),
.B(n_1675),
.Y(n_1785)
);

OAI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1690),
.A2(n_1351),
.B1(n_1352),
.B2(n_1349),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1485),
.A2(n_768),
.B1(n_1352),
.B2(n_1351),
.Y(n_1787)
);

OAI22xp33_ASAP7_75t_SL g1788 ( 
.A1(n_1459),
.A2(n_690),
.B1(n_692),
.B2(n_671),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1455),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1675),
.B(n_1375),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1500),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1481),
.Y(n_1792)
);

AO22x2_ASAP7_75t_L g1793 ( 
.A1(n_1499),
.A2(n_1692),
.B1(n_1679),
.B2(n_1682),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1461),
.B(n_1011),
.Y(n_1794)
);

OAI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1571),
.A2(n_1385),
.B1(n_1387),
.B2(n_1375),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1512),
.B(n_1218),
.Y(n_1796)
);

OA22x2_ASAP7_75t_L g1797 ( 
.A1(n_1564),
.A2(n_1387),
.B1(n_1389),
.B2(n_1385),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1481),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1512),
.A2(n_1389),
.B1(n_1397),
.B2(n_1394),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1515),
.B(n_1394),
.Y(n_1800)
);

OAI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1521),
.A2(n_1405),
.B1(n_1408),
.B2(n_1397),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1469),
.B(n_1670),
.Y(n_1802)
);

INVx3_ASAP7_75t_L g1803 ( 
.A(n_1561),
.Y(n_1803)
);

AOI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1448),
.A2(n_1408),
.B1(n_1414),
.B2(n_1405),
.Y(n_1804)
);

BUFx6f_ASAP7_75t_SL g1805 ( 
.A(n_1610),
.Y(n_1805)
);

OAI22xp33_ASAP7_75t_SL g1806 ( 
.A1(n_1501),
.A2(n_692),
.B1(n_695),
.B2(n_690),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1483),
.Y(n_1807)
);

AOI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1631),
.A2(n_1418),
.B1(n_1414),
.B2(n_1393),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1638),
.A2(n_1418),
.B1(n_1403),
.B2(n_1411),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1515),
.B(n_1219),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1638),
.A2(n_1415),
.B1(n_1413),
.B2(n_1384),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1483),
.Y(n_1812)
);

AND2x4_ASAP7_75t_L g1813 ( 
.A(n_1469),
.B(n_1012),
.Y(n_1813)
);

OAI22xp5_ASAP7_75t_SL g1814 ( 
.A1(n_1625),
.A2(n_733),
.B1(n_734),
.B2(n_732),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1572),
.B(n_1221),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1699),
.B(n_1221),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1699),
.B(n_1222),
.Y(n_1817)
);

OA22x2_ASAP7_75t_L g1818 ( 
.A1(n_1646),
.A2(n_1230),
.B1(n_1239),
.B2(n_1222),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1488),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1469),
.B(n_1670),
.Y(n_1820)
);

OAI22xp33_ASAP7_75t_R g1821 ( 
.A1(n_1695),
.A2(n_706),
.B1(n_711),
.B2(n_695),
.Y(n_1821)
);

OR2x6_ASAP7_75t_L g1822 ( 
.A(n_1667),
.B(n_706),
.Y(n_1822)
);

AOI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1501),
.A2(n_1239),
.B1(n_1241),
.B2(n_1230),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1488),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1453),
.B(n_1241),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1503),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1701),
.B(n_1243),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1701),
.B(n_1463),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1489),
.Y(n_1829)
);

AO22x2_ASAP7_75t_L g1830 ( 
.A1(n_1678),
.A2(n_717),
.B1(n_719),
.B2(n_711),
.Y(n_1830)
);

AOI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1503),
.A2(n_1246),
.B1(n_1251),
.B2(n_1243),
.Y(n_1831)
);

OA22x2_ASAP7_75t_L g1832 ( 
.A1(n_1507),
.A2(n_1510),
.B1(n_1482),
.B2(n_1729),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1509),
.Y(n_1833)
);

INVx1_ASAP7_75t_SL g1834 ( 
.A(n_1540),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1726),
.B(n_1730),
.Y(n_1835)
);

OAI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1691),
.A2(n_1251),
.B1(n_1257),
.B2(n_1246),
.Y(n_1836)
);

AND2x4_ASAP7_75t_L g1837 ( 
.A(n_1670),
.B(n_1012),
.Y(n_1837)
);

AO22x2_ASAP7_75t_L g1838 ( 
.A1(n_1678),
.A2(n_719),
.B1(n_730),
.B2(n_717),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1509),
.B(n_1257),
.Y(n_1839)
);

OAI22xp33_ASAP7_75t_SL g1840 ( 
.A1(n_1517),
.A2(n_735),
.B1(n_737),
.B2(n_730),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1726),
.B(n_1261),
.Y(n_1841)
);

BUFx2_ASAP7_75t_L g1842 ( 
.A(n_1540),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1552),
.Y(n_1843)
);

OAI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1733),
.A2(n_1702),
.B1(n_1707),
.B2(n_1693),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1489),
.Y(n_1845)
);

AO22x2_ASAP7_75t_L g1846 ( 
.A1(n_1679),
.A2(n_737),
.B1(n_750),
.B2(n_735),
.Y(n_1846)
);

OAI22xp33_ASAP7_75t_SL g1847 ( 
.A1(n_1517),
.A2(n_752),
.B1(n_754),
.B2(n_750),
.Y(n_1847)
);

OAI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1523),
.A2(n_1263),
.B1(n_1265),
.B2(n_1261),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1494),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1494),
.Y(n_1850)
);

AOI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1523),
.A2(n_1265),
.B1(n_1266),
.B2(n_1263),
.Y(n_1851)
);

INVx5_ASAP7_75t_L g1852 ( 
.A(n_1677),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1637),
.B(n_1266),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1726),
.B(n_1730),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1529),
.A2(n_1273),
.B1(n_1283),
.B2(n_1270),
.Y(n_1855)
);

OAI22xp33_ASAP7_75t_R g1856 ( 
.A1(n_1651),
.A2(n_754),
.B1(n_758),
.B2(n_752),
.Y(n_1856)
);

OAI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1529),
.A2(n_1273),
.B1(n_1283),
.B2(n_1270),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1730),
.B(n_1292),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_SL g1859 ( 
.A1(n_1518),
.A2(n_741),
.B1(n_744),
.B2(n_736),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1637),
.B(n_1292),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1570),
.B(n_1577),
.Y(n_1861)
);

OA22x2_ASAP7_75t_L g1862 ( 
.A1(n_1658),
.A2(n_1299),
.B1(n_1295),
.B2(n_765),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1694),
.B(n_1295),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1694),
.B(n_1299),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1694),
.B(n_546),
.Y(n_1865)
);

OAI22xp33_ASAP7_75t_SL g1866 ( 
.A1(n_1534),
.A2(n_765),
.B1(n_758),
.B2(n_751),
.Y(n_1866)
);

AO22x2_ASAP7_75t_L g1867 ( 
.A1(n_1682),
.A2(n_1687),
.B1(n_1725),
.B2(n_1686),
.Y(n_1867)
);

OA22x2_ASAP7_75t_L g1868 ( 
.A1(n_1604),
.A2(n_1719),
.B1(n_1660),
.B2(n_1617),
.Y(n_1868)
);

OAI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1534),
.A2(n_1333),
.B1(n_756),
.B2(n_759),
.Y(n_1869)
);

AND2x2_ASAP7_75t_SL g1870 ( 
.A(n_1472),
.B(n_552),
.Y(n_1870)
);

AND2x6_ASAP7_75t_L g1871 ( 
.A(n_1666),
.B(n_1674),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1684),
.B(n_546),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1719),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1535),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1496),
.Y(n_1875)
);

OAI22xp33_ASAP7_75t_L g1876 ( 
.A1(n_1535),
.A2(n_1333),
.B1(n_761),
.B2(n_763),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1496),
.Y(n_1877)
);

OAI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1539),
.A2(n_767),
.B1(n_769),
.B2(n_745),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1719),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1570),
.B(n_1015),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1684),
.B(n_546),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1647),
.B(n_1353),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1666),
.A2(n_552),
.B1(n_773),
.B2(n_772),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1684),
.B(n_575),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1696),
.B(n_1710),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1539),
.A2(n_778),
.B1(n_779),
.B2(n_776),
.Y(n_1886)
);

AO22x2_ASAP7_75t_L g1887 ( 
.A1(n_1686),
.A2(n_1019),
.B1(n_1020),
.B2(n_1015),
.Y(n_1887)
);

AOI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1545),
.A2(n_1020),
.B1(n_1021),
.B2(n_1019),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1655),
.B(n_1593),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1696),
.B(n_575),
.Y(n_1890)
);

AOI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1545),
.A2(n_1595),
.B1(n_1585),
.B2(n_1561),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1505),
.Y(n_1892)
);

AO22x2_ASAP7_75t_L g1893 ( 
.A1(n_1687),
.A2(n_1022),
.B1(n_1027),
.B2(n_1021),
.Y(n_1893)
);

OAI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1595),
.A2(n_1401),
.B1(n_875),
.B2(n_878),
.Y(n_1894)
);

AOI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1585),
.A2(n_1027),
.B1(n_1028),
.B2(n_1022),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1505),
.Y(n_1896)
);

INVx2_ASAP7_75t_SL g1897 ( 
.A(n_1676),
.Y(n_1897)
);

OAI22xp33_ASAP7_75t_SL g1898 ( 
.A1(n_1465),
.A2(n_1029),
.B1(n_1030),
.B2(n_1028),
.Y(n_1898)
);

AOI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1585),
.A2(n_1030),
.B1(n_1036),
.B2(n_1029),
.Y(n_1899)
);

OAI22xp33_ASAP7_75t_SL g1900 ( 
.A1(n_1466),
.A2(n_1039),
.B1(n_1047),
.B2(n_1036),
.Y(n_1900)
);

OAI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1479),
.A2(n_1401),
.B1(n_875),
.B2(n_878),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1696),
.B(n_575),
.Y(n_1902)
);

AO22x2_ASAP7_75t_L g1903 ( 
.A1(n_1725),
.A2(n_1047),
.B1(n_1050),
.B2(n_1039),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1607),
.A2(n_1054),
.B1(n_1055),
.B2(n_1050),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1710),
.B(n_575),
.Y(n_1905)
);

OAI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1487),
.A2(n_879),
.B1(n_883),
.B2(n_876),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1506),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1710),
.B(n_742),
.Y(n_1908)
);

AOI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1607),
.A2(n_1056),
.B1(n_1058),
.B2(n_1055),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1716),
.B(n_742),
.Y(n_1910)
);

NAND2xp33_ASAP7_75t_SL g1911 ( 
.A(n_1593),
.B(n_1056),
.Y(n_1911)
);

AOI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1607),
.A2(n_1061),
.B1(n_1062),
.B2(n_1058),
.Y(n_1912)
);

INVx3_ASAP7_75t_L g1913 ( 
.A(n_1609),
.Y(n_1913)
);

OAI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1490),
.A2(n_879),
.B1(n_883),
.B2(n_876),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1716),
.B(n_742),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1609),
.A2(n_1062),
.B1(n_1063),
.B2(n_1061),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1609),
.A2(n_1065),
.B1(n_1069),
.B2(n_1063),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1716),
.B(n_742),
.Y(n_1918)
);

OAI22xp33_ASAP7_75t_SL g1919 ( 
.A1(n_1555),
.A2(n_1069),
.B1(n_1073),
.B2(n_1065),
.Y(n_1919)
);

AO22x2_ASAP7_75t_L g1920 ( 
.A1(n_1727),
.A2(n_1075),
.B1(n_1078),
.B2(n_1073),
.Y(n_1920)
);

AOI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1576),
.A2(n_1078),
.B1(n_1079),
.B2(n_1075),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1731),
.B(n_1079),
.Y(n_1922)
);

OR2x6_ASAP7_75t_L g1923 ( 
.A(n_1722),
.B(n_1082),
.Y(n_1923)
);

AND2x2_ASAP7_75t_SL g1924 ( 
.A(n_1703),
.B(n_1082),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1731),
.B(n_1518),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1506),
.Y(n_1926)
);

AO22x2_ASAP7_75t_L g1927 ( 
.A1(n_1727),
.A2(n_1084),
.B1(n_1089),
.B2(n_1083),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1613),
.Y(n_1928)
);

AOI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1531),
.A2(n_1084),
.B1(n_1089),
.B2(n_1083),
.Y(n_1929)
);

AO22x2_ASAP7_75t_L g1930 ( 
.A1(n_1601),
.A2(n_1093),
.B1(n_1096),
.B2(n_1090),
.Y(n_1930)
);

OA22x2_ASAP7_75t_L g1931 ( 
.A1(n_1663),
.A2(n_1093),
.B1(n_1096),
.B2(n_1090),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1613),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1531),
.Y(n_1933)
);

AND2x2_ASAP7_75t_SL g1934 ( 
.A(n_1602),
.B(n_1142),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1613),
.Y(n_1935)
);

AOI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1538),
.A2(n_1104),
.B1(n_1105),
.B2(n_1103),
.Y(n_1936)
);

OAI22xp33_ASAP7_75t_L g1937 ( 
.A1(n_1560),
.A2(n_884),
.B1(n_889),
.B2(n_887),
.Y(n_1937)
);

INVx3_ASAP7_75t_L g1938 ( 
.A(n_1621),
.Y(n_1938)
);

INVx8_ASAP7_75t_L g1939 ( 
.A(n_1676),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1731),
.B(n_1103),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1700),
.B(n_1104),
.Y(n_1941)
);

OAI22xp33_ASAP7_75t_L g1942 ( 
.A1(n_1567),
.A2(n_884),
.B1(n_889),
.B2(n_887),
.Y(n_1942)
);

AOI22x1_ASAP7_75t_L g1943 ( 
.A1(n_1542),
.A2(n_1106),
.B1(n_1107),
.B2(n_1105),
.Y(n_1943)
);

OAI22xp5_ASAP7_75t_SL g1944 ( 
.A1(n_1566),
.A2(n_1107),
.B1(n_1108),
.B2(n_1106),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1621),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1700),
.B(n_1108),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1706),
.B(n_1111),
.Y(n_1947)
);

AND2x4_ASAP7_75t_L g1948 ( 
.A(n_1577),
.B(n_1111),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1621),
.Y(n_1949)
);

AOI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1538),
.A2(n_1113),
.B1(n_1114),
.B2(n_1112),
.Y(n_1950)
);

AO22x2_ASAP7_75t_L g1951 ( 
.A1(n_1632),
.A2(n_1113),
.B1(n_1114),
.B2(n_1112),
.Y(n_1951)
);

BUFx2_ASAP7_75t_L g1952 ( 
.A(n_1587),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1706),
.B(n_1116),
.Y(n_1953)
);

OAI22xp33_ASAP7_75t_R g1954 ( 
.A1(n_1526),
.A2(n_1117),
.B1(n_1122),
.B2(n_1116),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1574),
.A2(n_1122),
.B1(n_1123),
.B2(n_1117),
.Y(n_1955)
);

OAI22xp33_ASAP7_75t_SL g1956 ( 
.A1(n_1578),
.A2(n_1125),
.B1(n_1127),
.B2(n_1123),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1713),
.B(n_1125),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1602),
.B(n_1127),
.Y(n_1958)
);

NAND2xp33_ASAP7_75t_SL g1959 ( 
.A(n_1662),
.B(n_1128),
.Y(n_1959)
);

AOI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1574),
.A2(n_1584),
.B1(n_1588),
.B2(n_1582),
.Y(n_1960)
);

AOI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1584),
.A2(n_1129),
.B1(n_1139),
.B2(n_1128),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1594),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1640),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1640),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1662),
.B(n_1129),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1713),
.B(n_1139),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1612),
.A2(n_1142),
.B1(n_892),
.B2(n_896),
.Y(n_1967)
);

AOI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1612),
.A2(n_892),
.B1(n_896),
.B2(n_895),
.Y(n_1968)
);

AOI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1616),
.A2(n_895),
.B1(n_899),
.B2(n_898),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1714),
.B(n_898),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1640),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1656),
.Y(n_1972)
);

BUFx10_ASAP7_75t_L g1973 ( 
.A(n_1662),
.Y(n_1973)
);

OAI22xp33_ASAP7_75t_L g1974 ( 
.A1(n_1579),
.A2(n_899),
.B1(n_904),
.B2(n_902),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1656),
.Y(n_1975)
);

AOI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1616),
.A2(n_902),
.B1(n_912),
.B2(n_904),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1656),
.Y(n_1977)
);

OAI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1674),
.A2(n_912),
.B1(n_914),
.B2(n_913),
.Y(n_1978)
);

AOI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1623),
.A2(n_913),
.B1(n_918),
.B2(n_914),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1714),
.B(n_918),
.Y(n_1980)
);

AND2x4_ASAP7_75t_L g1981 ( 
.A(n_1579),
.B(n_922),
.Y(n_1981)
);

XOR2xp5_ASAP7_75t_L g1982 ( 
.A(n_1608),
.B(n_305),
.Y(n_1982)
);

XNOR2xp5_ASAP7_75t_L g1983 ( 
.A(n_1587),
.B(n_306),
.Y(n_1983)
);

INVx2_ASAP7_75t_SL g1984 ( 
.A(n_1676),
.Y(n_1984)
);

OAI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1623),
.A2(n_922),
.B1(n_925),
.B2(n_924),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1720),
.B(n_924),
.Y(n_1986)
);

AOI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1627),
.A2(n_925),
.B1(n_936),
.B2(n_929),
.Y(n_1987)
);

INVx3_ASAP7_75t_L g1988 ( 
.A(n_1659),
.Y(n_1988)
);

INVx1_ASAP7_75t_SL g1989 ( 
.A(n_1633),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1606),
.Y(n_1990)
);

OAI22xp33_ASAP7_75t_SL g1991 ( 
.A1(n_1627),
.A2(n_936),
.B1(n_938),
.B2(n_929),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1533),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1720),
.B(n_1721),
.Y(n_1993)
);

OAI22xp33_ASAP7_75t_L g1994 ( 
.A1(n_1606),
.A2(n_938),
.B1(n_940),
.B2(n_939),
.Y(n_1994)
);

AOI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1628),
.A2(n_939),
.B1(n_943),
.B2(n_940),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1533),
.Y(n_1996)
);

CKINVDCx6p67_ASAP7_75t_R g1997 ( 
.A(n_1556),
.Y(n_1997)
);

INVx2_ASAP7_75t_SL g1998 ( 
.A(n_1676),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1721),
.B(n_943),
.Y(n_1999)
);

AO22x2_ASAP7_75t_L g2000 ( 
.A1(n_1698),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1663),
.B(n_944),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1665),
.B(n_944),
.Y(n_2002)
);

OAI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1665),
.A2(n_1668),
.B1(n_1671),
.B2(n_1669),
.Y(n_2003)
);

AOI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1628),
.A2(n_945),
.B1(n_961),
.B2(n_960),
.Y(n_2004)
);

XNOR2xp5_ASAP7_75t_L g2005 ( 
.A(n_1608),
.B(n_1636),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1668),
.B(n_945),
.Y(n_2006)
);

AOI22xp5_ASAP7_75t_SL g2007 ( 
.A1(n_1566),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_2007)
);

OAI22xp33_ASAP7_75t_SL g2008 ( 
.A1(n_1629),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_2008)
);

AO22x2_ASAP7_75t_L g2009 ( 
.A1(n_1709),
.A2(n_13),
.B1(n_9),
.B2(n_10),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1669),
.B(n_960),
.Y(n_2010)
);

OAI22xp33_ASAP7_75t_SL g2011 ( 
.A1(n_1629),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1536),
.Y(n_2012)
);

OAI22xp33_ASAP7_75t_SL g2013 ( 
.A1(n_1464),
.A2(n_19),
.B1(n_15),
.B2(n_17),
.Y(n_2013)
);

OA22x2_ASAP7_75t_L g2014 ( 
.A1(n_1671),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1661),
.Y(n_2015)
);

AOI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1639),
.A2(n_961),
.B1(n_1133),
.B2(n_1064),
.Y(n_2016)
);

OAI22xp33_ASAP7_75t_SL g2017 ( 
.A1(n_1486),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_2017)
);

OAI22xp33_ASAP7_75t_SL g2018 ( 
.A1(n_1492),
.A2(n_28),
.B1(n_24),
.B2(n_27),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1542),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1672),
.B(n_1133),
.Y(n_2020)
);

XOR2xp5_ASAP7_75t_L g2021 ( 
.A(n_1636),
.B(n_307),
.Y(n_2021)
);

AOI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1642),
.A2(n_961),
.B1(n_1133),
.B2(n_1064),
.Y(n_2022)
);

BUFx3_ASAP7_75t_L g2023 ( 
.A(n_1610),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_L g2024 ( 
.A(n_1711),
.B(n_24),
.Y(n_2024)
);

OAI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1643),
.A2(n_1657),
.B1(n_1648),
.B2(n_1672),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1536),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1502),
.B(n_1133),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1537),
.Y(n_2028)
);

NAND3x1_ASAP7_75t_L g2029 ( 
.A(n_1630),
.B(n_27),
.C(n_28),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1542),
.Y(n_2030)
);

INVxp67_ASAP7_75t_SL g2031 ( 
.A(n_1553),
.Y(n_2031)
);

INVx3_ASAP7_75t_L g2032 ( 
.A(n_2019),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1770),
.Y(n_2033)
);

BUFx6f_ASAP7_75t_L g2034 ( 
.A(n_1843),
.Y(n_2034)
);

INVx4_ASAP7_75t_SL g2035 ( 
.A(n_1871),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1789),
.Y(n_2036)
);

INVx3_ASAP7_75t_L g2037 ( 
.A(n_2030),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1792),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1798),
.Y(n_2039)
);

INVx4_ASAP7_75t_L g2040 ( 
.A(n_1843),
.Y(n_2040)
);

BUFx4f_ASAP7_75t_L g2041 ( 
.A(n_1939),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1922),
.B(n_1511),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1928),
.Y(n_2043)
);

BUFx10_ASAP7_75t_L g2044 ( 
.A(n_1889),
.Y(n_2044)
);

BUFx2_ASAP7_75t_L g2045 ( 
.A(n_1735),
.Y(n_2045)
);

AOI22xp33_ASAP7_75t_L g2046 ( 
.A1(n_1746),
.A2(n_1543),
.B1(n_1554),
.B2(n_1537),
.Y(n_2046)
);

INVx3_ASAP7_75t_L g2047 ( 
.A(n_1765),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1932),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1935),
.Y(n_2049)
);

INVx3_ASAP7_75t_L g2050 ( 
.A(n_1765),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_SL g2051 ( 
.A(n_1835),
.B(n_1662),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1807),
.Y(n_2052)
);

OR2x6_ASAP7_75t_L g2053 ( 
.A(n_1854),
.B(n_1662),
.Y(n_2053)
);

AOI22xp33_ASAP7_75t_L g2054 ( 
.A1(n_1746),
.A2(n_1554),
.B1(n_1558),
.B2(n_1543),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1940),
.B(n_1683),
.Y(n_2055)
);

BUFx3_ASAP7_75t_L g2056 ( 
.A(n_1973),
.Y(n_2056)
);

BUFx2_ASAP7_75t_L g2057 ( 
.A(n_1735),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1945),
.Y(n_2058)
);

INVx5_ASAP7_75t_L g2059 ( 
.A(n_1852),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1812),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1819),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_1885),
.B(n_1683),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1824),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1829),
.Y(n_2064)
);

OR2x6_ASAP7_75t_L g2065 ( 
.A(n_1939),
.B(n_1683),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1845),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1849),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1739),
.B(n_1516),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1850),
.Y(n_2069)
);

BUFx3_ASAP7_75t_L g2070 ( 
.A(n_1973),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1941),
.B(n_1683),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1875),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1877),
.Y(n_2073)
);

INVxp33_ASAP7_75t_L g2074 ( 
.A(n_1828),
.Y(n_2074)
);

OAI22xp5_ASAP7_75t_L g2075 ( 
.A1(n_1743),
.A2(n_1712),
.B1(n_1673),
.B2(n_1722),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1892),
.Y(n_2076)
);

NOR2x1p5_ASAP7_75t_L g2077 ( 
.A(n_1997),
.B(n_1473),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1896),
.Y(n_2078)
);

XOR2xp5_ASAP7_75t_L g2079 ( 
.A(n_2005),
.B(n_1749),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1907),
.Y(n_2080)
);

INVxp33_ASAP7_75t_SL g2081 ( 
.A(n_1771),
.Y(n_2081)
);

BUFx6f_ASAP7_75t_L g2082 ( 
.A(n_1843),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1926),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1734),
.B(n_1528),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_2015),
.Y(n_2085)
);

INVx3_ASAP7_75t_L g2086 ( 
.A(n_1803),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_1805),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1752),
.B(n_1553),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1803),
.Y(n_2089)
);

NOR2x1p5_ASAP7_75t_L g2090 ( 
.A(n_1853),
.B(n_1473),
.Y(n_2090)
);

AO22x2_ASAP7_75t_L g2091 ( 
.A1(n_1738),
.A2(n_1477),
.B1(n_1673),
.B2(n_1688),
.Y(n_2091)
);

NOR2xp33_ASAP7_75t_L g2092 ( 
.A(n_1737),
.B(n_1688),
.Y(n_2092)
);

INVx3_ASAP7_75t_L g2093 ( 
.A(n_1913),
.Y(n_2093)
);

NAND2xp33_ASAP7_75t_SL g2094 ( 
.A(n_1993),
.B(n_1683),
.Y(n_2094)
);

AND3x2_ASAP7_75t_L g2095 ( 
.A(n_2024),
.B(n_1633),
.C(n_1723),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1988),
.Y(n_2096)
);

BUFx6f_ASAP7_75t_L g2097 ( 
.A(n_1939),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1988),
.Y(n_2098)
);

NAND2xp33_ASAP7_75t_SL g2099 ( 
.A(n_1841),
.B(n_1697),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1913),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1938),
.Y(n_2101)
);

OAI22xp33_ASAP7_75t_L g2102 ( 
.A1(n_1743),
.A2(n_1697),
.B1(n_1717),
.B2(n_1715),
.Y(n_2102)
);

HB1xp67_ASAP7_75t_L g2103 ( 
.A(n_1740),
.Y(n_2103)
);

INVx4_ASAP7_75t_L g2104 ( 
.A(n_1767),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1938),
.Y(n_2105)
);

BUFx6f_ASAP7_75t_L g2106 ( 
.A(n_1852),
.Y(n_2106)
);

HB1xp67_ASAP7_75t_L g2107 ( 
.A(n_1785),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_1805),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1949),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_1946),
.B(n_1697),
.Y(n_2110)
);

OR2x2_ASAP7_75t_L g2111 ( 
.A(n_1756),
.B(n_1573),
.Y(n_2111)
);

BUFx6f_ASAP7_75t_L g2112 ( 
.A(n_1852),
.Y(n_2112)
);

INVx2_ASAP7_75t_SL g2113 ( 
.A(n_1947),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1977),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1963),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1964),
.Y(n_2116)
);

OR2x2_ASAP7_75t_L g2117 ( 
.A(n_1756),
.B(n_1586),
.Y(n_2117)
);

BUFx10_ASAP7_75t_L g2118 ( 
.A(n_1741),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_SL g2119 ( 
.A(n_1924),
.B(n_1697),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1971),
.Y(n_2120)
);

AND2x2_ASAP7_75t_SL g2121 ( 
.A(n_1755),
.B(n_1715),
.Y(n_2121)
);

INVx2_ASAP7_75t_SL g2122 ( 
.A(n_1953),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1972),
.Y(n_2123)
);

BUFx6f_ASAP7_75t_L g2124 ( 
.A(n_1802),
.Y(n_2124)
);

AOI22xp33_ASAP7_75t_L g2125 ( 
.A1(n_1832),
.A2(n_1558),
.B1(n_1562),
.B2(n_1559),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1747),
.B(n_1553),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_L g2127 ( 
.A(n_1775),
.B(n_1688),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_L g2128 ( 
.A(n_1796),
.B(n_1715),
.Y(n_2128)
);

AOI22xp33_ASAP7_75t_L g2129 ( 
.A1(n_1933),
.A2(n_1977),
.B1(n_1813),
.B2(n_1753),
.Y(n_2129)
);

INVx4_ASAP7_75t_L g2130 ( 
.A(n_1767),
.Y(n_2130)
);

INVx3_ASAP7_75t_L g2131 ( 
.A(n_1975),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_SL g2132 ( 
.A(n_1934),
.B(n_1715),
.Y(n_2132)
);

NOR2xp33_ASAP7_75t_L g2133 ( 
.A(n_1825),
.B(n_1715),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1748),
.B(n_1599),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1782),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1791),
.B(n_1599),
.Y(n_2136)
);

INVx2_ASAP7_75t_SL g2137 ( 
.A(n_1957),
.Y(n_2137)
);

INVx4_ASAP7_75t_L g2138 ( 
.A(n_1767),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2031),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1992),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1996),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2012),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_1771),
.Y(n_2143)
);

AOI22xp33_ASAP7_75t_L g2144 ( 
.A1(n_1813),
.A2(n_1833),
.B1(n_1874),
.B2(n_1826),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1966),
.B(n_1599),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_2026),
.Y(n_2146)
);

INVx4_ASAP7_75t_L g2147 ( 
.A(n_1802),
.Y(n_2147)
);

AND3x2_ASAP7_75t_L g2148 ( 
.A(n_1952),
.B(n_1547),
.C(n_1732),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2028),
.Y(n_2149)
);

NAND3xp33_ASAP7_75t_L g2150 ( 
.A(n_1804),
.B(n_1728),
.C(n_1718),
.Y(n_2150)
);

INVx3_ASAP7_75t_L g2151 ( 
.A(n_1820),
.Y(n_2151)
);

BUFx3_ASAP7_75t_L g2152 ( 
.A(n_1735),
.Y(n_2152)
);

INVx3_ASAP7_75t_L g2153 ( 
.A(n_1820),
.Y(n_2153)
);

NOR2xp33_ASAP7_75t_L g2154 ( 
.A(n_1815),
.B(n_1717),
.Y(n_2154)
);

INVx3_ASAP7_75t_L g2155 ( 
.A(n_1745),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1768),
.Y(n_2156)
);

AND2x6_ASAP7_75t_L g2157 ( 
.A(n_1757),
.B(n_1717),
.Y(n_2157)
);

AOI22xp33_ASAP7_75t_L g2158 ( 
.A1(n_1962),
.A2(n_1562),
.B1(n_1569),
.B2(n_1559),
.Y(n_2158)
);

INVx4_ASAP7_75t_L g2159 ( 
.A(n_1861),
.Y(n_2159)
);

BUFx2_ASAP7_75t_L g2160 ( 
.A(n_1873),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_SL g2161 ( 
.A(n_1804),
.B(n_1717),
.Y(n_2161)
);

NAND3xp33_ASAP7_75t_L g2162 ( 
.A(n_1882),
.B(n_1718),
.C(n_1717),
.Y(n_2162)
);

BUFx6f_ASAP7_75t_SL g2163 ( 
.A(n_1751),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1769),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_1970),
.B(n_1980),
.Y(n_2165)
);

BUFx4f_ASAP7_75t_L g2166 ( 
.A(n_1871),
.Y(n_2166)
);

INVx4_ASAP7_75t_L g2167 ( 
.A(n_1861),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1981),
.Y(n_2168)
);

INVxp67_ASAP7_75t_SL g2169 ( 
.A(n_1990),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1772),
.Y(n_2170)
);

NOR2x1p5_ASAP7_75t_L g2171 ( 
.A(n_1860),
.B(n_1565),
.Y(n_2171)
);

INVx3_ASAP7_75t_L g2172 ( 
.A(n_1981),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1880),
.Y(n_2173)
);

OR2x2_ASAP7_75t_L g2174 ( 
.A(n_1958),
.B(n_1565),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1880),
.Y(n_2175)
);

AND2x6_ASAP7_75t_L g2176 ( 
.A(n_1757),
.B(n_1718),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1986),
.B(n_1622),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1948),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1948),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1943),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1754),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1999),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_1799),
.B(n_1718),
.Y(n_2183)
);

NOR2xp33_ASAP7_75t_L g2184 ( 
.A(n_1763),
.B(n_1718),
.Y(n_2184)
);

BUFx10_ASAP7_75t_L g2185 ( 
.A(n_1870),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1837),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_SL g2187 ( 
.A(n_1799),
.B(n_1724),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1837),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1872),
.B(n_1622),
.Y(n_2189)
);

BUFx6f_ASAP7_75t_SL g2190 ( 
.A(n_1751),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1754),
.Y(n_2191)
);

NAND2xp33_ASAP7_75t_R g2192 ( 
.A(n_1800),
.B(n_1685),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2010),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2020),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_1839),
.B(n_1724),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1759),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2027),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1759),
.Y(n_2198)
);

NOR2xp33_ASAP7_75t_L g2199 ( 
.A(n_1736),
.B(n_1724),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1794),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2001),
.B(n_1724),
.Y(n_2201)
);

INVx4_ASAP7_75t_L g2202 ( 
.A(n_1923),
.Y(n_2202)
);

HAxp5_ASAP7_75t_SL g2203 ( 
.A(n_1809),
.B(n_1685),
.CON(n_2203),
.SN(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2002),
.B(n_1724),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1881),
.B(n_1622),
.Y(n_2205)
);

AOI22xp5_ASAP7_75t_L g2206 ( 
.A1(n_1744),
.A2(n_1520),
.B1(n_1513),
.B2(n_1552),
.Y(n_2206)
);

HB1xp67_ASAP7_75t_L g2207 ( 
.A(n_1879),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1884),
.B(n_1644),
.Y(n_2208)
);

OAI21xp5_ASAP7_75t_L g2209 ( 
.A1(n_1891),
.A2(n_1689),
.B(n_1704),
.Y(n_2209)
);

BUFx6f_ASAP7_75t_L g2210 ( 
.A(n_1871),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2006),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1890),
.B(n_1644),
.Y(n_2212)
);

AOI22xp5_ASAP7_75t_L g2213 ( 
.A1(n_1764),
.A2(n_1520),
.B1(n_1513),
.B2(n_1552),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_SL g2214 ( 
.A(n_1823),
.B(n_1676),
.Y(n_2214)
);

NOR2xp33_ASAP7_75t_L g2215 ( 
.A(n_1758),
.B(n_1790),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1902),
.B(n_1905),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1908),
.B(n_1644),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_1823),
.B(n_1549),
.Y(n_2218)
);

AOI22xp33_ASAP7_75t_L g2219 ( 
.A1(n_1762),
.A2(n_1589),
.B1(n_1592),
.B2(n_1569),
.Y(n_2219)
);

NOR2xp33_ASAP7_75t_L g2220 ( 
.A(n_1758),
.B(n_1722),
.Y(n_2220)
);

BUFx3_ASAP7_75t_L g2221 ( 
.A(n_2023),
.Y(n_2221)
);

INVxp67_ASAP7_75t_SL g2222 ( 
.A(n_1891),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_1910),
.B(n_1589),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_1915),
.B(n_1918),
.Y(n_2224)
);

AOI22xp33_ASAP7_75t_L g2225 ( 
.A1(n_1762),
.A2(n_1597),
.B1(n_1598),
.B2(n_1592),
.Y(n_2225)
);

BUFx4f_ASAP7_75t_L g2226 ( 
.A(n_1923),
.Y(n_2226)
);

INVx3_ASAP7_75t_L g2227 ( 
.A(n_1794),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_SL g2228 ( 
.A(n_1831),
.B(n_1549),
.Y(n_2228)
);

INVxp67_ASAP7_75t_L g2229 ( 
.A(n_1816),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1923),
.B(n_1704),
.Y(n_2230)
);

AOI22xp33_ASAP7_75t_L g2231 ( 
.A1(n_1766),
.A2(n_1598),
.B1(n_1605),
.B2(n_1597),
.Y(n_2231)
);

AOI22xp5_ASAP7_75t_L g2232 ( 
.A1(n_1858),
.A2(n_1520),
.B1(n_1513),
.B2(n_1552),
.Y(n_2232)
);

BUFx10_ASAP7_75t_L g2233 ( 
.A(n_1751),
.Y(n_2233)
);

NOR2xp33_ASAP7_75t_L g2234 ( 
.A(n_1795),
.B(n_1722),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_SL g2235 ( 
.A(n_1831),
.B(n_1549),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_1851),
.B(n_1549),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1772),
.B(n_1605),
.Y(n_2237)
);

INVx6_ASAP7_75t_L g2238 ( 
.A(n_1822),
.Y(n_2238)
);

AND2x4_ASAP7_75t_L g2239 ( 
.A(n_1897),
.B(n_1984),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1991),
.Y(n_2240)
);

INVx2_ASAP7_75t_SL g2241 ( 
.A(n_1965),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1960),
.B(n_1611),
.Y(n_2242)
);

INVx3_ASAP7_75t_L g2243 ( 
.A(n_1931),
.Y(n_2243)
);

NOR2x1p5_ASAP7_75t_L g2244 ( 
.A(n_1817),
.B(n_1556),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1991),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_1827),
.B(n_1513),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1960),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1985),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1887),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_1887),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_SL g2251 ( 
.A(n_1851),
.B(n_1549),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_1844),
.B(n_1611),
.Y(n_2252)
);

INVxp67_ASAP7_75t_L g2253 ( 
.A(n_1865),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1893),
.Y(n_2254)
);

INVx8_ASAP7_75t_L g2255 ( 
.A(n_1822),
.Y(n_2255)
);

BUFx10_ASAP7_75t_L g2256 ( 
.A(n_1998),
.Y(n_2256)
);

CKINVDCx20_ASAP7_75t_R g2257 ( 
.A(n_1749),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1968),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1893),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1903),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_L g2261 ( 
.A(n_1784),
.B(n_1520),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_1783),
.B(n_1619),
.Y(n_2262)
);

INVx1_ASAP7_75t_SL g2263 ( 
.A(n_1989),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1968),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1903),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1969),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_1920),
.B(n_1689),
.Y(n_2267)
);

INVx3_ASAP7_75t_L g2268 ( 
.A(n_1868),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1969),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2025),
.Y(n_2270)
);

AOI22xp5_ASAP7_75t_L g2271 ( 
.A1(n_1793),
.A2(n_1649),
.B1(n_1619),
.B2(n_1532),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1920),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1927),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_1783),
.B(n_1649),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1927),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_SL g2276 ( 
.A(n_1855),
.B(n_1786),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1930),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_1793),
.B(n_1519),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1930),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1951),
.Y(n_2280)
);

INVx2_ASAP7_75t_SL g2281 ( 
.A(n_1863),
.Y(n_2281)
);

BUFx6f_ASAP7_75t_L g2282 ( 
.A(n_1822),
.Y(n_2282)
);

INVx4_ASAP7_75t_L g2283 ( 
.A(n_1776),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_SL g2284 ( 
.A(n_1855),
.B(n_1750),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1951),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2014),
.Y(n_2286)
);

INVx2_ASAP7_75t_SL g2287 ( 
.A(n_1864),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_1976),
.Y(n_2288)
);

BUFx3_ASAP7_75t_L g2289 ( 
.A(n_1842),
.Y(n_2289)
);

INVx5_ASAP7_75t_L g2290 ( 
.A(n_1776),
.Y(n_2290)
);

BUFx3_ASAP7_75t_L g2291 ( 
.A(n_1925),
.Y(n_2291)
);

INVx3_ASAP7_75t_L g2292 ( 
.A(n_2029),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_SL g2293 ( 
.A(n_1761),
.B(n_1732),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1780),
.B(n_1519),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1978),
.Y(n_2295)
);

BUFx3_ASAP7_75t_L g2296 ( 
.A(n_1810),
.Y(n_2296)
);

INVx2_ASAP7_75t_SL g2297 ( 
.A(n_1867),
.Y(n_2297)
);

CKINVDCx11_ASAP7_75t_R g2298 ( 
.A(n_1834),
.Y(n_2298)
);

INVx3_ASAP7_75t_L g2299 ( 
.A(n_1776),
.Y(n_2299)
);

AND2x4_ASAP7_75t_L g2300 ( 
.A(n_1780),
.B(n_1476),
.Y(n_2300)
);

INVxp67_ASAP7_75t_SL g2301 ( 
.A(n_2003),
.Y(n_2301)
);

AOI22xp33_ASAP7_75t_L g2302 ( 
.A1(n_1766),
.A2(n_1532),
.B1(n_1544),
.B2(n_1519),
.Y(n_2302)
);

NAND3xp33_ASAP7_75t_SL g2303 ( 
.A(n_1808),
.B(n_1809),
.C(n_1811),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_1787),
.B(n_1519),
.Y(n_2304)
);

BUFx6f_ASAP7_75t_L g2305 ( 
.A(n_1959),
.Y(n_2305)
);

INVx3_ASAP7_75t_L g2306 ( 
.A(n_1867),
.Y(n_2306)
);

INVx4_ASAP7_75t_L g2307 ( 
.A(n_2000),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_1848),
.B(n_1732),
.Y(n_2308)
);

AOI22xp33_ASAP7_75t_SL g2309 ( 
.A1(n_1944),
.A2(n_1681),
.B1(n_1677),
.B2(n_1532),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_1787),
.B(n_1519),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1976),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1979),
.Y(n_2312)
);

BUFx3_ASAP7_75t_L g2313 ( 
.A(n_1834),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_1836),
.B(n_1532),
.Y(n_2314)
);

OA22x2_ASAP7_75t_L g2315 ( 
.A1(n_1814),
.A2(n_1944),
.B1(n_1808),
.B2(n_1859),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_1895),
.B(n_1476),
.Y(n_2316)
);

AOI22xp33_ASAP7_75t_L g2317 ( 
.A1(n_1862),
.A2(n_1544),
.B1(n_1551),
.B2(n_1532),
.Y(n_2317)
);

AOI22xp5_ASAP7_75t_L g2318 ( 
.A1(n_1911),
.A2(n_1551),
.B1(n_1557),
.B2(n_1544),
.Y(n_2318)
);

AOI22xp33_ASAP7_75t_L g2319 ( 
.A1(n_1760),
.A2(n_1551),
.B1(n_1557),
.B2(n_1544),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_L g2320 ( 
.A(n_1857),
.B(n_1547),
.Y(n_2320)
);

NAND3xp33_ASAP7_75t_L g2321 ( 
.A(n_1886),
.B(n_1583),
.C(n_1580),
.Y(n_2321)
);

INVxp67_ASAP7_75t_SL g2322 ( 
.A(n_2004),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1979),
.Y(n_2323)
);

INVx3_ASAP7_75t_L g2324 ( 
.A(n_2034),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_SL g2325 ( 
.A(n_2121),
.B(n_1801),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2107),
.B(n_1811),
.Y(n_2326)
);

BUFx3_ASAP7_75t_L g2327 ( 
.A(n_2221),
.Y(n_2327)
);

AOI22xp33_ASAP7_75t_L g2328 ( 
.A1(n_2315),
.A2(n_1821),
.B1(n_2013),
.B2(n_2017),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2165),
.B(n_1760),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2096),
.Y(n_2330)
);

BUFx6f_ASAP7_75t_L g2331 ( 
.A(n_2097),
.Y(n_2331)
);

AND2x4_ASAP7_75t_L g2332 ( 
.A(n_2159),
.B(n_1895),
.Y(n_2332)
);

INVxp67_ASAP7_75t_L g2333 ( 
.A(n_2111),
.Y(n_2333)
);

AND2x6_ASAP7_75t_L g2334 ( 
.A(n_2267),
.B(n_2004),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2096),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2098),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2085),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_SL g2338 ( 
.A(n_2121),
.B(n_1777),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2211),
.B(n_1886),
.Y(n_2339)
);

OR2x6_ASAP7_75t_L g2340 ( 
.A(n_2255),
.B(n_1778),
.Y(n_2340)
);

OR2x2_ASAP7_75t_SL g2341 ( 
.A(n_2303),
.B(n_1856),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2085),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2135),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2038),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_L g2345 ( 
.A(n_2074),
.B(n_1742),
.Y(n_2345)
);

AND2x4_ASAP7_75t_L g2346 ( 
.A(n_2159),
.B(n_1899),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2165),
.B(n_1894),
.Y(n_2347)
);

NOR2xp33_ASAP7_75t_L g2348 ( 
.A(n_2074),
.B(n_1773),
.Y(n_2348)
);

BUFx6f_ASAP7_75t_L g2349 ( 
.A(n_2097),
.Y(n_2349)
);

CKINVDCx5p33_ASAP7_75t_R g2350 ( 
.A(n_2192),
.Y(n_2350)
);

NOR2xp33_ASAP7_75t_L g2351 ( 
.A(n_2229),
.B(n_1773),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2133),
.B(n_1866),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2068),
.B(n_1866),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2098),
.Y(n_2354)
);

NOR2xp33_ASAP7_75t_L g2355 ( 
.A(n_2092),
.B(n_2127),
.Y(n_2355)
);

INVx2_ASAP7_75t_SL g2356 ( 
.A(n_2313),
.Y(n_2356)
);

AO22x2_ASAP7_75t_L g2357 ( 
.A1(n_2307),
.A2(n_2009),
.B1(n_2000),
.B2(n_2007),
.Y(n_2357)
);

BUFx6f_ASAP7_75t_L g2358 ( 
.A(n_2097),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2039),
.Y(n_2359)
);

BUFx2_ASAP7_75t_L g2360 ( 
.A(n_2289),
.Y(n_2360)
);

CKINVDCx20_ASAP7_75t_R g2361 ( 
.A(n_2298),
.Y(n_2361)
);

INVx3_ASAP7_75t_L g2362 ( 
.A(n_2034),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2063),
.Y(n_2363)
);

INVx3_ASAP7_75t_L g2364 ( 
.A(n_2034),
.Y(n_2364)
);

INVx3_ASAP7_75t_L g2365 ( 
.A(n_2034),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2063),
.Y(n_2366)
);

AOI22xp5_ASAP7_75t_L g2367 ( 
.A1(n_2154),
.A2(n_1818),
.B1(n_1797),
.B2(n_1954),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2033),
.Y(n_2368)
);

BUFx6f_ASAP7_75t_L g2369 ( 
.A(n_2097),
.Y(n_2369)
);

AND2x6_ASAP7_75t_L g2370 ( 
.A(n_2267),
.B(n_2016),
.Y(n_2370)
);

INVxp67_ASAP7_75t_L g2371 ( 
.A(n_2111),
.Y(n_2371)
);

INVx4_ASAP7_75t_SL g2372 ( 
.A(n_2157),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2064),
.Y(n_2373)
);

AND2x4_ASAP7_75t_L g2374 ( 
.A(n_2159),
.B(n_1899),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2066),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2066),
.Y(n_2376)
);

NOR2xp33_ASAP7_75t_L g2377 ( 
.A(n_2117),
.B(n_1901),
.Y(n_2377)
);

INVx8_ASAP7_75t_L g2378 ( 
.A(n_2255),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_2097),
.Y(n_2379)
);

AND2x4_ASAP7_75t_L g2380 ( 
.A(n_2167),
.B(n_1904),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2067),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2211),
.B(n_1830),
.Y(n_2382)
);

OAI221xp5_ASAP7_75t_L g2383 ( 
.A1(n_2276),
.A2(n_1814),
.B1(n_1859),
.B2(n_2007),
.C(n_1774),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2067),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2078),
.Y(n_2385)
);

INVx4_ASAP7_75t_L g2386 ( 
.A(n_2056),
.Y(n_2386)
);

BUFx2_ASAP7_75t_L g2387 ( 
.A(n_2289),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2078),
.Y(n_2388)
);

BUFx2_ASAP7_75t_L g2389 ( 
.A(n_2296),
.Y(n_2389)
);

HB1xp67_ASAP7_75t_L g2390 ( 
.A(n_2071),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2084),
.B(n_1869),
.Y(n_2391)
);

AO22x2_ASAP7_75t_L g2392 ( 
.A1(n_2307),
.A2(n_2009),
.B1(n_2021),
.B2(n_1982),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2080),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2080),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2036),
.Y(n_2395)
);

AND3x4_ASAP7_75t_L g2396 ( 
.A(n_2296),
.B(n_1774),
.C(n_1778),
.Y(n_2396)
);

AND2x4_ASAP7_75t_L g2397 ( 
.A(n_2167),
.B(n_1904),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2201),
.B(n_1830),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2036),
.Y(n_2399)
);

HB1xp67_ASAP7_75t_L g2400 ( 
.A(n_2071),
.Y(n_2400)
);

NAND3xp33_ASAP7_75t_SL g2401 ( 
.A(n_2184),
.B(n_1921),
.C(n_1883),
.Y(n_2401)
);

BUFx3_ASAP7_75t_L g2402 ( 
.A(n_2221),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2182),
.B(n_1876),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_L g2404 ( 
.A(n_2117),
.B(n_1878),
.Y(n_2404)
);

NAND2x1p5_ASAP7_75t_L g2405 ( 
.A(n_2166),
.B(n_1476),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2182),
.B(n_1788),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2052),
.Y(n_2407)
);

OR2x2_ASAP7_75t_L g2408 ( 
.A(n_2263),
.B(n_1983),
.Y(n_2408)
);

INVx3_ASAP7_75t_L g2409 ( 
.A(n_2082),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2083),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2083),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2216),
.B(n_1788),
.Y(n_2412)
);

OA22x2_ASAP7_75t_L g2413 ( 
.A1(n_2307),
.A2(n_2284),
.B1(n_2143),
.B2(n_2095),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2043),
.Y(n_2414)
);

BUFx6f_ASAP7_75t_L g2415 ( 
.A(n_2210),
.Y(n_2415)
);

BUFx6f_ASAP7_75t_L g2416 ( 
.A(n_2210),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2052),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2224),
.B(n_1806),
.Y(n_2418)
);

BUFx6f_ASAP7_75t_L g2419 ( 
.A(n_2210),
.Y(n_2419)
);

NOR2xp33_ASAP7_75t_L g2420 ( 
.A(n_2301),
.B(n_1806),
.Y(n_2420)
);

INVx3_ASAP7_75t_L g2421 ( 
.A(n_2082),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2055),
.B(n_1840),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2201),
.B(n_1838),
.Y(n_2423)
);

BUFx3_ASAP7_75t_L g2424 ( 
.A(n_2152),
.Y(n_2424)
);

OR2x2_ASAP7_75t_SL g2425 ( 
.A(n_2150),
.B(n_1779),
.Y(n_2425)
);

BUFx6f_ASAP7_75t_L g2426 ( 
.A(n_2210),
.Y(n_2426)
);

CKINVDCx20_ASAP7_75t_R g2427 ( 
.A(n_2298),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2055),
.B(n_1840),
.Y(n_2428)
);

HB1xp67_ASAP7_75t_L g2429 ( 
.A(n_2110),
.Y(n_2429)
);

NAND3x1_ASAP7_75t_L g2430 ( 
.A(n_2320),
.B(n_1936),
.C(n_1929),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2060),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2060),
.Y(n_2432)
);

AOI22xp33_ASAP7_75t_L g2433 ( 
.A1(n_2315),
.A2(n_2013),
.B1(n_2018),
.B2(n_2017),
.Y(n_2433)
);

BUFx2_ASAP7_75t_L g2434 ( 
.A(n_2045),
.Y(n_2434)
);

BUFx2_ASAP7_75t_L g2435 ( 
.A(n_2045),
.Y(n_2435)
);

BUFx6f_ASAP7_75t_L g2436 ( 
.A(n_2210),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2048),
.Y(n_2437)
);

BUFx3_ASAP7_75t_L g2438 ( 
.A(n_2152),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2049),
.Y(n_2439)
);

BUFx3_ASAP7_75t_L g2440 ( 
.A(n_2057),
.Y(n_2440)
);

AND2x6_ASAP7_75t_L g2441 ( 
.A(n_2300),
.B(n_2016),
.Y(n_2441)
);

INVxp67_ASAP7_75t_L g2442 ( 
.A(n_2204),
.Y(n_2442)
);

AND2x2_ASAP7_75t_L g2443 ( 
.A(n_2204),
.B(n_1838),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2061),
.Y(n_2444)
);

AND2x4_ASAP7_75t_L g2445 ( 
.A(n_2167),
.B(n_1909),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2058),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_2102),
.B(n_2018),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_2222),
.B(n_1847),
.Y(n_2448)
);

BUFx4_ASAP7_75t_L g2449 ( 
.A(n_2148),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2128),
.B(n_1847),
.Y(n_2450)
);

XNOR2x2_ASAP7_75t_L g2451 ( 
.A(n_2315),
.B(n_1846),
.Y(n_2451)
);

AND2x4_ASAP7_75t_L g2452 ( 
.A(n_2281),
.B(n_1909),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2109),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2061),
.Y(n_2454)
);

NOR2xp33_ASAP7_75t_L g2455 ( 
.A(n_2113),
.B(n_2122),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2069),
.Y(n_2456)
);

CKINVDCx5p33_ASAP7_75t_R g2457 ( 
.A(n_2087),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2115),
.Y(n_2458)
);

AOI22xp33_ASAP7_75t_SL g2459 ( 
.A1(n_2157),
.A2(n_1846),
.B1(n_2011),
.B2(n_2008),
.Y(n_2459)
);

OR2x2_ASAP7_75t_L g2460 ( 
.A(n_2174),
.B(n_1929),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2116),
.Y(n_2461)
);

AND2x4_ASAP7_75t_L g2462 ( 
.A(n_2281),
.B(n_1912),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_2110),
.B(n_2113),
.Y(n_2463)
);

AO22x2_ASAP7_75t_L g2464 ( 
.A1(n_2292),
.A2(n_2011),
.B1(n_2008),
.B2(n_1781),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2069),
.Y(n_2465)
);

NOR2xp33_ASAP7_75t_L g2466 ( 
.A(n_2122),
.B(n_1898),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2072),
.Y(n_2467)
);

AND2x4_ASAP7_75t_L g2468 ( 
.A(n_2287),
.B(n_1912),
.Y(n_2468)
);

AND2x6_ASAP7_75t_L g2469 ( 
.A(n_2300),
.B(n_2022),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_SL g2470 ( 
.A(n_2047),
.B(n_2050),
.Y(n_2470)
);

NOR2xp33_ASAP7_75t_L g2471 ( 
.A(n_2137),
.B(n_1898),
.Y(n_2471)
);

INVx4_ASAP7_75t_L g2472 ( 
.A(n_2056),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2137),
.B(n_1779),
.Y(n_2473)
);

BUFx2_ASAP7_75t_L g2474 ( 
.A(n_2057),
.Y(n_2474)
);

OR2x2_ASAP7_75t_L g2475 ( 
.A(n_2174),
.B(n_1936),
.Y(n_2475)
);

AND2x4_ASAP7_75t_L g2476 ( 
.A(n_2287),
.B(n_2147),
.Y(n_2476)
);

INVx2_ASAP7_75t_SL g2477 ( 
.A(n_2103),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2072),
.Y(n_2478)
);

INVxp33_ASAP7_75t_L g2479 ( 
.A(n_2199),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_SL g2480 ( 
.A(n_2047),
.B(n_1544),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2120),
.Y(n_2481)
);

AND2x4_ASAP7_75t_L g2482 ( 
.A(n_2147),
.B(n_1916),
.Y(n_2482)
);

AOI22xp33_ASAP7_75t_L g2483 ( 
.A1(n_2247),
.A2(n_1919),
.B1(n_1956),
.B2(n_1900),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2123),
.Y(n_2484)
);

INVx1_ASAP7_75t_SL g2485 ( 
.A(n_2160),
.Y(n_2485)
);

OAI221xp5_ASAP7_75t_L g2486 ( 
.A1(n_2253),
.A2(n_1961),
.B1(n_1955),
.B2(n_1950),
.C(n_1916),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2073),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2270),
.B(n_1921),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2073),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2076),
.Y(n_2490)
);

AOI22xp5_ASAP7_75t_L g2491 ( 
.A1(n_2234),
.A2(n_1681),
.B1(n_1781),
.B2(n_1974),
.Y(n_2491)
);

AND2x6_ASAP7_75t_L g2492 ( 
.A(n_2300),
.B(n_2022),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2076),
.Y(n_2493)
);

AND2x4_ASAP7_75t_L g2494 ( 
.A(n_2147),
.B(n_1917),
.Y(n_2494)
);

BUFx2_ASAP7_75t_L g2495 ( 
.A(n_2160),
.Y(n_2495)
);

BUFx6f_ASAP7_75t_L g2496 ( 
.A(n_2124),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2140),
.Y(n_2497)
);

AND2x4_ASAP7_75t_L g2498 ( 
.A(n_2186),
.B(n_1917),
.Y(n_2498)
);

AND2x4_ASAP7_75t_L g2499 ( 
.A(n_2186),
.B(n_1950),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2215),
.B(n_1955),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2140),
.Y(n_2501)
);

NAND2x1p5_ASAP7_75t_L g2502 ( 
.A(n_2166),
.B(n_1659),
.Y(n_2502)
);

INVx3_ASAP7_75t_L g2503 ( 
.A(n_2082),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2142),
.Y(n_2504)
);

AOI22xp5_ASAP7_75t_L g2505 ( 
.A1(n_2161),
.A2(n_1681),
.B1(n_1994),
.B2(n_1677),
.Y(n_2505)
);

INVx3_ASAP7_75t_L g2506 ( 
.A(n_2082),
.Y(n_2506)
);

AND2x4_ASAP7_75t_L g2507 ( 
.A(n_2188),
.B(n_1961),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2142),
.Y(n_2508)
);

AND2x4_ASAP7_75t_L g2509 ( 
.A(n_2188),
.B(n_1888),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2141),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2146),
.Y(n_2511)
);

NOR2xp33_ASAP7_75t_L g2512 ( 
.A(n_2183),
.B(n_1900),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2146),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2141),
.Y(n_2514)
);

INVx3_ASAP7_75t_L g2515 ( 
.A(n_2040),
.Y(n_2515)
);

BUFx2_ASAP7_75t_L g2516 ( 
.A(n_2291),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2247),
.B(n_2042),
.Y(n_2517)
);

CKINVDCx5p33_ASAP7_75t_R g2518 ( 
.A(n_2087),
.Y(n_2518)
);

INVx3_ASAP7_75t_L g2519 ( 
.A(n_2040),
.Y(n_2519)
);

AND2x4_ASAP7_75t_L g2520 ( 
.A(n_2291),
.B(n_1888),
.Y(n_2520)
);

HB1xp67_ASAP7_75t_L g2521 ( 
.A(n_2297),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2101),
.Y(n_2522)
);

HB1xp67_ASAP7_75t_L g2523 ( 
.A(n_2297),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2149),
.Y(n_2524)
);

CKINVDCx5p33_ASAP7_75t_R g2525 ( 
.A(n_2108),
.Y(n_2525)
);

NOR2xp33_ASAP7_75t_L g2526 ( 
.A(n_2187),
.B(n_1919),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_SL g2527 ( 
.A(n_2047),
.B(n_1551),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2118),
.B(n_1967),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_SL g2529 ( 
.A(n_2050),
.B(n_1551),
.Y(n_2529)
);

OR2x6_ASAP7_75t_L g2530 ( 
.A(n_2255),
.B(n_1581),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2131),
.Y(n_2531)
);

NAND3xp33_ASAP7_75t_L g2532 ( 
.A(n_2203),
.B(n_1967),
.C(n_1987),
.Y(n_2532)
);

AND2x4_ASAP7_75t_L g2533 ( 
.A(n_2202),
.B(n_1987),
.Y(n_2533)
);

NAND3xp33_ASAP7_75t_L g2534 ( 
.A(n_2203),
.B(n_1995),
.C(n_1914),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2131),
.Y(n_2535)
);

AND2x6_ASAP7_75t_L g2536 ( 
.A(n_2170),
.B(n_1995),
.Y(n_2536)
);

INVxp67_ASAP7_75t_SL g2537 ( 
.A(n_2177),
.Y(n_2537)
);

BUFx6f_ASAP7_75t_L g2538 ( 
.A(n_2124),
.Y(n_2538)
);

BUFx2_ASAP7_75t_L g2539 ( 
.A(n_2207),
.Y(n_2539)
);

INVx4_ASAP7_75t_L g2540 ( 
.A(n_2070),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2101),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2114),
.Y(n_2542)
);

AND2x4_ASAP7_75t_L g2543 ( 
.A(n_2202),
.B(n_1470),
.Y(n_2543)
);

OAI22xp5_ASAP7_75t_SL g2544 ( 
.A1(n_2257),
.A2(n_1956),
.B1(n_31),
.B2(n_29),
.Y(n_2544)
);

INVx5_ASAP7_75t_L g2545 ( 
.A(n_2106),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2114),
.Y(n_2546)
);

BUFx2_ASAP7_75t_L g2547 ( 
.A(n_2279),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_SL g2548 ( 
.A(n_2050),
.B(n_2086),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2131),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2145),
.B(n_1681),
.Y(n_2550)
);

AND2x2_ASAP7_75t_L g2551 ( 
.A(n_2118),
.B(n_1590),
.Y(n_2551)
);

INVxp67_ASAP7_75t_SL g2552 ( 
.A(n_2139),
.Y(n_2552)
);

BUFx3_ASAP7_75t_L g2553 ( 
.A(n_2070),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2355),
.B(n_2246),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2500),
.B(n_2326),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2355),
.B(n_2286),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2552),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_SL g2558 ( 
.A(n_2517),
.B(n_2162),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_2391),
.B(n_2119),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2368),
.Y(n_2560)
);

INVx2_ASAP7_75t_SL g2561 ( 
.A(n_2327),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2420),
.B(n_2286),
.Y(n_2562)
);

NOR2x1p5_ASAP7_75t_L g2563 ( 
.A(n_2460),
.B(n_2108),
.Y(n_2563)
);

AOI22xp5_ASAP7_75t_L g2564 ( 
.A1(n_2348),
.A2(n_2351),
.B1(n_2345),
.B2(n_2383),
.Y(n_2564)
);

AOI22xp33_ASAP7_75t_L g2565 ( 
.A1(n_2532),
.A2(n_2292),
.B1(n_2176),
.B2(n_2157),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2368),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2420),
.B(n_2118),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_SL g2568 ( 
.A(n_2372),
.B(n_2223),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2552),
.B(n_2132),
.Y(n_2569)
);

AOI22xp5_ASAP7_75t_L g2570 ( 
.A1(n_2348),
.A2(n_2081),
.B1(n_2195),
.B2(n_2261),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2339),
.B(n_2144),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2398),
.B(n_2173),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_SL g2573 ( 
.A(n_2372),
.B(n_2075),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_SL g2574 ( 
.A(n_2372),
.B(n_2304),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2353),
.B(n_2243),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2390),
.B(n_2243),
.Y(n_2576)
);

AOI22xp5_ASAP7_75t_L g2577 ( 
.A1(n_2351),
.A2(n_2081),
.B1(n_2099),
.B2(n_2220),
.Y(n_2577)
);

AND2x6_ASAP7_75t_L g2578 ( 
.A(n_2415),
.B(n_2277),
.Y(n_2578)
);

HB1xp67_ASAP7_75t_L g2579 ( 
.A(n_2485),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2423),
.B(n_2175),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2390),
.B(n_2243),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2400),
.B(n_2249),
.Y(n_2582)
);

AND2x4_ASAP7_75t_L g2583 ( 
.A(n_2424),
.B(n_2202),
.Y(n_2583)
);

NOR2xp33_ASAP7_75t_L g2584 ( 
.A(n_2479),
.B(n_2292),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2400),
.B(n_2249),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2352),
.B(n_2310),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_SL g2587 ( 
.A(n_2450),
.B(n_2189),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2429),
.B(n_2537),
.Y(n_2588)
);

BUFx3_ASAP7_75t_L g2589 ( 
.A(n_2327),
.Y(n_2589)
);

INVx3_ASAP7_75t_L g2590 ( 
.A(n_2515),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2343),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_SL g2592 ( 
.A(n_2448),
.B(n_2205),
.Y(n_2592)
);

CKINVDCx20_ASAP7_75t_R g2593 ( 
.A(n_2361),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_L g2594 ( 
.A(n_2479),
.B(n_2044),
.Y(n_2594)
);

INVx2_ASAP7_75t_SL g2595 ( 
.A(n_2402),
.Y(n_2595)
);

AOI22xp5_ASAP7_75t_L g2596 ( 
.A1(n_2345),
.A2(n_2099),
.B1(n_2051),
.B2(n_2257),
.Y(n_2596)
);

AOI22xp33_ASAP7_75t_L g2597 ( 
.A1(n_2328),
.A2(n_2176),
.B1(n_2157),
.B2(n_2091),
.Y(n_2597)
);

NAND2x1_ASAP7_75t_L g2598 ( 
.A(n_2515),
.B(n_2086),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2429),
.B(n_2250),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2537),
.B(n_2250),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2344),
.Y(n_2601)
);

NAND2xp33_ASAP7_75t_L g2602 ( 
.A(n_2378),
.B(n_2157),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2395),
.Y(n_2603)
);

HB1xp67_ASAP7_75t_L g2604 ( 
.A(n_2495),
.Y(n_2604)
);

AOI22xp5_ASAP7_75t_SL g2605 ( 
.A1(n_2427),
.A2(n_2079),
.B1(n_2143),
.B2(n_2157),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2443),
.B(n_2178),
.Y(n_2606)
);

AOI22xp5_ASAP7_75t_L g2607 ( 
.A1(n_2404),
.A2(n_2293),
.B1(n_2214),
.B2(n_2308),
.Y(n_2607)
);

NOR2xp33_ASAP7_75t_L g2608 ( 
.A(n_2333),
.B(n_2044),
.Y(n_2608)
);

O2A1O1Ixp33_ASAP7_75t_L g2609 ( 
.A1(n_2325),
.A2(n_2268),
.B(n_2285),
.C(n_2275),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2448),
.B(n_2254),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_SL g2611 ( 
.A(n_2325),
.B(n_2208),
.Y(n_2611)
);

NOR2xp33_ASAP7_75t_L g2612 ( 
.A(n_2333),
.B(n_2044),
.Y(n_2612)
);

AOI22xp33_ASAP7_75t_L g2613 ( 
.A1(n_2328),
.A2(n_2176),
.B1(n_2091),
.B2(n_2272),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2442),
.B(n_2254),
.Y(n_2614)
);

NOR2xp33_ASAP7_75t_L g2615 ( 
.A(n_2371),
.B(n_2306),
.Y(n_2615)
);

AND2x2_ASAP7_75t_SL g2616 ( 
.A(n_2433),
.B(n_2226),
.Y(n_2616)
);

AOI22xp5_ASAP7_75t_L g2617 ( 
.A1(n_2404),
.A2(n_2350),
.B1(n_2377),
.B2(n_2338),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2399),
.Y(n_2618)
);

INVx3_ASAP7_75t_L g2619 ( 
.A(n_2519),
.Y(n_2619)
);

NAND2xp33_ASAP7_75t_L g2620 ( 
.A(n_2378),
.B(n_2176),
.Y(n_2620)
);

AOI22xp33_ASAP7_75t_L g2621 ( 
.A1(n_2534),
.A2(n_2176),
.B1(n_2091),
.B2(n_2170),
.Y(n_2621)
);

NAND3xp33_ASAP7_75t_SL g2622 ( 
.A(n_2367),
.B(n_2079),
.C(n_2129),
.Y(n_2622)
);

AOI21xp5_ASAP7_75t_L g2623 ( 
.A1(n_2550),
.A2(n_2059),
.B(n_2212),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2359),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2442),
.B(n_2259),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2363),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2551),
.B(n_2259),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2366),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2399),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2488),
.B(n_2260),
.Y(n_2630)
);

O2A1O1Ixp33_ASAP7_75t_L g2631 ( 
.A1(n_2338),
.A2(n_2447),
.B(n_2377),
.C(n_2347),
.Y(n_2631)
);

AOI22xp5_ASAP7_75t_L g2632 ( 
.A1(n_2430),
.A2(n_2053),
.B1(n_2176),
.B2(n_2153),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2463),
.B(n_2260),
.Y(n_2633)
);

O2A1O1Ixp5_ASAP7_75t_L g2634 ( 
.A1(n_2447),
.A2(n_2094),
.B(n_2228),
.C(n_2218),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2382),
.B(n_2265),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2475),
.B(n_2179),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2371),
.B(n_2520),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2499),
.B(n_2265),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2499),
.B(n_2273),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2507),
.B(n_2452),
.Y(n_2640)
);

AND2x6_ASAP7_75t_SL g2641 ( 
.A(n_2340),
.B(n_2053),
.Y(n_2641)
);

INVx3_ASAP7_75t_L g2642 ( 
.A(n_2496),
.Y(n_2642)
);

AND2x2_ASAP7_75t_SL g2643 ( 
.A(n_2433),
.B(n_2226),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2507),
.B(n_2273),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2452),
.B(n_2227),
.Y(n_2645)
);

AOI22xp33_ASAP7_75t_L g2646 ( 
.A1(n_2451),
.A2(n_2091),
.B1(n_2268),
.B2(n_2277),
.Y(n_2646)
);

AOI22xp5_ASAP7_75t_L g2647 ( 
.A1(n_2413),
.A2(n_2053),
.B1(n_2153),
.B2(n_2151),
.Y(n_2647)
);

INVx2_ASAP7_75t_SL g2648 ( 
.A(n_2402),
.Y(n_2648)
);

AOI22xp33_ASAP7_75t_L g2649 ( 
.A1(n_2544),
.A2(n_2268),
.B1(n_2280),
.B2(n_2245),
.Y(n_2649)
);

NAND3xp33_ASAP7_75t_SL g2650 ( 
.A(n_2396),
.B(n_2274),
.C(n_2262),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_SL g2651 ( 
.A(n_2412),
.B(n_2217),
.Y(n_2651)
);

INVxp67_ASAP7_75t_L g2652 ( 
.A(n_2539),
.Y(n_2652)
);

AND2x2_ASAP7_75t_L g2653 ( 
.A(n_2520),
.B(n_2181),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2373),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2375),
.Y(n_2655)
);

NOR2xp33_ASAP7_75t_L g2656 ( 
.A(n_2341),
.B(n_2306),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2376),
.Y(n_2657)
);

INVx4_ASAP7_75t_L g2658 ( 
.A(n_2378),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2462),
.B(n_2468),
.Y(n_2659)
);

OR2x6_ASAP7_75t_L g2660 ( 
.A(n_2360),
.B(n_2255),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2381),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2462),
.B(n_2227),
.Y(n_2662)
);

OR2x2_ASAP7_75t_L g2663 ( 
.A(n_2408),
.B(n_2191),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2528),
.B(n_2196),
.Y(n_2664)
);

CKINVDCx5p33_ASAP7_75t_R g2665 ( 
.A(n_2457),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2468),
.B(n_2227),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2384),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_SL g2668 ( 
.A(n_2418),
.B(n_2062),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2466),
.B(n_2168),
.Y(n_2669)
);

AOI22xp5_ASAP7_75t_L g2670 ( 
.A1(n_2413),
.A2(n_2053),
.B1(n_2153),
.B2(n_2151),
.Y(n_2670)
);

AOI22xp33_ASAP7_75t_L g2671 ( 
.A1(n_2459),
.A2(n_2536),
.B1(n_2401),
.B2(n_2526),
.Y(n_2671)
);

AND2x6_ASAP7_75t_L g2672 ( 
.A(n_2415),
.B(n_2280),
.Y(n_2672)
);

NOR2xp33_ASAP7_75t_L g2673 ( 
.A(n_2403),
.B(n_2306),
.Y(n_2673)
);

INVx3_ASAP7_75t_L g2674 ( 
.A(n_2496),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2466),
.B(n_2168),
.Y(n_2675)
);

AND2x2_ASAP7_75t_SL g2676 ( 
.A(n_2512),
.B(n_2226),
.Y(n_2676)
);

NOR2xp33_ASAP7_75t_L g2677 ( 
.A(n_2329),
.B(n_2172),
.Y(n_2677)
);

AO22x1_ASAP7_75t_L g2678 ( 
.A1(n_2396),
.A2(n_2290),
.B1(n_2282),
.B2(n_2299),
.Y(n_2678)
);

BUFx3_ASAP7_75t_L g2679 ( 
.A(n_2387),
.Y(n_2679)
);

NOR2xp33_ASAP7_75t_L g2680 ( 
.A(n_2521),
.B(n_2523),
.Y(n_2680)
);

BUFx6f_ASAP7_75t_L g2681 ( 
.A(n_2331),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2385),
.Y(n_2682)
);

AOI22xp5_ASAP7_75t_L g2683 ( 
.A1(n_2482),
.A2(n_2151),
.B1(n_2244),
.B2(n_2190),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2471),
.B(n_2455),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2407),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_SL g2686 ( 
.A(n_2512),
.B(n_2314),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2417),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2417),
.Y(n_2688)
);

BUFx3_ASAP7_75t_L g2689 ( 
.A(n_2553),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2431),
.Y(n_2690)
);

BUFx3_ASAP7_75t_L g2691 ( 
.A(n_2553),
.Y(n_2691)
);

OR2x6_ASAP7_75t_L g2692 ( 
.A(n_2516),
.B(n_2238),
.Y(n_2692)
);

INVx3_ASAP7_75t_L g2693 ( 
.A(n_2496),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_SL g2694 ( 
.A(n_2526),
.B(n_2094),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2471),
.B(n_2172),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_SL g2696 ( 
.A(n_2422),
.B(n_2242),
.Y(n_2696)
);

AOI22xp33_ASAP7_75t_L g2697 ( 
.A1(n_2459),
.A2(n_2240),
.B1(n_2245),
.B2(n_2258),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2455),
.B(n_2172),
.Y(n_2698)
);

NOR2xp33_ASAP7_75t_L g2699 ( 
.A(n_2521),
.B(n_2169),
.Y(n_2699)
);

BUFx6f_ASAP7_75t_SL g2700 ( 
.A(n_2424),
.Y(n_2700)
);

NOR2xp33_ASAP7_75t_L g2701 ( 
.A(n_2523),
.B(n_2185),
.Y(n_2701)
);

OR2x2_ASAP7_75t_L g2702 ( 
.A(n_2477),
.B(n_2198),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2509),
.B(n_2258),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2431),
.Y(n_2704)
);

AND2x6_ASAP7_75t_SL g2705 ( 
.A(n_2340),
.B(n_2077),
.Y(n_2705)
);

OAI22xp5_ASAP7_75t_L g2706 ( 
.A1(n_2482),
.A2(n_2238),
.B1(n_2206),
.B2(n_2316),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2509),
.B(n_2264),
.Y(n_2707)
);

NOR2xp33_ASAP7_75t_L g2708 ( 
.A(n_2486),
.B(n_2185),
.Y(n_2708)
);

INVx4_ASAP7_75t_L g2709 ( 
.A(n_2545),
.Y(n_2709)
);

OAI21xp5_ASAP7_75t_L g2710 ( 
.A1(n_2401),
.A2(n_2321),
.B(n_2252),
.Y(n_2710)
);

AOI21xp5_ASAP7_75t_L g2711 ( 
.A1(n_2480),
.A2(n_2059),
.B(n_2088),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2498),
.B(n_2264),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2498),
.B(n_2266),
.Y(n_2713)
);

AND2x2_ASAP7_75t_L g2714 ( 
.A(n_2389),
.B(n_2200),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2428),
.B(n_2266),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2388),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2432),
.Y(n_2717)
);

OAI22xp5_ASAP7_75t_L g2718 ( 
.A1(n_2494),
.A2(n_2238),
.B1(n_2316),
.B2(n_2213),
.Y(n_2718)
);

NAND2xp33_ASAP7_75t_L g2719 ( 
.A(n_2496),
.B(n_2282),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2434),
.B(n_2299),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2432),
.Y(n_2721)
);

AOI22xp33_ASAP7_75t_L g2722 ( 
.A1(n_2536),
.A2(n_2240),
.B1(n_2311),
.B2(n_2269),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_2536),
.B(n_2269),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2393),
.Y(n_2724)
);

AOI22xp5_ASAP7_75t_L g2725 ( 
.A1(n_2494),
.A2(n_2163),
.B1(n_2190),
.B2(n_2238),
.Y(n_2725)
);

NOR2xp33_ASAP7_75t_L g2726 ( 
.A(n_2356),
.B(n_2185),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2394),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2435),
.B(n_2299),
.Y(n_2728)
);

AOI22xp5_ASAP7_75t_L g2729 ( 
.A1(n_2332),
.A2(n_2163),
.B1(n_2190),
.B2(n_2124),
.Y(n_2729)
);

OAI22x1_ASAP7_75t_R g2730 ( 
.A1(n_2427),
.A2(n_2171),
.B1(n_2090),
.B2(n_2163),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2474),
.B(n_2283),
.Y(n_2731)
);

INVxp67_ASAP7_75t_L g2732 ( 
.A(n_2547),
.Y(n_2732)
);

OAI22xp5_ASAP7_75t_SL g2733 ( 
.A1(n_2340),
.A2(n_2283),
.B1(n_2282),
.B2(n_2290),
.Y(n_2733)
);

A2O1A1Ixp33_ASAP7_75t_L g2734 ( 
.A1(n_2406),
.A2(n_2295),
.B(n_2312),
.C(n_2311),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2536),
.B(n_2312),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2536),
.B(n_2323),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2684),
.B(n_2483),
.Y(n_2737)
);

AOI22xp5_ASAP7_75t_L g2738 ( 
.A1(n_2564),
.A2(n_2392),
.B1(n_2533),
.B2(n_2346),
.Y(n_2738)
);

NOR2x1p5_ASAP7_75t_L g2739 ( 
.A(n_2622),
.B(n_2518),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2591),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2715),
.B(n_2483),
.Y(n_2741)
);

INVxp67_ASAP7_75t_L g2742 ( 
.A(n_2579),
.Y(n_2742)
);

INVx3_ASAP7_75t_L g2743 ( 
.A(n_2658),
.Y(n_2743)
);

CKINVDCx11_ASAP7_75t_R g2744 ( 
.A(n_2593),
.Y(n_2744)
);

AOI22xp5_ASAP7_75t_L g2745 ( 
.A1(n_2577),
.A2(n_2392),
.B1(n_2533),
.B2(n_2346),
.Y(n_2745)
);

AND2x6_ASAP7_75t_L g2746 ( 
.A(n_2632),
.B(n_2230),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2555),
.B(n_2473),
.Y(n_2747)
);

INVx2_ASAP7_75t_SL g2748 ( 
.A(n_2689),
.Y(n_2748)
);

INVx3_ASAP7_75t_L g2749 ( 
.A(n_2658),
.Y(n_2749)
);

AND2x6_ASAP7_75t_L g2750 ( 
.A(n_2647),
.B(n_2230),
.Y(n_2750)
);

AND2x2_ASAP7_75t_L g2751 ( 
.A(n_2637),
.B(n_2392),
.Y(n_2751)
);

AND2x4_ASAP7_75t_L g2752 ( 
.A(n_2583),
.B(n_2438),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2560),
.Y(n_2753)
);

OAI22xp5_ASAP7_75t_L g2754 ( 
.A1(n_2649),
.A2(n_2357),
.B1(n_2425),
.B2(n_2323),
.Y(n_2754)
);

INVx3_ASAP7_75t_L g2755 ( 
.A(n_2709),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2566),
.Y(n_2756)
);

INVx3_ASAP7_75t_L g2757 ( 
.A(n_2709),
.Y(n_2757)
);

BUFx3_ASAP7_75t_L g2758 ( 
.A(n_2691),
.Y(n_2758)
);

AND2x2_ASAP7_75t_L g2759 ( 
.A(n_2664),
.B(n_2440),
.Y(n_2759)
);

OAI22xp33_ASAP7_75t_L g2760 ( 
.A1(n_2617),
.A2(n_2491),
.B1(n_2414),
.B2(n_2439),
.Y(n_2760)
);

BUFx3_ASAP7_75t_L g2761 ( 
.A(n_2589),
.Y(n_2761)
);

BUFx2_ASAP7_75t_L g2762 ( 
.A(n_2679),
.Y(n_2762)
);

AO22x1_ASAP7_75t_L g2763 ( 
.A1(n_2594),
.A2(n_2290),
.B1(n_2525),
.B2(n_2476),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_2583),
.B(n_2438),
.Y(n_2764)
);

OAI21xp5_ASAP7_75t_L g2765 ( 
.A1(n_2710),
.A2(n_2278),
.B(n_2271),
.Y(n_2765)
);

INVx2_ASAP7_75t_SL g2766 ( 
.A(n_2561),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2631),
.B(n_2337),
.Y(n_2767)
);

NOR2xp33_ASAP7_75t_L g2768 ( 
.A(n_2567),
.B(n_2332),
.Y(n_2768)
);

HB1xp67_ASAP7_75t_L g2769 ( 
.A(n_2588),
.Y(n_2769)
);

INVxp67_ASAP7_75t_SL g2770 ( 
.A(n_2557),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2559),
.B(n_2342),
.Y(n_2771)
);

AND2x4_ASAP7_75t_L g2772 ( 
.A(n_2692),
.B(n_2440),
.Y(n_2772)
);

BUFx6f_ASAP7_75t_L g2773 ( 
.A(n_2681),
.Y(n_2773)
);

OAI22xp5_ASAP7_75t_L g2774 ( 
.A1(n_2649),
.A2(n_2357),
.B1(n_2464),
.B2(n_2288),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2559),
.B(n_2441),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2601),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2603),
.Y(n_2777)
);

BUFx6f_ASAP7_75t_L g2778 ( 
.A(n_2681),
.Y(n_2778)
);

BUFx2_ASAP7_75t_L g2779 ( 
.A(n_2579),
.Y(n_2779)
);

AOI22xp33_ASAP7_75t_L g2780 ( 
.A1(n_2650),
.A2(n_2357),
.B1(n_2464),
.B2(n_2441),
.Y(n_2780)
);

AOI22xp5_ASAP7_75t_L g2781 ( 
.A1(n_2570),
.A2(n_2380),
.B1(n_2397),
.B2(n_2374),
.Y(n_2781)
);

OR2x2_ASAP7_75t_L g2782 ( 
.A(n_2562),
.B(n_2437),
.Y(n_2782)
);

AND2x4_ASAP7_75t_L g2783 ( 
.A(n_2692),
.B(n_2476),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2624),
.Y(n_2784)
);

BUFx2_ASAP7_75t_L g2785 ( 
.A(n_2604),
.Y(n_2785)
);

BUFx3_ASAP7_75t_L g2786 ( 
.A(n_2595),
.Y(n_2786)
);

INVx6_ASAP7_75t_L g2787 ( 
.A(n_2692),
.Y(n_2787)
);

INVxp67_ASAP7_75t_L g2788 ( 
.A(n_2680),
.Y(n_2788)
);

INVxp67_ASAP7_75t_L g2789 ( 
.A(n_2680),
.Y(n_2789)
);

BUFx3_ASAP7_75t_L g2790 ( 
.A(n_2648),
.Y(n_2790)
);

BUFx2_ASAP7_75t_L g2791 ( 
.A(n_2604),
.Y(n_2791)
);

HB1xp67_ASAP7_75t_L g2792 ( 
.A(n_2723),
.Y(n_2792)
);

AND2x4_ASAP7_75t_SL g2793 ( 
.A(n_2731),
.B(n_2386),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2610),
.B(n_2441),
.Y(n_2794)
);

AOI22xp33_ASAP7_75t_L g2795 ( 
.A1(n_2671),
.A2(n_2464),
.B1(n_2469),
.B2(n_2441),
.Y(n_2795)
);

AOI22xp5_ASAP7_75t_L g2796 ( 
.A1(n_2708),
.A2(n_2380),
.B1(n_2397),
.B2(n_2374),
.Y(n_2796)
);

AOI22xp5_ASAP7_75t_L g2797 ( 
.A1(n_2708),
.A2(n_2445),
.B1(n_2283),
.B2(n_2282),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2554),
.B(n_2441),
.Y(n_2798)
);

BUFx6f_ASAP7_75t_L g2799 ( 
.A(n_2681),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2626),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_SL g2801 ( 
.A(n_2607),
.B(n_2290),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2618),
.Y(n_2802)
);

NOR2xp33_ASAP7_75t_L g2803 ( 
.A(n_2659),
.B(n_2445),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2628),
.Y(n_2804)
);

NOR2xp33_ASAP7_75t_L g2805 ( 
.A(n_2640),
.B(n_2282),
.Y(n_2805)
);

AOI22xp33_ASAP7_75t_L g2806 ( 
.A1(n_2671),
.A2(n_2492),
.B1(n_2469),
.B2(n_2446),
.Y(n_2806)
);

NOR2xp33_ASAP7_75t_L g2807 ( 
.A(n_2584),
.B(n_2453),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2629),
.Y(n_2808)
);

INVx4_ASAP7_75t_L g2809 ( 
.A(n_2700),
.Y(n_2809)
);

O2A1O1Ixp33_ASAP7_75t_L g2810 ( 
.A1(n_2694),
.A2(n_2248),
.B(n_2461),
.C(n_2458),
.Y(n_2810)
);

NAND2x1p5_ASAP7_75t_L g2811 ( 
.A(n_2574),
.B(n_2545),
.Y(n_2811)
);

BUFx4f_ASAP7_75t_L g2812 ( 
.A(n_2660),
.Y(n_2812)
);

BUFx2_ASAP7_75t_L g2813 ( 
.A(n_2652),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2654),
.Y(n_2814)
);

INVxp67_ASAP7_75t_SL g2815 ( 
.A(n_2600),
.Y(n_2815)
);

OR2x6_ASAP7_75t_L g2816 ( 
.A(n_2733),
.B(n_2065),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_SL g2817 ( 
.A(n_2676),
.B(n_2233),
.Y(n_2817)
);

AND2x4_ASAP7_75t_L g2818 ( 
.A(n_2660),
.B(n_2386),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2655),
.Y(n_2819)
);

BUFx6f_ASAP7_75t_L g2820 ( 
.A(n_2660),
.Y(n_2820)
);

INVx3_ASAP7_75t_L g2821 ( 
.A(n_2590),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2657),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_SL g2823 ( 
.A(n_2596),
.B(n_2305),
.Y(n_2823)
);

BUFx8_ASAP7_75t_L g2824 ( 
.A(n_2700),
.Y(n_2824)
);

BUFx3_ASAP7_75t_L g2825 ( 
.A(n_2665),
.Y(n_2825)
);

INVx2_ASAP7_75t_SL g2826 ( 
.A(n_2563),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2685),
.Y(n_2827)
);

INVx3_ASAP7_75t_L g2828 ( 
.A(n_2590),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2687),
.Y(n_2829)
);

BUFx2_ASAP7_75t_L g2830 ( 
.A(n_2652),
.Y(n_2830)
);

OR2x6_ASAP7_75t_L g2831 ( 
.A(n_2678),
.B(n_2065),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2661),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2734),
.B(n_2469),
.Y(n_2833)
);

BUFx6f_ASAP7_75t_L g2834 ( 
.A(n_2720),
.Y(n_2834)
);

NAND2x1p5_ASAP7_75t_L g2835 ( 
.A(n_2574),
.B(n_2545),
.Y(n_2835)
);

OR2x6_ASAP7_75t_L g2836 ( 
.A(n_2573),
.B(n_2065),
.Y(n_2836)
);

OR2x6_ASAP7_75t_L g2837 ( 
.A(n_2573),
.B(n_2065),
.Y(n_2837)
);

INVx4_ASAP7_75t_L g2838 ( 
.A(n_2642),
.Y(n_2838)
);

NOR2xp33_ASAP7_75t_L g2839 ( 
.A(n_2584),
.B(n_2481),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2667),
.Y(n_2840)
);

INVx4_ASAP7_75t_L g2841 ( 
.A(n_2642),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2682),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2636),
.B(n_2484),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2688),
.Y(n_2844)
);

INVx4_ASAP7_75t_L g2845 ( 
.A(n_2674),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2716),
.Y(n_2846)
);

INVx3_ASAP7_75t_L g2847 ( 
.A(n_2619),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2734),
.B(n_2469),
.Y(n_2848)
);

HB1xp67_ASAP7_75t_L g2849 ( 
.A(n_2735),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2724),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2673),
.B(n_2492),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2722),
.B(n_2492),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2727),
.Y(n_2853)
);

CKINVDCx5p33_ASAP7_75t_R g2854 ( 
.A(n_2705),
.Y(n_2854)
);

BUFx3_ASAP7_75t_L g2855 ( 
.A(n_2728),
.Y(n_2855)
);

NOR2xp33_ASAP7_75t_L g2856 ( 
.A(n_2571),
.B(n_2124),
.Y(n_2856)
);

O2A1O1Ixp33_ASAP7_75t_L g2857 ( 
.A1(n_2694),
.A2(n_2248),
.B(n_2236),
.C(n_2235),
.Y(n_2857)
);

NOR2xp33_ASAP7_75t_L g2858 ( 
.A(n_2556),
.B(n_2124),
.Y(n_2858)
);

CKINVDCx20_ASAP7_75t_R g2859 ( 
.A(n_2730),
.Y(n_2859)
);

INVxp67_ASAP7_75t_L g2860 ( 
.A(n_2615),
.Y(n_2860)
);

CKINVDCx5p33_ASAP7_75t_R g2861 ( 
.A(n_2594),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2690),
.Y(n_2862)
);

AOI22xp33_ASAP7_75t_L g2863 ( 
.A1(n_2686),
.A2(n_2492),
.B1(n_2334),
.B2(n_2411),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2576),
.Y(n_2864)
);

AND2x4_ASAP7_75t_L g2865 ( 
.A(n_2653),
.B(n_2472),
.Y(n_2865)
);

INVxp67_ASAP7_75t_L g2866 ( 
.A(n_2615),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_SL g2867 ( 
.A(n_2608),
.B(n_2233),
.Y(n_2867)
);

AND2x4_ASAP7_75t_L g2868 ( 
.A(n_2572),
.B(n_2472),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2581),
.Y(n_2869)
);

BUFx6f_ASAP7_75t_L g2870 ( 
.A(n_2714),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2704),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2717),
.Y(n_2872)
);

INVx2_ASAP7_75t_SL g2873 ( 
.A(n_2702),
.Y(n_2873)
);

BUFx6f_ASAP7_75t_L g2874 ( 
.A(n_2674),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2721),
.Y(n_2875)
);

BUFx6f_ASAP7_75t_L g2876 ( 
.A(n_2693),
.Y(n_2876)
);

INVxp67_ASAP7_75t_L g2877 ( 
.A(n_2663),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_2614),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2625),
.Y(n_2879)
);

HB1xp67_ASAP7_75t_L g2880 ( 
.A(n_2736),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2582),
.Y(n_2881)
);

INVx2_ASAP7_75t_SL g2882 ( 
.A(n_2580),
.Y(n_2882)
);

INVx3_ASAP7_75t_L g2883 ( 
.A(n_2619),
.Y(n_2883)
);

AND2x4_ASAP7_75t_SL g2884 ( 
.A(n_2606),
.B(n_2540),
.Y(n_2884)
);

HB1xp67_ASAP7_75t_L g2885 ( 
.A(n_2585),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2722),
.B(n_2492),
.Y(n_2886)
);

HB1xp67_ASAP7_75t_L g2887 ( 
.A(n_2599),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2635),
.Y(n_2888)
);

INVx2_ASAP7_75t_SL g2889 ( 
.A(n_2693),
.Y(n_2889)
);

INVxp67_ASAP7_75t_L g2890 ( 
.A(n_2699),
.Y(n_2890)
);

BUFx2_ASAP7_75t_L g2891 ( 
.A(n_2732),
.Y(n_2891)
);

AOI21xp5_ASAP7_75t_L g2892 ( 
.A1(n_2602),
.A2(n_2209),
.B(n_2294),
.Y(n_2892)
);

BUFx2_ASAP7_75t_L g2893 ( 
.A(n_2732),
.Y(n_2893)
);

CKINVDCx5p33_ASAP7_75t_R g2894 ( 
.A(n_2608),
.Y(n_2894)
);

AOI211xp5_ASAP7_75t_L g2895 ( 
.A1(n_2656),
.A2(n_2251),
.B(n_1937),
.C(n_1942),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2638),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2639),
.Y(n_2897)
);

HB1xp67_ASAP7_75t_L g2898 ( 
.A(n_2569),
.Y(n_2898)
);

INVx6_ASAP7_75t_L g2899 ( 
.A(n_2641),
.Y(n_2899)
);

AND3x1_ASAP7_75t_SL g2900 ( 
.A(n_2605),
.B(n_2497),
.C(n_2410),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2644),
.Y(n_2901)
);

OR2x6_ASAP7_75t_L g2902 ( 
.A(n_2718),
.B(n_2530),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2697),
.B(n_2501),
.Y(n_2903)
);

AND2x6_ASAP7_75t_L g2904 ( 
.A(n_2670),
.B(n_2415),
.Y(n_2904)
);

NAND3xp33_ASAP7_75t_L g2905 ( 
.A(n_2565),
.B(n_2125),
.C(n_2317),
.Y(n_2905)
);

INVx3_ASAP7_75t_L g2906 ( 
.A(n_2578),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2627),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2656),
.B(n_2510),
.Y(n_2908)
);

INVx3_ASAP7_75t_L g2909 ( 
.A(n_2578),
.Y(n_2909)
);

INVx3_ASAP7_75t_L g2910 ( 
.A(n_2578),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2712),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2770),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2770),
.Y(n_2913)
);

AND2x4_ASAP7_75t_L g2914 ( 
.A(n_2855),
.B(n_2729),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2769),
.Y(n_2915)
);

AOI21xp5_ASAP7_75t_L g2916 ( 
.A1(n_2801),
.A2(n_2620),
.B(n_2719),
.Y(n_2916)
);

AOI21xp5_ASAP7_75t_L g2917 ( 
.A1(n_2801),
.A2(n_2565),
.B(n_2686),
.Y(n_2917)
);

AOI21xp5_ASAP7_75t_L g2918 ( 
.A1(n_2767),
.A2(n_2558),
.B(n_2592),
.Y(n_2918)
);

AOI33xp33_ASAP7_75t_L g2919 ( 
.A1(n_2780),
.A2(n_2621),
.A3(n_2613),
.B1(n_2697),
.B2(n_2597),
.B3(n_2646),
.Y(n_2919)
);

AOI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2892),
.A2(n_2823),
.B(n_2857),
.Y(n_2920)
);

NOR2xp33_ASAP7_75t_SL g2921 ( 
.A(n_2809),
.B(n_2540),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2769),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2753),
.Y(n_2923)
);

OAI22xp5_ASAP7_75t_L g2924 ( 
.A1(n_2806),
.A2(n_2597),
.B1(n_2613),
.B2(n_2616),
.Y(n_2924)
);

A2O1A1Ixp33_ASAP7_75t_L g2925 ( 
.A1(n_2738),
.A2(n_2634),
.B(n_2643),
.C(n_2616),
.Y(n_2925)
);

AOI21x1_ASAP7_75t_L g2926 ( 
.A1(n_2763),
.A2(n_2611),
.B(n_2651),
.Y(n_2926)
);

OAI21xp5_ASAP7_75t_L g2927 ( 
.A1(n_2857),
.A2(n_2611),
.B(n_2586),
.Y(n_2927)
);

AOI21xp5_ASAP7_75t_L g2928 ( 
.A1(n_2892),
.A2(n_2568),
.B(n_2651),
.Y(n_2928)
);

INVx1_ASAP7_75t_SL g2929 ( 
.A(n_2779),
.Y(n_2929)
);

OAI22x1_ASAP7_75t_L g2930 ( 
.A1(n_2745),
.A2(n_2683),
.B1(n_2612),
.B2(n_2725),
.Y(n_2930)
);

A2O1A1Ixp33_ASAP7_75t_L g2931 ( 
.A1(n_2806),
.A2(n_2643),
.B(n_2609),
.C(n_2677),
.Y(n_2931)
);

AOI21xp5_ASAP7_75t_L g2932 ( 
.A1(n_2823),
.A2(n_2568),
.B(n_2587),
.Y(n_2932)
);

OAI22xp5_ASAP7_75t_L g2933 ( 
.A1(n_2795),
.A2(n_2621),
.B1(n_2646),
.B2(n_2703),
.Y(n_2933)
);

HB1xp67_ASAP7_75t_L g2934 ( 
.A(n_2785),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2911),
.B(n_2707),
.Y(n_2935)
);

AND2x2_ASAP7_75t_L g2936 ( 
.A(n_2747),
.B(n_2677),
.Y(n_2936)
);

AND2x2_ASAP7_75t_L g2937 ( 
.A(n_2751),
.B(n_2759),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2756),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2901),
.B(n_2713),
.Y(n_2939)
);

AOI21xp5_ASAP7_75t_L g2940 ( 
.A1(n_2815),
.A2(n_2587),
.B(n_2586),
.Y(n_2940)
);

AOI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2815),
.A2(n_2706),
.B(n_2711),
.Y(n_2941)
);

AOI22xp33_ASAP7_75t_SL g2942 ( 
.A1(n_2750),
.A2(n_2672),
.B1(n_2334),
.B2(n_2669),
.Y(n_2942)
);

OA22x2_ASAP7_75t_L g2943 ( 
.A1(n_2754),
.A2(n_2630),
.B1(n_2575),
.B2(n_2675),
.Y(n_2943)
);

AOI21xp5_ASAP7_75t_L g2944 ( 
.A1(n_2831),
.A2(n_2696),
.B(n_2623),
.Y(n_2944)
);

O2A1O1Ixp33_ASAP7_75t_L g2945 ( 
.A1(n_2760),
.A2(n_2668),
.B(n_2696),
.C(n_2695),
.Y(n_2945)
);

BUFx2_ASAP7_75t_L g2946 ( 
.A(n_2772),
.Y(n_2946)
);

NOR2xp33_ASAP7_75t_L g2947 ( 
.A(n_2861),
.B(n_2894),
.Y(n_2947)
);

O2A1O1Ixp33_ASAP7_75t_L g2948 ( 
.A1(n_2760),
.A2(n_2668),
.B(n_2662),
.C(n_2666),
.Y(n_2948)
);

NAND3xp33_ASAP7_75t_L g2949 ( 
.A(n_2895),
.B(n_2645),
.C(n_2701),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2898),
.B(n_2633),
.Y(n_2950)
);

NOR2x1_ASAP7_75t_R g2951 ( 
.A(n_2744),
.B(n_2449),
.Y(n_2951)
);

NOR2xp67_ASAP7_75t_L g2952 ( 
.A(n_2826),
.B(n_2726),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_L g2953 ( 
.A(n_2896),
.B(n_2698),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2834),
.B(n_2699),
.Y(n_2954)
);

AOI21xp5_ASAP7_75t_L g2955 ( 
.A1(n_2810),
.A2(n_2041),
.B(n_2302),
.Y(n_2955)
);

AOI21xp5_ASAP7_75t_L g2956 ( 
.A1(n_2810),
.A2(n_2527),
.B(n_2480),
.Y(n_2956)
);

NOR2xp33_ASAP7_75t_L g2957 ( 
.A(n_2834),
.B(n_2233),
.Y(n_2957)
);

AOI22xp5_ASAP7_75t_L g2958 ( 
.A1(n_2739),
.A2(n_2305),
.B1(n_2672),
.B2(n_2241),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_SL g2959 ( 
.A(n_2768),
.B(n_2514),
.Y(n_2959)
);

NOR2xp33_ASAP7_75t_SL g2960 ( 
.A(n_2809),
.B(n_2104),
.Y(n_2960)
);

AOI21xp5_ASAP7_75t_L g2961 ( 
.A1(n_2765),
.A2(n_2529),
.B(n_2527),
.Y(n_2961)
);

AOI21xp5_ASAP7_75t_L g2962 ( 
.A1(n_2771),
.A2(n_2405),
.B(n_2309),
.Y(n_2962)
);

AOI22xp5_ASAP7_75t_L g2963 ( 
.A1(n_2899),
.A2(n_2305),
.B1(n_2672),
.B2(n_2241),
.Y(n_2963)
);

OAI21x1_ASAP7_75t_L g2964 ( 
.A1(n_2811),
.A2(n_2502),
.B(n_2180),
.Y(n_2964)
);

NOR2xp33_ASAP7_75t_L g2965 ( 
.A(n_2870),
.B(n_2104),
.Y(n_2965)
);

NOR2xp33_ASAP7_75t_L g2966 ( 
.A(n_2870),
.B(n_2104),
.Y(n_2966)
);

NOR2x1_ASAP7_75t_L g2967 ( 
.A(n_2867),
.B(n_2524),
.Y(n_2967)
);

AOI21xp5_ASAP7_75t_L g2968 ( 
.A1(n_2775),
.A2(n_2405),
.B(n_2505),
.Y(n_2968)
);

A2O1A1Ixp33_ASAP7_75t_SL g2969 ( 
.A1(n_2856),
.A2(n_2807),
.B(n_2839),
.C(n_2858),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2777),
.Y(n_2970)
);

OAI22xp5_ASAP7_75t_L g2971 ( 
.A1(n_2795),
.A2(n_2780),
.B1(n_2754),
.B2(n_2774),
.Y(n_2971)
);

INVx2_ASAP7_75t_SL g2972 ( 
.A(n_2758),
.Y(n_2972)
);

NOR2xp33_ASAP7_75t_L g2973 ( 
.A(n_2870),
.B(n_2130),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2897),
.B(n_2672),
.Y(n_2974)
);

O2A1O1Ixp33_ASAP7_75t_L g2975 ( 
.A1(n_2807),
.A2(n_2288),
.B(n_2237),
.C(n_1906),
.Y(n_2975)
);

AO32x2_ASAP7_75t_L g2976 ( 
.A1(n_2774),
.A2(n_2138),
.A3(n_2130),
.B1(n_2040),
.B2(n_2672),
.Y(n_2976)
);

O2A1O1Ixp33_ASAP7_75t_L g2977 ( 
.A1(n_2839),
.A2(n_2470),
.B(n_2548),
.C(n_2322),
.Y(n_2977)
);

NOR2xp33_ASAP7_75t_L g2978 ( 
.A(n_2762),
.B(n_2138),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2843),
.B(n_2522),
.Y(n_2979)
);

CKINVDCx8_ASAP7_75t_R g2980 ( 
.A(n_2752),
.Y(n_2980)
);

BUFx6f_ASAP7_75t_L g2981 ( 
.A(n_2761),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_SL g2982 ( 
.A(n_2782),
.B(n_2538),
.Y(n_2982)
);

O2A1O1Ixp33_ASAP7_75t_L g2983 ( 
.A1(n_2877),
.A2(n_2742),
.B(n_2817),
.C(n_2890),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2907),
.B(n_2444),
.Y(n_2984)
);

INVx2_ASAP7_75t_SL g2985 ( 
.A(n_2786),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_SL g2986 ( 
.A(n_2797),
.B(n_2538),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2877),
.B(n_2444),
.Y(n_2987)
);

HB1xp67_ASAP7_75t_L g2988 ( 
.A(n_2791),
.Y(n_2988)
);

NOR2xp33_ASAP7_75t_L g2989 ( 
.A(n_2865),
.B(n_2538),
.Y(n_2989)
);

A2O1A1Ixp33_ASAP7_75t_L g2990 ( 
.A1(n_2781),
.A2(n_2318),
.B(n_2232),
.C(n_2305),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_SL g2991 ( 
.A(n_2858),
.B(n_2538),
.Y(n_2991)
);

INVx3_ASAP7_75t_L g2992 ( 
.A(n_2874),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2878),
.B(n_2454),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2879),
.B(n_2454),
.Y(n_2994)
);

OAI321xp33_ASAP7_75t_L g2995 ( 
.A1(n_2833),
.A2(n_2319),
.A3(n_2219),
.B1(n_2231),
.B2(n_2225),
.C(n_2054),
.Y(n_2995)
);

OAI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_2890),
.A2(n_2139),
.B1(n_2046),
.B2(n_2193),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2802),
.Y(n_2997)
);

OAI22xp5_ASAP7_75t_L g2998 ( 
.A1(n_2788),
.A2(n_2194),
.B1(n_2193),
.B2(n_2456),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2881),
.B(n_2456),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2864),
.B(n_2465),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2808),
.Y(n_3001)
);

INVxp67_ASAP7_75t_L g3002 ( 
.A(n_2891),
.Y(n_3002)
);

OAI21xp33_ASAP7_75t_SL g3003 ( 
.A1(n_2816),
.A2(n_2548),
.B(n_2530),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2869),
.B(n_2465),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2776),
.Y(n_3005)
);

AOI22xp5_ASAP7_75t_L g3006 ( 
.A1(n_2899),
.A2(n_2305),
.B1(n_2194),
.B2(n_2158),
.Y(n_3006)
);

AOI21xp5_ASAP7_75t_L g3007 ( 
.A1(n_2833),
.A2(n_2059),
.B(n_2598),
.Y(n_3007)
);

NOR2xp33_ASAP7_75t_L g3008 ( 
.A(n_2825),
.B(n_2415),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2888),
.B(n_2467),
.Y(n_3009)
);

A2O1A1Ixp33_ASAP7_75t_L g3010 ( 
.A1(n_2803),
.A2(n_2239),
.B(n_2100),
.C(n_2105),
.Y(n_3010)
);

AOI21xp5_ASAP7_75t_L g3011 ( 
.A1(n_2848),
.A2(n_2816),
.B(n_2798),
.Y(n_3011)
);

AOI21xp5_ASAP7_75t_L g3012 ( 
.A1(n_2848),
.A2(n_2059),
.B(n_2197),
.Y(n_3012)
);

OAI21xp5_ASAP7_75t_L g3013 ( 
.A1(n_2905),
.A2(n_2197),
.B(n_2334),
.Y(n_3013)
);

OAI22x1_ASAP7_75t_L g3014 ( 
.A1(n_2860),
.A2(n_2535),
.B1(n_2531),
.B2(n_2549),
.Y(n_3014)
);

AOI21xp5_ASAP7_75t_L g3015 ( 
.A1(n_2816),
.A2(n_2134),
.B(n_2126),
.Y(n_3015)
);

AOI21xp5_ASAP7_75t_L g3016 ( 
.A1(n_2798),
.A2(n_2136),
.B(n_2530),
.Y(n_3016)
);

OAI22xp5_ASAP7_75t_L g3017 ( 
.A1(n_2788),
.A2(n_2478),
.B1(n_2487),
.B2(n_2467),
.Y(n_3017)
);

INVx4_ASAP7_75t_L g3018 ( 
.A(n_2884),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2885),
.B(n_2478),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_SL g3020 ( 
.A(n_2868),
.B(n_2256),
.Y(n_3020)
);

AOI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2836),
.A2(n_2543),
.B(n_2349),
.Y(n_3021)
);

AOI21xp5_ASAP7_75t_L g3022 ( 
.A1(n_2836),
.A2(n_2837),
.B(n_2902),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2885),
.B(n_2487),
.Y(n_3023)
);

OAI22xp5_ASAP7_75t_L g3024 ( 
.A1(n_2789),
.A2(n_2490),
.B1(n_2493),
.B2(n_2489),
.Y(n_3024)
);

AOI21xp5_ASAP7_75t_L g3025 ( 
.A1(n_2836),
.A2(n_2543),
.B(n_2349),
.Y(n_3025)
);

AO21x1_ASAP7_75t_L g3026 ( 
.A1(n_2903),
.A2(n_2502),
.B(n_2239),
.Y(n_3026)
);

BUFx2_ASAP7_75t_L g3027 ( 
.A(n_2772),
.Y(n_3027)
);

OAI22xp5_ASAP7_75t_L g3028 ( 
.A1(n_2789),
.A2(n_2490),
.B1(n_2493),
.B2(n_2489),
.Y(n_3028)
);

AOI21xp5_ASAP7_75t_L g3029 ( 
.A1(n_2837),
.A2(n_2349),
.B(n_2331),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2827),
.Y(n_3030)
);

OAI22xp5_ASAP7_75t_L g3031 ( 
.A1(n_2863),
.A2(n_2508),
.B1(n_2511),
.B2(n_2504),
.Y(n_3031)
);

OAI21xp5_ASAP7_75t_L g3032 ( 
.A1(n_2856),
.A2(n_2334),
.B(n_2370),
.Y(n_3032)
);

OAI22xp5_ASAP7_75t_L g3033 ( 
.A1(n_2863),
.A2(n_2508),
.B1(n_2511),
.B2(n_2504),
.Y(n_3033)
);

AOI21xp5_ASAP7_75t_L g3034 ( 
.A1(n_2837),
.A2(n_2358),
.B(n_2349),
.Y(n_3034)
);

AOI21x1_ASAP7_75t_L g3035 ( 
.A1(n_2737),
.A2(n_2335),
.B(n_2330),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2887),
.B(n_2513),
.Y(n_3036)
);

AOI21xp5_ASAP7_75t_L g3037 ( 
.A1(n_2902),
.A2(n_2369),
.B(n_2358),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_2829),
.Y(n_3038)
);

O2A1O1Ixp33_ASAP7_75t_SL g3039 ( 
.A1(n_2903),
.A2(n_2089),
.B(n_2513),
.C(n_2362),
.Y(n_3039)
);

OAI22xp5_ASAP7_75t_L g3040 ( 
.A1(n_2860),
.A2(n_2089),
.B1(n_2541),
.B2(n_2522),
.Y(n_3040)
);

INVx3_ASAP7_75t_L g3041 ( 
.A(n_2874),
.Y(n_3041)
);

OA22x2_ASAP7_75t_L g3042 ( 
.A1(n_2796),
.A2(n_2362),
.B1(n_2364),
.B2(n_2324),
.Y(n_3042)
);

BUFx12f_ASAP7_75t_L g3043 ( 
.A(n_2824),
.Y(n_3043)
);

OR2x2_ASAP7_75t_L g3044 ( 
.A(n_2792),
.B(n_2849),
.Y(n_3044)
);

INVx3_ASAP7_75t_SL g3045 ( 
.A(n_2854),
.Y(n_3045)
);

O2A1O1Ixp33_ASAP7_75t_L g3046 ( 
.A1(n_2742),
.A2(n_2093),
.B(n_2542),
.C(n_2546),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2849),
.B(n_2334),
.Y(n_3047)
);

OAI22xp5_ASAP7_75t_L g3048 ( 
.A1(n_2866),
.A2(n_2737),
.B1(n_2741),
.B2(n_2852),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2880),
.B(n_2370),
.Y(n_3049)
);

NOR2xp33_ASAP7_75t_SL g3050 ( 
.A(n_2859),
.B(n_2358),
.Y(n_3050)
);

AOI21xp5_ASAP7_75t_L g3051 ( 
.A1(n_2812),
.A2(n_2379),
.B(n_2369),
.Y(n_3051)
);

A2O1A1Ixp33_ASAP7_75t_L g3052 ( 
.A1(n_2812),
.A2(n_2093),
.B(n_2364),
.C(n_2324),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2880),
.B(n_2370),
.Y(n_3053)
);

NOR2xp33_ASAP7_75t_L g3054 ( 
.A(n_2873),
.B(n_2416),
.Y(n_3054)
);

AOI21xp5_ASAP7_75t_L g3055 ( 
.A1(n_2741),
.A2(n_2379),
.B(n_2369),
.Y(n_3055)
);

AOI22xp33_ASAP7_75t_L g3056 ( 
.A1(n_2750),
.A2(n_2899),
.B1(n_2746),
.B2(n_2851),
.Y(n_3056)
);

NOR2xp33_ASAP7_75t_L g3057 ( 
.A(n_2882),
.B(n_2416),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_2908),
.B(n_2370),
.Y(n_3058)
);

AND2x2_ASAP7_75t_L g3059 ( 
.A(n_2805),
.B(n_2365),
.Y(n_3059)
);

NOR2xp33_ASAP7_75t_L g3060 ( 
.A(n_2813),
.B(n_2416),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2805),
.B(n_2370),
.Y(n_3061)
);

OAI22xp5_ASAP7_75t_L g3062 ( 
.A1(n_2852),
.A2(n_2354),
.B1(n_2336),
.B2(n_2037),
.Y(n_3062)
);

HB1xp67_ASAP7_75t_L g3063 ( 
.A(n_2893),
.Y(n_3063)
);

OAI21xp33_ASAP7_75t_L g3064 ( 
.A1(n_2794),
.A2(n_2164),
.B(n_2156),
.Y(n_3064)
);

O2A1O1Ixp33_ASAP7_75t_L g3065 ( 
.A1(n_2794),
.A2(n_2037),
.B(n_2032),
.C(n_2156),
.Y(n_3065)
);

OAI21xp33_ASAP7_75t_L g3066 ( 
.A1(n_2886),
.A2(n_2740),
.B(n_2784),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2830),
.B(n_2844),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2800),
.Y(n_3068)
);

AOI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_2886),
.A2(n_2112),
.B(n_2106),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2862),
.Y(n_3070)
);

INVx4_ASAP7_75t_L g3071 ( 
.A(n_2793),
.Y(n_3071)
);

NOR2xp33_ASAP7_75t_L g3072 ( 
.A(n_2764),
.B(n_2419),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2871),
.B(n_2354),
.Y(n_3073)
);

AOI22x1_ASAP7_75t_L g3074 ( 
.A1(n_2811),
.A2(n_2426),
.B1(n_2436),
.B2(n_2419),
.Y(n_3074)
);

BUFx2_ASAP7_75t_L g3075 ( 
.A(n_2818),
.Y(n_3075)
);

BUFx2_ASAP7_75t_L g3076 ( 
.A(n_2818),
.Y(n_3076)
);

NOR2xp33_ASAP7_75t_L g3077 ( 
.A(n_2748),
.B(n_2419),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2804),
.Y(n_3078)
);

BUFx6f_ASAP7_75t_L g3079 ( 
.A(n_2773),
.Y(n_3079)
);

AOI22xp5_ASAP7_75t_L g3080 ( 
.A1(n_2900),
.A2(n_1681),
.B1(n_1677),
.B2(n_2256),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_2872),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_SL g3082 ( 
.A(n_2949),
.B(n_2820),
.Y(n_3082)
);

AOI21xp5_ASAP7_75t_L g3083 ( 
.A1(n_2920),
.A2(n_2835),
.B(n_2906),
.Y(n_3083)
);

OAI21x1_ASAP7_75t_L g3084 ( 
.A1(n_3012),
.A2(n_2835),
.B(n_2906),
.Y(n_3084)
);

AOI21xp33_ASAP7_75t_L g3085 ( 
.A1(n_2969),
.A2(n_2819),
.B(n_2814),
.Y(n_3085)
);

INVxp67_ASAP7_75t_L g3086 ( 
.A(n_3063),
.Y(n_3086)
);

OAI21x1_ASAP7_75t_L g3087 ( 
.A1(n_3007),
.A2(n_2910),
.B(n_2909),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_3048),
.B(n_2750),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_3048),
.B(n_2750),
.Y(n_3089)
);

AOI21xp33_ASAP7_75t_L g3090 ( 
.A1(n_2945),
.A2(n_2948),
.B(n_2943),
.Y(n_3090)
);

NAND3xp33_ASAP7_75t_L g3091 ( 
.A(n_2940),
.B(n_2824),
.C(n_2820),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_SL g3092 ( 
.A(n_2952),
.B(n_2820),
.Y(n_3092)
);

OAI22xp5_ASAP7_75t_L g3093 ( 
.A1(n_2971),
.A2(n_2787),
.B1(n_2832),
.B2(n_2822),
.Y(n_3093)
);

BUFx2_ASAP7_75t_L g3094 ( 
.A(n_2946),
.Y(n_3094)
);

OAI21x1_ASAP7_75t_SL g3095 ( 
.A1(n_2916),
.A2(n_2842),
.B(n_2840),
.Y(n_3095)
);

CKINVDCx20_ASAP7_75t_R g3096 ( 
.A(n_3045),
.Y(n_3096)
);

OAI21x1_ASAP7_75t_L g3097 ( 
.A1(n_2944),
.A2(n_2850),
.B(n_2846),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2915),
.B(n_2746),
.Y(n_3098)
);

AOI21xp5_ASAP7_75t_L g3099 ( 
.A1(n_2955),
.A2(n_2783),
.B(n_2757),
.Y(n_3099)
);

AO21x2_ASAP7_75t_L g3100 ( 
.A1(n_3016),
.A2(n_3069),
.B(n_2918),
.Y(n_3100)
);

AOI21xp5_ASAP7_75t_L g3101 ( 
.A1(n_2941),
.A2(n_2757),
.B(n_2755),
.Y(n_3101)
);

OAI21x1_ASAP7_75t_L g3102 ( 
.A1(n_3035),
.A2(n_2853),
.B(n_2828),
.Y(n_3102)
);

AOI21xp5_ASAP7_75t_L g3103 ( 
.A1(n_2995),
.A2(n_2755),
.B(n_2749),
.Y(n_3103)
);

AO31x2_ASAP7_75t_L g3104 ( 
.A1(n_3026),
.A2(n_2838),
.A3(n_2845),
.B(n_2841),
.Y(n_3104)
);

OR2x2_ASAP7_75t_L g3105 ( 
.A(n_3044),
.B(n_2875),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2922),
.B(n_2746),
.Y(n_3106)
);

OAI21x1_ASAP7_75t_L g3107 ( 
.A1(n_2928),
.A2(n_2828),
.B(n_2821),
.Y(n_3107)
);

NAND2x1_ASAP7_75t_L g3108 ( 
.A(n_2912),
.B(n_2913),
.Y(n_3108)
);

AOI211x1_ASAP7_75t_L g3109 ( 
.A1(n_3067),
.A2(n_32),
.B(n_29),
.C(n_30),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_3081),
.Y(n_3110)
);

OAI21x1_ASAP7_75t_L g3111 ( 
.A1(n_3055),
.A2(n_2847),
.B(n_2821),
.Y(n_3111)
);

O2A1O1Ixp5_ASAP7_75t_L g3112 ( 
.A1(n_2927),
.A2(n_2925),
.B(n_2926),
.C(n_2932),
.Y(n_3112)
);

BUFx2_ASAP7_75t_L g3113 ( 
.A(n_3027),
.Y(n_3113)
);

AOI211x1_ASAP7_75t_L g3114 ( 
.A1(n_2971),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2950),
.B(n_2746),
.Y(n_3115)
);

O2A1O1Ixp5_ASAP7_75t_L g3116 ( 
.A1(n_2927),
.A2(n_2841),
.B(n_2845),
.C(n_2838),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_3005),
.Y(n_3117)
);

OAI21x1_ASAP7_75t_L g3118 ( 
.A1(n_2964),
.A2(n_2883),
.B(n_2847),
.Y(n_3118)
);

NAND2x1p5_ASAP7_75t_L g3119 ( 
.A(n_2967),
.B(n_2743),
.Y(n_3119)
);

INVxp67_ASAP7_75t_L g3120 ( 
.A(n_2934),
.Y(n_3120)
);

OAI21xp5_ASAP7_75t_L g3121 ( 
.A1(n_2990),
.A2(n_2904),
.B(n_2883),
.Y(n_3121)
);

INVxp67_ASAP7_75t_L g3122 ( 
.A(n_2988),
.Y(n_3122)
);

INVx2_ASAP7_75t_SL g3123 ( 
.A(n_2981),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_3066),
.B(n_2904),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2935),
.B(n_2904),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2939),
.B(n_2904),
.Y(n_3126)
);

OAI22xp5_ASAP7_75t_L g3127 ( 
.A1(n_2924),
.A2(n_2931),
.B1(n_2933),
.B2(n_2942),
.Y(n_3127)
);

AOI21xp5_ASAP7_75t_L g3128 ( 
.A1(n_2995),
.A2(n_2426),
.B(n_2419),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_3068),
.B(n_2787),
.Y(n_3129)
);

INVx2_ASAP7_75t_SL g3130 ( 
.A(n_2981),
.Y(n_3130)
);

OAI21x1_ASAP7_75t_L g3131 ( 
.A1(n_2956),
.A2(n_2032),
.B(n_1581),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_3078),
.Y(n_3132)
);

AO21x2_ASAP7_75t_L g3133 ( 
.A1(n_3039),
.A2(n_2164),
.B(n_1614),
.Y(n_3133)
);

AOI21xp5_ASAP7_75t_L g3134 ( 
.A1(n_2961),
.A2(n_2436),
.B(n_2426),
.Y(n_3134)
);

OAI22xp5_ASAP7_75t_L g3135 ( 
.A1(n_2924),
.A2(n_2787),
.B1(n_2766),
.B2(n_2790),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_SL g3136 ( 
.A(n_2958),
.B(n_2874),
.Y(n_3136)
);

AOI21xp5_ASAP7_75t_L g3137 ( 
.A1(n_3010),
.A2(n_2436),
.B(n_2889),
.Y(n_3137)
);

AOI21xp5_ASAP7_75t_L g3138 ( 
.A1(n_3037),
.A2(n_2112),
.B(n_2106),
.Y(n_3138)
);

INVxp67_ASAP7_75t_L g3139 ( 
.A(n_2929),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2917),
.B(n_2876),
.Y(n_3140)
);

OAI21xp5_ASAP7_75t_L g3141 ( 
.A1(n_3015),
.A2(n_2155),
.B(n_2409),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_3011),
.B(n_2876),
.Y(n_3142)
);

AND2x2_ASAP7_75t_L g3143 ( 
.A(n_2937),
.B(n_2876),
.Y(n_3143)
);

BUFx2_ASAP7_75t_L g3144 ( 
.A(n_3075),
.Y(n_3144)
);

A2O1A1Ixp33_ASAP7_75t_L g3145 ( 
.A1(n_2919),
.A2(n_2421),
.B(n_2506),
.C(n_2503),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2923),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_2936),
.B(n_2773),
.Y(n_3147)
);

OAI22xp5_ASAP7_75t_L g3148 ( 
.A1(n_2933),
.A2(n_2799),
.B1(n_2778),
.B2(n_2421),
.Y(n_3148)
);

O2A1O1Ixp5_ASAP7_75t_L g3149 ( 
.A1(n_2959),
.A2(n_2503),
.B(n_2506),
.C(n_2155),
.Y(n_3149)
);

OAI21xp5_ASAP7_75t_L g3150 ( 
.A1(n_2962),
.A2(n_2155),
.B(n_1624),
.Y(n_3150)
);

AOI21xp5_ASAP7_75t_L g3151 ( 
.A1(n_3032),
.A2(n_2799),
.B(n_2778),
.Y(n_3151)
);

AOI21xp5_ASAP7_75t_L g3152 ( 
.A1(n_3032),
.A2(n_2799),
.B(n_2778),
.Y(n_3152)
);

BUFx2_ASAP7_75t_L g3153 ( 
.A(n_3076),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2929),
.B(n_35),
.Y(n_3154)
);

INVx3_ASAP7_75t_L g3155 ( 
.A(n_3079),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3019),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2953),
.B(n_2943),
.Y(n_3157)
);

AOI221x1_ASAP7_75t_L g3158 ( 
.A1(n_2930),
.A2(n_3034),
.B1(n_3029),
.B2(n_3014),
.C(n_3054),
.Y(n_3158)
);

BUFx6f_ASAP7_75t_L g3159 ( 
.A(n_2981),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_3023),
.B(n_35),
.Y(n_3160)
);

INVx4_ASAP7_75t_L g3161 ( 
.A(n_3071),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_3036),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_2954),
.B(n_37),
.Y(n_3163)
);

CKINVDCx14_ASAP7_75t_R g3164 ( 
.A(n_3043),
.Y(n_3164)
);

AOI21xp5_ASAP7_75t_L g3165 ( 
.A1(n_3013),
.A2(n_2035),
.B(n_1495),
.Y(n_3165)
);

OAI21x1_ASAP7_75t_L g3166 ( 
.A1(n_2968),
.A2(n_1495),
.B(n_1475),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_3047),
.B(n_38),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_2938),
.Y(n_3168)
);

A2O1A1Ixp33_ASAP7_75t_L g3169 ( 
.A1(n_3003),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_3169)
);

AOI21xp5_ASAP7_75t_L g3170 ( 
.A1(n_2977),
.A2(n_2035),
.B(n_1495),
.Y(n_3170)
);

OAI21x1_ASAP7_75t_L g3171 ( 
.A1(n_3065),
.A2(n_1546),
.B(n_1475),
.Y(n_3171)
);

AOI221xp5_ASAP7_75t_L g3172 ( 
.A1(n_2983),
.A2(n_1596),
.B1(n_1600),
.B2(n_1568),
.C(n_1557),
.Y(n_3172)
);

OAI21xp5_ASAP7_75t_L g3173 ( 
.A1(n_2975),
.A2(n_1654),
.B(n_1546),
.Y(n_3173)
);

OAI22x1_ASAP7_75t_L g3174 ( 
.A1(n_3002),
.A2(n_42),
.B1(n_39),
.B2(n_41),
.Y(n_3174)
);

AOI21x1_ASAP7_75t_L g3175 ( 
.A1(n_3021),
.A2(n_1591),
.B(n_1575),
.Y(n_3175)
);

AO21x1_ASAP7_75t_L g3176 ( 
.A1(n_2991),
.A2(n_43),
.B(n_44),
.Y(n_3176)
);

AND2x4_ASAP7_75t_L g3177 ( 
.A(n_3022),
.B(n_2035),
.Y(n_3177)
);

BUFx3_ASAP7_75t_L g3178 ( 
.A(n_2972),
.Y(n_3178)
);

AO31x2_ASAP7_75t_L g3179 ( 
.A1(n_3062),
.A2(n_1454),
.A3(n_2256),
.B(n_1654),
.Y(n_3179)
);

OAI22xp5_ASAP7_75t_L g3180 ( 
.A1(n_3056),
.A2(n_2963),
.B1(n_3042),
.B2(n_3058),
.Y(n_3180)
);

AOI21x1_ASAP7_75t_L g3181 ( 
.A1(n_3025),
.A2(n_1645),
.B(n_1654),
.Y(n_3181)
);

OAI21xp5_ASAP7_75t_L g3182 ( 
.A1(n_3006),
.A2(n_1654),
.B(n_1645),
.Y(n_3182)
);

OAI21x1_ASAP7_75t_L g3183 ( 
.A1(n_3017),
.A2(n_1645),
.B(n_1456),
.Y(n_3183)
);

AOI21xp5_ASAP7_75t_L g3184 ( 
.A1(n_2986),
.A2(n_1568),
.B(n_1557),
.Y(n_3184)
);

OAI21x1_ASAP7_75t_L g3185 ( 
.A1(n_3017),
.A2(n_1456),
.B(n_1449),
.Y(n_3185)
);

OAI21x1_ASAP7_75t_L g3186 ( 
.A1(n_3024),
.A2(n_1456),
.B(n_1449),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2970),
.Y(n_3187)
);

AO31x2_ASAP7_75t_L g3188 ( 
.A1(n_3062),
.A2(n_1454),
.A3(n_1654),
.B(n_46),
.Y(n_3188)
);

OAI21x1_ASAP7_75t_SL g3189 ( 
.A1(n_3046),
.A2(n_44),
.B(n_45),
.Y(n_3189)
);

OAI21xp5_ASAP7_75t_L g3190 ( 
.A1(n_3064),
.A2(n_1654),
.B(n_1449),
.Y(n_3190)
);

OAI21xp5_ASAP7_75t_L g3191 ( 
.A1(n_2998),
.A2(n_1504),
.B(n_45),
.Y(n_3191)
);

OAI21x1_ASAP7_75t_L g3192 ( 
.A1(n_3024),
.A2(n_1568),
.B(n_1557),
.Y(n_3192)
);

OAI21x1_ASAP7_75t_L g3193 ( 
.A1(n_3028),
.A2(n_1596),
.B(n_1568),
.Y(n_3193)
);

OAI21x1_ASAP7_75t_L g3194 ( 
.A1(n_3028),
.A2(n_1600),
.B(n_1596),
.Y(n_3194)
);

AOI21xp33_ASAP7_75t_L g3195 ( 
.A1(n_2998),
.A2(n_46),
.B(n_47),
.Y(n_3195)
);

O2A1O1Ixp5_ASAP7_75t_L g3196 ( 
.A1(n_2982),
.A2(n_50),
.B(n_47),
.C(n_49),
.Y(n_3196)
);

A2O1A1Ixp33_ASAP7_75t_L g3197 ( 
.A1(n_3080),
.A2(n_51),
.B(n_49),
.C(n_50),
.Y(n_3197)
);

OAI21x1_ASAP7_75t_L g3198 ( 
.A1(n_3074),
.A2(n_1600),
.B(n_1596),
.Y(n_3198)
);

AND2x2_ASAP7_75t_L g3199 ( 
.A(n_3059),
.B(n_51),
.Y(n_3199)
);

OAI21xp5_ASAP7_75t_L g3200 ( 
.A1(n_3052),
.A2(n_3033),
.B(n_3031),
.Y(n_3200)
);

OAI21x1_ASAP7_75t_SL g3201 ( 
.A1(n_2974),
.A2(n_52),
.B(n_54),
.Y(n_3201)
);

AOI21xp5_ASAP7_75t_L g3202 ( 
.A1(n_3051),
.A2(n_1603),
.B(n_1600),
.Y(n_3202)
);

AND2x2_ASAP7_75t_L g3203 ( 
.A(n_2914),
.B(n_52),
.Y(n_3203)
);

AO22x2_ASAP7_75t_L g3204 ( 
.A1(n_3049),
.A2(n_58),
.B1(n_55),
.B2(n_56),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3053),
.B(n_60),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2997),
.Y(n_3206)
);

NOR2xp67_ASAP7_75t_SL g3207 ( 
.A(n_2980),
.B(n_1603),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3001),
.Y(n_3208)
);

BUFx2_ASAP7_75t_L g3209 ( 
.A(n_2914),
.Y(n_3209)
);

AO31x2_ASAP7_75t_L g3210 ( 
.A1(n_3031),
.A2(n_62),
.A3(n_60),
.B(n_61),
.Y(n_3210)
);

OA22x2_ASAP7_75t_L g3211 ( 
.A1(n_3020),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2987),
.B(n_3030),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_3038),
.B(n_64),
.Y(n_3213)
);

OAI22xp5_ASAP7_75t_L g3214 ( 
.A1(n_3042),
.A2(n_67),
.B1(n_64),
.B2(n_65),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_L g3215 ( 
.A(n_3070),
.B(n_65),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_3000),
.B(n_68),
.Y(n_3216)
);

OAI21x1_ASAP7_75t_L g3217 ( 
.A1(n_3033),
.A2(n_1615),
.B(n_1603),
.Y(n_3217)
);

A2O1A1Ixp33_ASAP7_75t_L g3218 ( 
.A1(n_2957),
.A2(n_71),
.B(n_68),
.C(n_70),
.Y(n_3218)
);

OAI21x1_ASAP7_75t_L g3219 ( 
.A1(n_3040),
.A2(n_1615),
.B(n_1603),
.Y(n_3219)
);

AO21x1_ASAP7_75t_L g3220 ( 
.A1(n_3060),
.A2(n_70),
.B(n_71),
.Y(n_3220)
);

OAI21x1_ASAP7_75t_L g3221 ( 
.A1(n_3040),
.A2(n_1615),
.B(n_1603),
.Y(n_3221)
);

OAI21xp5_ASAP7_75t_L g3222 ( 
.A1(n_2996),
.A2(n_1504),
.B(n_72),
.Y(n_3222)
);

INVx5_ASAP7_75t_L g3223 ( 
.A(n_3079),
.Y(n_3223)
);

OAI21x1_ASAP7_75t_L g3224 ( 
.A1(n_2996),
.A2(n_1650),
.B(n_1641),
.Y(n_3224)
);

NAND2x1p5_ASAP7_75t_L g3225 ( 
.A(n_3071),
.B(n_1641),
.Y(n_3225)
);

OA21x2_ASAP7_75t_L g3226 ( 
.A1(n_3061),
.A2(n_72),
.B(n_73),
.Y(n_3226)
);

OAI21x1_ASAP7_75t_L g3227 ( 
.A1(n_3073),
.A2(n_1650),
.B(n_1641),
.Y(n_3227)
);

AOI21xp5_ASAP7_75t_L g3228 ( 
.A1(n_2960),
.A2(n_1652),
.B(n_1650),
.Y(n_3228)
);

HB1xp67_ASAP7_75t_L g3229 ( 
.A(n_2979),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_3004),
.B(n_2984),
.Y(n_3230)
);

AO21x1_ASAP7_75t_L g3231 ( 
.A1(n_3009),
.A2(n_73),
.B(n_74),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_2999),
.B(n_74),
.Y(n_3232)
);

INVx3_ASAP7_75t_L g3233 ( 
.A(n_2992),
.Y(n_3233)
);

NOR2x1_ASAP7_75t_L g3234 ( 
.A(n_2947),
.B(n_961),
.Y(n_3234)
);

INVx2_ASAP7_75t_L g3235 ( 
.A(n_2992),
.Y(n_3235)
);

OR2x6_ASAP7_75t_L g3236 ( 
.A(n_3018),
.B(n_1650),
.Y(n_3236)
);

OAI22xp5_ASAP7_75t_L g3237 ( 
.A1(n_2985),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_3237)
);

OAI21x1_ASAP7_75t_L g3238 ( 
.A1(n_2993),
.A2(n_2994),
.B(n_3041),
.Y(n_3238)
);

AOI21xp5_ASAP7_75t_L g3239 ( 
.A1(n_2965),
.A2(n_1652),
.B(n_1650),
.Y(n_3239)
);

OAI21xp5_ASAP7_75t_L g3240 ( 
.A1(n_2978),
.A2(n_1504),
.B(n_77),
.Y(n_3240)
);

INVx2_ASAP7_75t_L g3241 ( 
.A(n_2976),
.Y(n_3241)
);

OAI21xp5_ASAP7_75t_L g3242 ( 
.A1(n_2966),
.A2(n_1504),
.B(n_80),
.Y(n_3242)
);

AND2x2_ASAP7_75t_L g3243 ( 
.A(n_3008),
.B(n_80),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_3057),
.B(n_81),
.Y(n_3244)
);

OR2x6_ASAP7_75t_L g3245 ( 
.A(n_3018),
.B(n_1652),
.Y(n_3245)
);

OA21x2_ASAP7_75t_L g3246 ( 
.A1(n_2973),
.A2(n_81),
.B(n_82),
.Y(n_3246)
);

HB1xp67_ASAP7_75t_L g3247 ( 
.A(n_3077),
.Y(n_3247)
);

INVx6_ASAP7_75t_SL g3248 ( 
.A(n_2951),
.Y(n_3248)
);

AND2x4_ASAP7_75t_L g3249 ( 
.A(n_2989),
.B(n_308),
.Y(n_3249)
);

AOI21xp33_ASAP7_75t_L g3250 ( 
.A1(n_2921),
.A2(n_83),
.B(n_84),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_3072),
.B(n_83),
.Y(n_3251)
);

O2A1O1Ixp33_ASAP7_75t_L g3252 ( 
.A1(n_3050),
.A2(n_86),
.B(n_84),
.C(n_85),
.Y(n_3252)
);

OAI21x1_ASAP7_75t_L g3253 ( 
.A1(n_2976),
.A2(n_1653),
.B(n_310),
.Y(n_3253)
);

OAI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_2920),
.A2(n_1504),
.B(n_85),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_SL g3255 ( 
.A(n_2949),
.B(n_1470),
.Y(n_3255)
);

OAI21xp5_ASAP7_75t_L g3256 ( 
.A1(n_3254),
.A2(n_86),
.B(n_89),
.Y(n_3256)
);

AOI21xp5_ASAP7_75t_L g3257 ( 
.A1(n_3254),
.A2(n_1467),
.B(n_1447),
.Y(n_3257)
);

AOI21x1_ASAP7_75t_L g3258 ( 
.A1(n_3234),
.A2(n_89),
.B(n_91),
.Y(n_3258)
);

AOI21xp5_ASAP7_75t_L g3259 ( 
.A1(n_3170),
.A2(n_1467),
.B(n_1447),
.Y(n_3259)
);

OAI21xp5_ASAP7_75t_L g3260 ( 
.A1(n_3169),
.A2(n_92),
.B(n_93),
.Y(n_3260)
);

OAI22xp5_ASAP7_75t_L g3261 ( 
.A1(n_3127),
.A2(n_1064),
.B1(n_1133),
.B2(n_961),
.Y(n_3261)
);

AOI22xp5_ASAP7_75t_L g3262 ( 
.A1(n_3127),
.A2(n_1498),
.B1(n_1470),
.B2(n_1497),
.Y(n_3262)
);

AOI21xp5_ASAP7_75t_L g3263 ( 
.A1(n_3228),
.A2(n_1491),
.B(n_1470),
.Y(n_3263)
);

OAI21x1_ASAP7_75t_L g3264 ( 
.A1(n_3198),
.A2(n_322),
.B(n_321),
.Y(n_3264)
);

OAI21xp5_ASAP7_75t_L g3265 ( 
.A1(n_3112),
.A2(n_93),
.B(n_94),
.Y(n_3265)
);

OA21x2_ASAP7_75t_L g3266 ( 
.A1(n_3158),
.A2(n_95),
.B(n_96),
.Y(n_3266)
);

BUFx10_ASAP7_75t_L g3267 ( 
.A(n_3159),
.Y(n_3267)
);

OAI21x1_ASAP7_75t_L g3268 ( 
.A1(n_3224),
.A2(n_326),
.B(n_324),
.Y(n_3268)
);

OAI21x1_ASAP7_75t_L g3269 ( 
.A1(n_3227),
.A2(n_331),
.B(n_327),
.Y(n_3269)
);

AOI21x1_ASAP7_75t_SL g3270 ( 
.A1(n_3142),
.A2(n_95),
.B(n_97),
.Y(n_3270)
);

OR2x2_ASAP7_75t_L g3271 ( 
.A(n_3115),
.B(n_98),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_3117),
.Y(n_3272)
);

OAI22xp5_ASAP7_75t_L g3273 ( 
.A1(n_3197),
.A2(n_1064),
.B1(n_102),
.B2(n_99),
.Y(n_3273)
);

AND2x2_ASAP7_75t_L g3274 ( 
.A(n_3094),
.B(n_99),
.Y(n_3274)
);

OAI21x1_ASAP7_75t_L g3275 ( 
.A1(n_3185),
.A2(n_335),
.B(n_334),
.Y(n_3275)
);

AO32x2_ASAP7_75t_L g3276 ( 
.A1(n_3093),
.A2(n_101),
.A3(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_3276)
);

BUFx2_ASAP7_75t_L g3277 ( 
.A(n_3247),
.Y(n_3277)
);

OAI21x1_ASAP7_75t_L g3278 ( 
.A1(n_3186),
.A2(n_338),
.B(n_337),
.Y(n_3278)
);

NAND3x1_ASAP7_75t_L g3279 ( 
.A(n_3240),
.B(n_3154),
.C(n_3157),
.Y(n_3279)
);

OAI22x1_ASAP7_75t_L g3280 ( 
.A1(n_3120),
.A2(n_107),
.B1(n_101),
.B2(n_104),
.Y(n_3280)
);

AOI21x1_ASAP7_75t_L g3281 ( 
.A1(n_3082),
.A2(n_108),
.B(n_109),
.Y(n_3281)
);

O2A1O1Ixp33_ASAP7_75t_L g3282 ( 
.A1(n_3218),
.A2(n_112),
.B(n_108),
.C(n_109),
.Y(n_3282)
);

NAND3xp33_ASAP7_75t_L g3283 ( 
.A(n_3090),
.B(n_1064),
.C(n_1023),
.Y(n_3283)
);

OA21x2_ASAP7_75t_L g3284 ( 
.A1(n_3090),
.A2(n_112),
.B(n_113),
.Y(n_3284)
);

NOR2x1_ASAP7_75t_R g3285 ( 
.A(n_3161),
.B(n_780),
.Y(n_3285)
);

BUFx4_ASAP7_75t_SL g3286 ( 
.A(n_3096),
.Y(n_3286)
);

NOR2xp33_ASAP7_75t_SL g3287 ( 
.A(n_3161),
.B(n_780),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_3156),
.B(n_114),
.Y(n_3288)
);

INVxp67_ASAP7_75t_L g3289 ( 
.A(n_3229),
.Y(n_3289)
);

AOI221xp5_ASAP7_75t_L g3290 ( 
.A1(n_3237),
.A2(n_116),
.B1(n_117),
.B2(n_119),
.C(n_120),
.Y(n_3290)
);

OAI21x1_ASAP7_75t_L g3291 ( 
.A1(n_3192),
.A2(n_3194),
.B(n_3193),
.Y(n_3291)
);

BUFx3_ASAP7_75t_L g3292 ( 
.A(n_3159),
.Y(n_3292)
);

OAI21x1_ASAP7_75t_L g3293 ( 
.A1(n_3219),
.A2(n_343),
.B(n_340),
.Y(n_3293)
);

AND2x2_ASAP7_75t_L g3294 ( 
.A(n_3113),
.B(n_117),
.Y(n_3294)
);

AOI21xp5_ASAP7_75t_L g3295 ( 
.A1(n_3165),
.A2(n_1497),
.B(n_1491),
.Y(n_3295)
);

A2O1A1Ixp33_ASAP7_75t_L g3296 ( 
.A1(n_3252),
.A2(n_122),
.B(n_119),
.C(n_120),
.Y(n_3296)
);

CKINVDCx11_ASAP7_75t_R g3297 ( 
.A(n_3159),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_3162),
.B(n_123),
.Y(n_3298)
);

AOI22xp5_ASAP7_75t_L g3299 ( 
.A1(n_3093),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_3299)
);

NOR2x1_ASAP7_75t_R g3300 ( 
.A(n_3248),
.B(n_780),
.Y(n_3300)
);

OAI21xp5_ASAP7_75t_L g3301 ( 
.A1(n_3091),
.A2(n_124),
.B(n_126),
.Y(n_3301)
);

AOI21xp5_ASAP7_75t_L g3302 ( 
.A1(n_3100),
.A2(n_1497),
.B(n_1491),
.Y(n_3302)
);

OAI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_3240),
.A2(n_127),
.B(n_128),
.Y(n_3303)
);

AOI21xp5_ASAP7_75t_L g3304 ( 
.A1(n_3100),
.A2(n_1498),
.B(n_1023),
.Y(n_3304)
);

AOI22xp33_ASAP7_75t_SL g3305 ( 
.A1(n_3242),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_3305)
);

AOI22xp5_ASAP7_75t_L g3306 ( 
.A1(n_3135),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_3306)
);

AO31x2_ASAP7_75t_L g3307 ( 
.A1(n_3214),
.A2(n_133),
.A3(n_134),
.B(n_135),
.Y(n_3307)
);

A2O1A1Ixp33_ASAP7_75t_L g3308 ( 
.A1(n_3242),
.A2(n_134),
.B(n_136),
.C(n_137),
.Y(n_3308)
);

OA21x2_ASAP7_75t_L g3309 ( 
.A1(n_3097),
.A2(n_136),
.B(n_137),
.Y(n_3309)
);

AND2x4_ASAP7_75t_L g3310 ( 
.A(n_3122),
.B(n_138),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3086),
.B(n_139),
.Y(n_3311)
);

OAI21x1_ASAP7_75t_L g3312 ( 
.A1(n_3221),
.A2(n_3217),
.B(n_3101),
.Y(n_3312)
);

INVx3_ASAP7_75t_L g3313 ( 
.A(n_3119),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_3132),
.Y(n_3314)
);

AO31x2_ASAP7_75t_L g3315 ( 
.A1(n_3214),
.A2(n_140),
.A3(n_141),
.B(n_143),
.Y(n_3315)
);

AOI21xp5_ASAP7_75t_L g3316 ( 
.A1(n_3222),
.A2(n_1498),
.B(n_1023),
.Y(n_3316)
);

O2A1O1Ixp33_ASAP7_75t_L g3317 ( 
.A1(n_3237),
.A2(n_140),
.B(n_141),
.C(n_144),
.Y(n_3317)
);

CKINVDCx20_ASAP7_75t_R g3318 ( 
.A(n_3164),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_3222),
.A2(n_1498),
.B(n_1023),
.Y(n_3319)
);

INVx4_ASAP7_75t_SL g3320 ( 
.A(n_3210),
.Y(n_3320)
);

AOI22xp5_ASAP7_75t_L g3321 ( 
.A1(n_3135),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3110),
.Y(n_3322)
);

AO31x2_ASAP7_75t_L g3323 ( 
.A1(n_3241),
.A2(n_147),
.A3(n_149),
.B(n_151),
.Y(n_3323)
);

AOI21xp5_ASAP7_75t_L g3324 ( 
.A1(n_3190),
.A2(n_1023),
.B(n_780),
.Y(n_3324)
);

CKINVDCx5p33_ASAP7_75t_R g3325 ( 
.A(n_3248),
.Y(n_3325)
);

OAI21x1_ASAP7_75t_L g3326 ( 
.A1(n_3083),
.A2(n_347),
.B(n_346),
.Y(n_3326)
);

AOI22xp5_ASAP7_75t_L g3327 ( 
.A1(n_3180),
.A2(n_780),
.B1(n_152),
.B2(n_153),
.Y(n_3327)
);

A2O1A1Ixp33_ASAP7_75t_L g3328 ( 
.A1(n_3191),
.A2(n_147),
.B(n_154),
.C(n_156),
.Y(n_3328)
);

A2O1A1Ixp33_ASAP7_75t_L g3329 ( 
.A1(n_3191),
.A2(n_156),
.B(n_157),
.C(n_158),
.Y(n_3329)
);

NAND3xp33_ASAP7_75t_L g3330 ( 
.A(n_3109),
.B(n_780),
.C(n_159),
.Y(n_3330)
);

BUFx3_ASAP7_75t_L g3331 ( 
.A(n_3178),
.Y(n_3331)
);

NOR2xp33_ASAP7_75t_L g3332 ( 
.A(n_3092),
.B(n_159),
.Y(n_3332)
);

OAI21xp5_ASAP7_75t_L g3333 ( 
.A1(n_3255),
.A2(n_160),
.B(n_161),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3108),
.Y(n_3334)
);

AO31x2_ASAP7_75t_L g3335 ( 
.A1(n_3231),
.A2(n_162),
.A3(n_163),
.B(n_165),
.Y(n_3335)
);

OR2x6_ASAP7_75t_L g3336 ( 
.A(n_3099),
.B(n_3121),
.Y(n_3336)
);

AO31x2_ASAP7_75t_L g3337 ( 
.A1(n_3137),
.A2(n_165),
.A3(n_167),
.B(n_169),
.Y(n_3337)
);

OAI21x1_ASAP7_75t_L g3338 ( 
.A1(n_3134),
.A2(n_355),
.B(n_350),
.Y(n_3338)
);

AOI21xp5_ASAP7_75t_L g3339 ( 
.A1(n_3190),
.A2(n_167),
.B(n_169),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_3157),
.B(n_170),
.Y(n_3340)
);

AOI21xp5_ASAP7_75t_L g3341 ( 
.A1(n_3200),
.A2(n_170),
.B(n_171),
.Y(n_3341)
);

HB1xp67_ASAP7_75t_L g3342 ( 
.A(n_3139),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_SL g3343 ( 
.A(n_3142),
.B(n_356),
.Y(n_3343)
);

AND2x2_ASAP7_75t_L g3344 ( 
.A(n_3144),
.B(n_3153),
.Y(n_3344)
);

AOI21xp5_ASAP7_75t_L g3345 ( 
.A1(n_3200),
.A2(n_171),
.B(n_173),
.Y(n_3345)
);

BUFx6f_ASAP7_75t_L g3346 ( 
.A(n_3223),
.Y(n_3346)
);

INVx3_ASAP7_75t_L g3347 ( 
.A(n_3119),
.Y(n_3347)
);

OAI21x1_ASAP7_75t_L g3348 ( 
.A1(n_3084),
.A2(n_366),
.B(n_361),
.Y(n_3348)
);

AOI21xp5_ASAP7_75t_L g3349 ( 
.A1(n_3141),
.A2(n_173),
.B(n_174),
.Y(n_3349)
);

NAND3xp33_ASAP7_75t_SL g3350 ( 
.A(n_3220),
.B(n_174),
.C(n_175),
.Y(n_3350)
);

AOI21xp5_ASAP7_75t_L g3351 ( 
.A1(n_3141),
.A2(n_175),
.B(n_176),
.Y(n_3351)
);

AOI21xp5_ASAP7_75t_L g3352 ( 
.A1(n_3128),
.A2(n_176),
.B(n_177),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_3105),
.Y(n_3353)
);

NAND3xp33_ASAP7_75t_L g3354 ( 
.A(n_3250),
.B(n_178),
.C(n_179),
.Y(n_3354)
);

O2A1O1Ixp33_ASAP7_75t_SL g3355 ( 
.A1(n_3250),
.A2(n_178),
.B(n_179),
.C(n_180),
.Y(n_3355)
);

AOI21xp5_ASAP7_75t_L g3356 ( 
.A1(n_3121),
.A2(n_180),
.B(n_182),
.Y(n_3356)
);

OR2x2_ASAP7_75t_L g3357 ( 
.A(n_3115),
.B(n_184),
.Y(n_3357)
);

INVx3_ASAP7_75t_L g3358 ( 
.A(n_3235),
.Y(n_3358)
);

OAI21x1_ASAP7_75t_L g3359 ( 
.A1(n_3087),
.A2(n_370),
.B(n_369),
.Y(n_3359)
);

A2O1A1Ixp33_ASAP7_75t_L g3360 ( 
.A1(n_3196),
.A2(n_184),
.B(n_185),
.C(n_186),
.Y(n_3360)
);

AO221x2_ASAP7_75t_L g3361 ( 
.A1(n_3174),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.C(n_188),
.Y(n_3361)
);

AOI21xp5_ASAP7_75t_L g3362 ( 
.A1(n_3173),
.A2(n_189),
.B(n_190),
.Y(n_3362)
);

INVxp67_ASAP7_75t_L g3363 ( 
.A(n_3147),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3209),
.B(n_189),
.Y(n_3364)
);

AO21x1_ASAP7_75t_L g3365 ( 
.A1(n_3085),
.A2(n_190),
.B(n_192),
.Y(n_3365)
);

AOI21xp5_ASAP7_75t_L g3366 ( 
.A1(n_3173),
.A2(n_193),
.B(n_195),
.Y(n_3366)
);

OR2x2_ASAP7_75t_L g3367 ( 
.A(n_3088),
.B(n_196),
.Y(n_3367)
);

O2A1O1Ixp33_ASAP7_75t_L g3368 ( 
.A1(n_3195),
.A2(n_197),
.B(n_198),
.C(n_199),
.Y(n_3368)
);

OAI21xp5_ASAP7_75t_L g3369 ( 
.A1(n_3085),
.A2(n_197),
.B(n_200),
.Y(n_3369)
);

AND2x2_ASAP7_75t_L g3370 ( 
.A(n_3143),
.B(n_200),
.Y(n_3370)
);

OAI22x1_ASAP7_75t_L g3371 ( 
.A1(n_3088),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_3371)
);

AOI21xp5_ASAP7_75t_L g3372 ( 
.A1(n_3172),
.A2(n_202),
.B(n_203),
.Y(n_3372)
);

INVx3_ASAP7_75t_L g3373 ( 
.A(n_3233),
.Y(n_3373)
);

AND2x4_ASAP7_75t_L g3374 ( 
.A(n_3177),
.B(n_204),
.Y(n_3374)
);

INVx2_ASAP7_75t_L g3375 ( 
.A(n_3187),
.Y(n_3375)
);

OA21x2_ASAP7_75t_L g3376 ( 
.A1(n_3140),
.A2(n_205),
.B(n_206),
.Y(n_3376)
);

INVx3_ASAP7_75t_L g3377 ( 
.A(n_3233),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_3212),
.B(n_206),
.Y(n_3378)
);

NOR2x1_ASAP7_75t_L g3379 ( 
.A(n_3140),
.B(n_207),
.Y(n_3379)
);

NAND3xp33_ASAP7_75t_L g3380 ( 
.A(n_3114),
.B(n_3195),
.C(n_3167),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3212),
.B(n_208),
.Y(n_3381)
);

NOR2xp67_ASAP7_75t_L g3382 ( 
.A(n_3206),
.B(n_209),
.Y(n_3382)
);

AOI21xp5_ASAP7_75t_SL g3383 ( 
.A1(n_3246),
.A2(n_446),
.B(n_445),
.Y(n_3383)
);

NOR2xp67_ASAP7_75t_L g3384 ( 
.A(n_3208),
.B(n_209),
.Y(n_3384)
);

A2O1A1Ixp33_ASAP7_75t_L g3385 ( 
.A1(n_3089),
.A2(n_210),
.B(n_211),
.C(n_212),
.Y(n_3385)
);

AOI21xp5_ASAP7_75t_L g3386 ( 
.A1(n_3103),
.A2(n_210),
.B(n_213),
.Y(n_3386)
);

OAI22x1_ASAP7_75t_L g3387 ( 
.A1(n_3089),
.A2(n_214),
.B1(n_217),
.B2(n_218),
.Y(n_3387)
);

CKINVDCx5p33_ASAP7_75t_R g3388 ( 
.A(n_3123),
.Y(n_3388)
);

AO32x2_ASAP7_75t_L g3389 ( 
.A1(n_3180),
.A2(n_214),
.A3(n_218),
.B1(n_219),
.B2(n_221),
.Y(n_3389)
);

AOI21xp5_ASAP7_75t_L g3390 ( 
.A1(n_3149),
.A2(n_219),
.B(n_221),
.Y(n_3390)
);

AOI21xp5_ASAP7_75t_L g3391 ( 
.A1(n_3184),
.A2(n_222),
.B(n_223),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_3125),
.B(n_222),
.Y(n_3392)
);

AOI21xp5_ASAP7_75t_L g3393 ( 
.A1(n_3202),
.A2(n_223),
.B(n_224),
.Y(n_3393)
);

AOI21x1_ASAP7_75t_L g3394 ( 
.A1(n_3204),
.A2(n_225),
.B(n_227),
.Y(n_3394)
);

CKINVDCx5p33_ASAP7_75t_R g3395 ( 
.A(n_3130),
.Y(n_3395)
);

A2O1A1Ixp33_ASAP7_75t_L g3396 ( 
.A1(n_3253),
.A2(n_225),
.B(n_227),
.C(n_228),
.Y(n_3396)
);

O2A1O1Ixp33_ASAP7_75t_L g3397 ( 
.A1(n_3189),
.A2(n_229),
.B(n_231),
.C(n_232),
.Y(n_3397)
);

BUFx3_ASAP7_75t_L g3398 ( 
.A(n_3155),
.Y(n_3398)
);

AOI21xp5_ASAP7_75t_L g3399 ( 
.A1(n_3150),
.A2(n_229),
.B(n_231),
.Y(n_3399)
);

AOI221x1_ASAP7_75t_L g3400 ( 
.A1(n_3204),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.C(n_237),
.Y(n_3400)
);

OAI21x1_ASAP7_75t_L g3401 ( 
.A1(n_3131),
.A2(n_443),
.B(n_435),
.Y(n_3401)
);

AOI221xp5_ASAP7_75t_SL g3402 ( 
.A1(n_3167),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.C(n_238),
.Y(n_3402)
);

AOI31xp67_ASAP7_75t_L g3403 ( 
.A1(n_3211),
.A2(n_239),
.A3(n_240),
.B(n_241),
.Y(n_3403)
);

INVx2_ASAP7_75t_L g3404 ( 
.A(n_3146),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3168),
.Y(n_3405)
);

OAI21x1_ASAP7_75t_L g3406 ( 
.A1(n_3302),
.A2(n_3095),
.B(n_3107),
.Y(n_3406)
);

OAI221xp5_ASAP7_75t_L g3407 ( 
.A1(n_3303),
.A2(n_3211),
.B1(n_3205),
.B2(n_3226),
.C(n_3251),
.Y(n_3407)
);

CKINVDCx20_ASAP7_75t_R g3408 ( 
.A(n_3318),
.Y(n_3408)
);

INVx2_ASAP7_75t_L g3409 ( 
.A(n_3358),
.Y(n_3409)
);

OAI221xp5_ASAP7_75t_L g3410 ( 
.A1(n_3301),
.A2(n_3205),
.B1(n_3226),
.B2(n_3251),
.C(n_3244),
.Y(n_3410)
);

CKINVDCx16_ASAP7_75t_R g3411 ( 
.A(n_3331),
.Y(n_3411)
);

BUFx2_ASAP7_75t_R g3412 ( 
.A(n_3325),
.Y(n_3412)
);

OAI21x1_ASAP7_75t_L g3413 ( 
.A1(n_3312),
.A2(n_3102),
.B(n_3111),
.Y(n_3413)
);

OAI21x1_ASAP7_75t_SL g3414 ( 
.A1(n_3394),
.A2(n_3176),
.B(n_3129),
.Y(n_3414)
);

OAI21x1_ASAP7_75t_SL g3415 ( 
.A1(n_3365),
.A2(n_3129),
.B(n_3201),
.Y(n_3415)
);

AOI22xp33_ASAP7_75t_L g3416 ( 
.A1(n_3256),
.A2(n_3177),
.B1(n_3204),
.B2(n_3126),
.Y(n_3416)
);

INVx6_ASAP7_75t_L g3417 ( 
.A(n_3267),
.Y(n_3417)
);

OAI21x1_ASAP7_75t_L g3418 ( 
.A1(n_3291),
.A2(n_3118),
.B(n_3238),
.Y(n_3418)
);

AOI22xp33_ASAP7_75t_L g3419 ( 
.A1(n_3341),
.A2(n_3203),
.B1(n_3136),
.B2(n_3124),
.Y(n_3419)
);

OR2x6_ASAP7_75t_L g3420 ( 
.A(n_3336),
.B(n_3124),
.Y(n_3420)
);

AO21x2_ASAP7_75t_L g3421 ( 
.A1(n_3304),
.A2(n_3133),
.B(n_3160),
.Y(n_3421)
);

AOI21x1_ASAP7_75t_L g3422 ( 
.A1(n_3340),
.A2(n_3246),
.B(n_3160),
.Y(n_3422)
);

AO31x2_ASAP7_75t_L g3423 ( 
.A1(n_3400),
.A2(n_3098),
.A3(n_3106),
.B(n_3148),
.Y(n_3423)
);

AO21x2_ASAP7_75t_L g3424 ( 
.A1(n_3265),
.A2(n_3133),
.B(n_3213),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3405),
.B(n_3098),
.Y(n_3425)
);

OAI21xp5_ASAP7_75t_L g3426 ( 
.A1(n_3345),
.A2(n_3148),
.B(n_3116),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_3314),
.B(n_3106),
.Y(n_3427)
);

INVx4_ASAP7_75t_L g3428 ( 
.A(n_3297),
.Y(n_3428)
);

BUFx10_ASAP7_75t_L g3429 ( 
.A(n_3332),
.Y(n_3429)
);

CKINVDCx11_ASAP7_75t_R g3430 ( 
.A(n_3267),
.Y(n_3430)
);

AOI21xp5_ASAP7_75t_L g3431 ( 
.A1(n_3257),
.A2(n_3150),
.B(n_3239),
.Y(n_3431)
);

OAI21xp5_ASAP7_75t_L g3432 ( 
.A1(n_3399),
.A2(n_3152),
.B(n_3151),
.Y(n_3432)
);

OAI21xp5_ASAP7_75t_L g3433 ( 
.A1(n_3356),
.A2(n_3244),
.B(n_3216),
.Y(n_3433)
);

OR2x2_ASAP7_75t_L g3434 ( 
.A(n_3353),
.B(n_3230),
.Y(n_3434)
);

BUFx8_ASAP7_75t_L g3435 ( 
.A(n_3274),
.Y(n_3435)
);

HB1xp67_ASAP7_75t_L g3436 ( 
.A(n_3277),
.Y(n_3436)
);

NAND3xp33_ASAP7_75t_L g3437 ( 
.A(n_3308),
.B(n_3216),
.C(n_3232),
.Y(n_3437)
);

NAND3xp33_ASAP7_75t_L g3438 ( 
.A(n_3402),
.B(n_3232),
.C(n_3213),
.Y(n_3438)
);

INVxp67_ASAP7_75t_L g3439 ( 
.A(n_3342),
.Y(n_3439)
);

NOR2x1_ASAP7_75t_SL g3440 ( 
.A(n_3336),
.B(n_3236),
.Y(n_3440)
);

O2A1O1Ixp33_ASAP7_75t_L g3441 ( 
.A1(n_3328),
.A2(n_3329),
.B(n_3385),
.C(n_3296),
.Y(n_3441)
);

AOI22x1_ASAP7_75t_L g3442 ( 
.A1(n_3280),
.A2(n_3243),
.B1(n_3163),
.B2(n_3199),
.Y(n_3442)
);

CKINVDCx11_ASAP7_75t_R g3443 ( 
.A(n_3310),
.Y(n_3443)
);

AOI21x1_ASAP7_75t_L g3444 ( 
.A1(n_3382),
.A2(n_3215),
.B(n_3207),
.Y(n_3444)
);

OAI211xp5_ASAP7_75t_L g3445 ( 
.A1(n_3327),
.A2(n_3305),
.B(n_3321),
.C(n_3306),
.Y(n_3445)
);

CKINVDCx20_ASAP7_75t_R g3446 ( 
.A(n_3388),
.Y(n_3446)
);

OR2x6_ASAP7_75t_L g3447 ( 
.A(n_3383),
.B(n_3236),
.Y(n_3447)
);

BUFx6f_ASAP7_75t_L g3448 ( 
.A(n_3346),
.Y(n_3448)
);

AO21x2_ASAP7_75t_L g3449 ( 
.A1(n_3259),
.A2(n_3350),
.B(n_3362),
.Y(n_3449)
);

OAI21x1_ASAP7_75t_L g3450 ( 
.A1(n_3295),
.A2(n_3183),
.B(n_3175),
.Y(n_3450)
);

OAI21xp5_ASAP7_75t_L g3451 ( 
.A1(n_3279),
.A2(n_3215),
.B(n_3182),
.Y(n_3451)
);

NOR2xp33_ASAP7_75t_L g3452 ( 
.A(n_3271),
.B(n_3249),
.Y(n_3452)
);

INVx1_ASAP7_75t_SL g3453 ( 
.A(n_3344),
.Y(n_3453)
);

AO31x2_ASAP7_75t_L g3454 ( 
.A1(n_3334),
.A2(n_3230),
.A3(n_3138),
.B(n_3145),
.Y(n_3454)
);

OAI22xp5_ASAP7_75t_L g3455 ( 
.A1(n_3299),
.A2(n_3182),
.B1(n_3223),
.B2(n_3236),
.Y(n_3455)
);

AOI22xp33_ASAP7_75t_L g3456 ( 
.A1(n_3260),
.A2(n_3361),
.B1(n_3380),
.B2(n_3366),
.Y(n_3456)
);

OAI21x1_ASAP7_75t_L g3457 ( 
.A1(n_3359),
.A2(n_3181),
.B(n_3166),
.Y(n_3457)
);

OAI21xp5_ASAP7_75t_L g3458 ( 
.A1(n_3349),
.A2(n_3225),
.B(n_3249),
.Y(n_3458)
);

OAI21x1_ASAP7_75t_L g3459 ( 
.A1(n_3348),
.A2(n_3309),
.B(n_3263),
.Y(n_3459)
);

AO31x2_ASAP7_75t_L g3460 ( 
.A1(n_3396),
.A2(n_3210),
.A3(n_3179),
.B(n_3188),
.Y(n_3460)
);

AND2x2_ASAP7_75t_L g3461 ( 
.A(n_3289),
.B(n_3363),
.Y(n_3461)
);

INVx4_ASAP7_75t_SL g3462 ( 
.A(n_3337),
.Y(n_3462)
);

BUFx2_ASAP7_75t_SL g3463 ( 
.A(n_3398),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_SL g3464 ( 
.A(n_3379),
.B(n_3155),
.Y(n_3464)
);

AOI221xp5_ASAP7_75t_L g3465 ( 
.A1(n_3282),
.A2(n_239),
.B1(n_242),
.B2(n_243),
.C(n_244),
.Y(n_3465)
);

INVx2_ASAP7_75t_L g3466 ( 
.A(n_3375),
.Y(n_3466)
);

HB1xp67_ASAP7_75t_L g3467 ( 
.A(n_3272),
.Y(n_3467)
);

INVx2_ASAP7_75t_SL g3468 ( 
.A(n_3395),
.Y(n_3468)
);

A2O1A1Ixp33_ASAP7_75t_L g3469 ( 
.A1(n_3317),
.A2(n_3223),
.B(n_3210),
.C(n_246),
.Y(n_3469)
);

O2A1O1Ixp33_ASAP7_75t_L g3470 ( 
.A1(n_3355),
.A2(n_3245),
.B(n_243),
.C(n_246),
.Y(n_3470)
);

OA21x2_ASAP7_75t_L g3471 ( 
.A1(n_3392),
.A2(n_3171),
.B(n_3104),
.Y(n_3471)
);

BUFx6f_ASAP7_75t_L g3472 ( 
.A(n_3346),
.Y(n_3472)
);

NAND2x1p5_ASAP7_75t_L g3473 ( 
.A(n_3313),
.B(n_3223),
.Y(n_3473)
);

BUFx3_ASAP7_75t_L g3474 ( 
.A(n_3292),
.Y(n_3474)
);

INVx3_ASAP7_75t_L g3475 ( 
.A(n_3347),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3322),
.Y(n_3476)
);

NOR2xp33_ASAP7_75t_SL g3477 ( 
.A(n_3300),
.B(n_3245),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3404),
.Y(n_3478)
);

NAND2x1p5_ASAP7_75t_L g3479 ( 
.A(n_3347),
.B(n_3104),
.Y(n_3479)
);

NOR2xp33_ASAP7_75t_L g3480 ( 
.A(n_3357),
.B(n_3367),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3320),
.B(n_3188),
.Y(n_3481)
);

OAI21x1_ASAP7_75t_L g3482 ( 
.A1(n_3326),
.A2(n_3179),
.B(n_3188),
.Y(n_3482)
);

AND2x2_ASAP7_75t_L g3483 ( 
.A(n_3373),
.B(n_3245),
.Y(n_3483)
);

OAI221xp5_ASAP7_75t_L g3484 ( 
.A1(n_3306),
.A2(n_242),
.B1(n_248),
.B2(n_249),
.C(n_252),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3320),
.B(n_252),
.Y(n_3485)
);

NAND2x1p5_ASAP7_75t_L g3486 ( 
.A(n_3346),
.B(n_372),
.Y(n_3486)
);

AO31x2_ASAP7_75t_L g3487 ( 
.A1(n_3371),
.A2(n_254),
.A3(n_258),
.B(n_259),
.Y(n_3487)
);

AND2x4_ASAP7_75t_L g3488 ( 
.A(n_3377),
.B(n_259),
.Y(n_3488)
);

OR2x6_ASAP7_75t_L g3489 ( 
.A(n_3316),
.B(n_3319),
.Y(n_3489)
);

NOR2x1_ASAP7_75t_L g3490 ( 
.A(n_3376),
.B(n_261),
.Y(n_3490)
);

OAI21x1_ASAP7_75t_L g3491 ( 
.A1(n_3269),
.A2(n_261),
.B(n_262),
.Y(n_3491)
);

INVx8_ASAP7_75t_L g3492 ( 
.A(n_3374),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3376),
.B(n_265),
.Y(n_3493)
);

OAI21x1_ASAP7_75t_L g3494 ( 
.A1(n_3401),
.A2(n_267),
.B(n_268),
.Y(n_3494)
);

NOR4xp25_ASAP7_75t_L g3495 ( 
.A(n_3397),
.B(n_269),
.C(n_270),
.D(n_271),
.Y(n_3495)
);

OAI21x1_ASAP7_75t_L g3496 ( 
.A1(n_3268),
.A2(n_271),
.B(n_272),
.Y(n_3496)
);

NAND2x1p5_ASAP7_75t_L g3497 ( 
.A(n_3266),
.B(n_382),
.Y(n_3497)
);

INVx2_ASAP7_75t_SL g3498 ( 
.A(n_3286),
.Y(n_3498)
);

NAND3xp33_ASAP7_75t_L g3499 ( 
.A(n_3386),
.B(n_273),
.C(n_274),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3323),
.Y(n_3500)
);

AOI22xp33_ASAP7_75t_SL g3501 ( 
.A1(n_3361),
.A2(n_273),
.B1(n_275),
.B2(n_276),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3294),
.B(n_278),
.Y(n_3502)
);

OA21x2_ASAP7_75t_L g3503 ( 
.A1(n_3378),
.A2(n_279),
.B(n_280),
.Y(n_3503)
);

INVx1_ASAP7_75t_SL g3504 ( 
.A(n_3379),
.Y(n_3504)
);

OR2x2_ASAP7_75t_L g3505 ( 
.A(n_3311),
.B(n_3381),
.Y(n_3505)
);

OAI21x1_ASAP7_75t_L g3506 ( 
.A1(n_3293),
.A2(n_280),
.B(n_281),
.Y(n_3506)
);

BUFx6f_ASAP7_75t_SL g3507 ( 
.A(n_3310),
.Y(n_3507)
);

OAI21xp5_ASAP7_75t_L g3508 ( 
.A1(n_3351),
.A2(n_282),
.B(n_283),
.Y(n_3508)
);

OAI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_3352),
.A2(n_3354),
.B(n_3369),
.Y(n_3509)
);

INVx2_ASAP7_75t_L g3510 ( 
.A(n_3337),
.Y(n_3510)
);

AND2x4_ASAP7_75t_L g3511 ( 
.A(n_3384),
.B(n_283),
.Y(n_3511)
);

AOI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_3324),
.A2(n_393),
.B(n_428),
.Y(n_3512)
);

OA21x2_ASAP7_75t_L g3513 ( 
.A1(n_3418),
.A2(n_3298),
.B(n_3288),
.Y(n_3513)
);

AOI21xp5_ASAP7_75t_L g3514 ( 
.A1(n_3509),
.A2(n_3368),
.B(n_3266),
.Y(n_3514)
);

NAND4xp25_ASAP7_75t_L g3515 ( 
.A(n_3456),
.B(n_3290),
.C(n_3321),
.D(n_3299),
.Y(n_3515)
);

OAI22xp5_ASAP7_75t_L g3516 ( 
.A1(n_3416),
.A2(n_3330),
.B1(n_3360),
.B2(n_3339),
.Y(n_3516)
);

AOI21x1_ASAP7_75t_L g3517 ( 
.A1(n_3485),
.A2(n_3384),
.B(n_3258),
.Y(n_3517)
);

INVx2_ASAP7_75t_SL g3518 ( 
.A(n_3428),
.Y(n_3518)
);

CKINVDCx5p33_ASAP7_75t_R g3519 ( 
.A(n_3408),
.Y(n_3519)
);

INVx3_ASAP7_75t_L g3520 ( 
.A(n_3448),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_3504),
.Y(n_3521)
);

A2O1A1Ixp33_ASAP7_75t_L g3522 ( 
.A1(n_3441),
.A2(n_3333),
.B(n_3273),
.C(n_3372),
.Y(n_3522)
);

OR2x6_ASAP7_75t_L g3523 ( 
.A(n_3463),
.B(n_3403),
.Y(n_3523)
);

OAI21x1_ASAP7_75t_L g3524 ( 
.A1(n_3479),
.A2(n_3281),
.B(n_3270),
.Y(n_3524)
);

INVx2_ASAP7_75t_L g3525 ( 
.A(n_3504),
.Y(n_3525)
);

AOI21x1_ASAP7_75t_L g3526 ( 
.A1(n_3485),
.A2(n_3284),
.B(n_3387),
.Y(n_3526)
);

AOI21x1_ASAP7_75t_L g3527 ( 
.A1(n_3493),
.A2(n_3284),
.B(n_3390),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3425),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3425),
.Y(n_3529)
);

OA21x2_ASAP7_75t_L g3530 ( 
.A1(n_3481),
.A2(n_3264),
.B(n_3275),
.Y(n_3530)
);

AO21x2_ASAP7_75t_L g3531 ( 
.A1(n_3493),
.A2(n_3393),
.B(n_3283),
.Y(n_3531)
);

INVx3_ASAP7_75t_L g3532 ( 
.A(n_3448),
.Y(n_3532)
);

INVx1_ASAP7_75t_SL g3533 ( 
.A(n_3412),
.Y(n_3533)
);

CKINVDCx11_ASAP7_75t_R g3534 ( 
.A(n_3446),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3427),
.Y(n_3535)
);

OAI21x1_ASAP7_75t_L g3536 ( 
.A1(n_3479),
.A2(n_3278),
.B(n_3338),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3439),
.B(n_3364),
.Y(n_3537)
);

INVxp67_ASAP7_75t_L g3538 ( 
.A(n_3490),
.Y(n_3538)
);

CKINVDCx20_ASAP7_75t_R g3539 ( 
.A(n_3411),
.Y(n_3539)
);

AO21x2_ASAP7_75t_L g3540 ( 
.A1(n_3481),
.A2(n_3391),
.B(n_3343),
.Y(n_3540)
);

NOR2xp33_ASAP7_75t_L g3541 ( 
.A(n_3429),
.B(n_3370),
.Y(n_3541)
);

AO31x2_ASAP7_75t_L g3542 ( 
.A1(n_3510),
.A2(n_3261),
.A3(n_3389),
.B(n_3276),
.Y(n_3542)
);

NAND3xp33_ASAP7_75t_L g3543 ( 
.A(n_3509),
.B(n_3262),
.C(n_3287),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3500),
.Y(n_3544)
);

A2O1A1Ixp33_ASAP7_75t_L g3545 ( 
.A1(n_3470),
.A2(n_3445),
.B(n_3508),
.C(n_3501),
.Y(n_3545)
);

OAI21x1_ASAP7_75t_SL g3546 ( 
.A1(n_3440),
.A2(n_3276),
.B(n_3389),
.Y(n_3546)
);

BUFx6f_ASAP7_75t_L g3547 ( 
.A(n_3448),
.Y(n_3547)
);

A2O1A1Ixp33_ASAP7_75t_L g3548 ( 
.A1(n_3508),
.A2(n_3389),
.B(n_3276),
.C(n_3315),
.Y(n_3548)
);

OAI21x1_ASAP7_75t_L g3549 ( 
.A1(n_3413),
.A2(n_3337),
.B(n_3285),
.Y(n_3549)
);

AOI21x1_ASAP7_75t_L g3550 ( 
.A1(n_3464),
.A2(n_3335),
.B(n_3315),
.Y(n_3550)
);

HB1xp67_ASAP7_75t_L g3551 ( 
.A(n_3462),
.Y(n_3551)
);

OA21x2_ASAP7_75t_L g3552 ( 
.A1(n_3459),
.A2(n_3335),
.B(n_3315),
.Y(n_3552)
);

AO221x2_ASAP7_75t_L g3553 ( 
.A1(n_3433),
.A2(n_3432),
.B1(n_3426),
.B2(n_3451),
.C(n_3437),
.Y(n_3553)
);

OAI21xp5_ASAP7_75t_L g3554 ( 
.A1(n_3499),
.A2(n_3307),
.B(n_3335),
.Y(n_3554)
);

INVx2_ASAP7_75t_L g3555 ( 
.A(n_3466),
.Y(n_3555)
);

HB1xp67_ASAP7_75t_L g3556 ( 
.A(n_3462),
.Y(n_3556)
);

BUFx8_ASAP7_75t_SL g3557 ( 
.A(n_3507),
.Y(n_3557)
);

OR2x6_ASAP7_75t_L g3558 ( 
.A(n_3447),
.B(n_3285),
.Y(n_3558)
);

OAI21x1_ASAP7_75t_L g3559 ( 
.A1(n_3422),
.A2(n_3473),
.B(n_3406),
.Y(n_3559)
);

AOI21xp5_ASAP7_75t_L g3560 ( 
.A1(n_3469),
.A2(n_284),
.B(n_285),
.Y(n_3560)
);

AND2x2_ASAP7_75t_L g3561 ( 
.A(n_3453),
.B(n_287),
.Y(n_3561)
);

OA21x2_ASAP7_75t_L g3562 ( 
.A1(n_3432),
.A2(n_287),
.B(n_290),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3467),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3476),
.Y(n_3564)
);

OA21x2_ASAP7_75t_L g3565 ( 
.A1(n_3451),
.A2(n_290),
.B(n_291),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3461),
.B(n_293),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3478),
.Y(n_3567)
);

AO21x2_ASAP7_75t_L g3568 ( 
.A1(n_3414),
.A2(n_295),
.B(n_296),
.Y(n_3568)
);

BUFx3_ASAP7_75t_L g3569 ( 
.A(n_3428),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3434),
.Y(n_3570)
);

INVx2_ASAP7_75t_L g3571 ( 
.A(n_3462),
.Y(n_3571)
);

OAI21x1_ASAP7_75t_SL g3572 ( 
.A1(n_3415),
.A2(n_295),
.B(n_296),
.Y(n_3572)
);

AOI21xp5_ASAP7_75t_L g3573 ( 
.A1(n_3489),
.A2(n_298),
.B(n_299),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3436),
.Y(n_3574)
);

AO31x2_ASAP7_75t_L g3575 ( 
.A1(n_3455),
.A2(n_298),
.A3(n_300),
.B(n_301),
.Y(n_3575)
);

OAI21x1_ASAP7_75t_SL g3576 ( 
.A1(n_3444),
.A2(n_302),
.B(n_304),
.Y(n_3576)
);

AOI21xp5_ASAP7_75t_L g3577 ( 
.A1(n_3489),
.A2(n_302),
.B(n_373),
.Y(n_3577)
);

AOI21xp5_ASAP7_75t_L g3578 ( 
.A1(n_3489),
.A2(n_375),
.B(n_377),
.Y(n_3578)
);

NOR2x1_ASAP7_75t_SL g3579 ( 
.A(n_3420),
.B(n_380),
.Y(n_3579)
);

OR2x2_ASAP7_75t_L g3580 ( 
.A(n_3505),
.B(n_385),
.Y(n_3580)
);

AOI22xp33_ASAP7_75t_SL g3581 ( 
.A1(n_3410),
.A2(n_3484),
.B1(n_3407),
.B2(n_3433),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3409),
.Y(n_3582)
);

AO21x2_ASAP7_75t_L g3583 ( 
.A1(n_3431),
.A2(n_388),
.B(n_395),
.Y(n_3583)
);

CKINVDCx5p33_ASAP7_75t_R g3584 ( 
.A(n_3430),
.Y(n_3584)
);

INVx2_ASAP7_75t_L g3585 ( 
.A(n_3503),
.Y(n_3585)
);

NOR2xp33_ASAP7_75t_L g3586 ( 
.A(n_3429),
.B(n_397),
.Y(n_3586)
);

OA21x2_ASAP7_75t_L g3587 ( 
.A1(n_3426),
.A2(n_398),
.B(n_404),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_3503),
.Y(n_3588)
);

CKINVDCx11_ASAP7_75t_R g3589 ( 
.A(n_3443),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3480),
.B(n_3423),
.Y(n_3590)
);

AOI21x1_ASAP7_75t_L g3591 ( 
.A1(n_3511),
.A2(n_407),
.B(n_409),
.Y(n_3591)
);

INVx2_ASAP7_75t_L g3592 ( 
.A(n_3475),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3423),
.B(n_411),
.Y(n_3593)
);

BUFx3_ASAP7_75t_L g3594 ( 
.A(n_3498),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_3423),
.B(n_413),
.Y(n_3595)
);

OA21x2_ASAP7_75t_L g3596 ( 
.A1(n_3482),
.A2(n_414),
.B(n_415),
.Y(n_3596)
);

AND2x2_ASAP7_75t_L g3597 ( 
.A(n_3474),
.B(n_417),
.Y(n_3597)
);

INVx2_ASAP7_75t_L g3598 ( 
.A(n_3471),
.Y(n_3598)
);

OAI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3495),
.A2(n_425),
.B(n_426),
.Y(n_3599)
);

HB1xp67_ASAP7_75t_L g3600 ( 
.A(n_3471),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3483),
.Y(n_3601)
);

BUFx2_ASAP7_75t_L g3602 ( 
.A(n_3472),
.Y(n_3602)
);

BUFx2_ASAP7_75t_L g3603 ( 
.A(n_3472),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3472),
.Y(n_3604)
);

AOI21xp5_ASAP7_75t_L g3605 ( 
.A1(n_3449),
.A2(n_433),
.B(n_3465),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_3473),
.Y(n_3606)
);

AO31x2_ASAP7_75t_L g3607 ( 
.A1(n_3455),
.A2(n_3452),
.A3(n_3512),
.B(n_3460),
.Y(n_3607)
);

AOI22xp33_ASAP7_75t_L g3608 ( 
.A1(n_3484),
.A2(n_3465),
.B1(n_3410),
.B2(n_3438),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3460),
.Y(n_3609)
);

CKINVDCx14_ASAP7_75t_R g3610 ( 
.A(n_3589),
.Y(n_3610)
);

BUFx2_ASAP7_75t_SL g3611 ( 
.A(n_3539),
.Y(n_3611)
);

BUFx12f_ASAP7_75t_L g3612 ( 
.A(n_3589),
.Y(n_3612)
);

OAI21xp33_ASAP7_75t_L g3613 ( 
.A1(n_3581),
.A2(n_3419),
.B(n_3438),
.Y(n_3613)
);

OAI22xp5_ASAP7_75t_SL g3614 ( 
.A1(n_3539),
.A2(n_3412),
.B1(n_3447),
.B2(n_3468),
.Y(n_3614)
);

AOI22xp33_ASAP7_75t_L g3615 ( 
.A1(n_3553),
.A2(n_3424),
.B1(n_3458),
.B2(n_3442),
.Y(n_3615)
);

INVx6_ASAP7_75t_L g3616 ( 
.A(n_3569),
.Y(n_3616)
);

AOI22xp5_ASAP7_75t_L g3617 ( 
.A1(n_3553),
.A2(n_3424),
.B1(n_3477),
.B2(n_3458),
.Y(n_3617)
);

OAI21xp33_ASAP7_75t_L g3618 ( 
.A1(n_3608),
.A2(n_3497),
.B(n_3511),
.Y(n_3618)
);

INVx3_ASAP7_75t_L g3619 ( 
.A(n_3557),
.Y(n_3619)
);

AOI22xp33_ASAP7_75t_L g3620 ( 
.A1(n_3553),
.A2(n_3507),
.B1(n_3492),
.B2(n_3435),
.Y(n_3620)
);

AND2x4_ASAP7_75t_SL g3621 ( 
.A(n_3558),
.B(n_3488),
.Y(n_3621)
);

NOR2xp33_ASAP7_75t_L g3622 ( 
.A(n_3569),
.B(n_3435),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_3585),
.B(n_3454),
.Y(n_3623)
);

AOI22xp33_ASAP7_75t_SL g3624 ( 
.A1(n_3516),
.A2(n_3477),
.B1(n_3502),
.B2(n_3492),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_3547),
.Y(n_3625)
);

BUFx12f_ASAP7_75t_L g3626 ( 
.A(n_3534),
.Y(n_3626)
);

OAI21xp5_ASAP7_75t_SL g3627 ( 
.A1(n_3608),
.A2(n_3486),
.B(n_3487),
.Y(n_3627)
);

AOI22xp33_ASAP7_75t_SL g3628 ( 
.A1(n_3546),
.A2(n_3494),
.B1(n_3491),
.B2(n_3496),
.Y(n_3628)
);

AOI22xp33_ASAP7_75t_L g3629 ( 
.A1(n_3605),
.A2(n_3599),
.B1(n_3514),
.B2(n_3560),
.Y(n_3629)
);

AOI22xp33_ASAP7_75t_L g3630 ( 
.A1(n_3562),
.A2(n_3417),
.B1(n_3421),
.B2(n_3506),
.Y(n_3630)
);

OAI21xp5_ASAP7_75t_SL g3631 ( 
.A1(n_3545),
.A2(n_3522),
.B(n_3538),
.Y(n_3631)
);

OAI22xp5_ASAP7_75t_L g3632 ( 
.A1(n_3545),
.A2(n_3487),
.B1(n_3454),
.B2(n_3460),
.Y(n_3632)
);

CKINVDCx5p33_ASAP7_75t_R g3633 ( 
.A(n_3534),
.Y(n_3633)
);

NAND3xp33_ASAP7_75t_L g3634 ( 
.A(n_3554),
.B(n_3487),
.C(n_3457),
.Y(n_3634)
);

CKINVDCx20_ASAP7_75t_R g3635 ( 
.A(n_3519),
.Y(n_3635)
);

OAI22xp33_ASAP7_75t_SL g3636 ( 
.A1(n_3538),
.A2(n_3450),
.B1(n_3590),
.B2(n_3585),
.Y(n_3636)
);

AOI22xp33_ASAP7_75t_L g3637 ( 
.A1(n_3587),
.A2(n_3565),
.B1(n_3531),
.B2(n_3543),
.Y(n_3637)
);

AOI22xp33_ASAP7_75t_L g3638 ( 
.A1(n_3587),
.A2(n_3565),
.B1(n_3531),
.B2(n_3568),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3570),
.Y(n_3639)
);

OAI21xp5_ASAP7_75t_SL g3640 ( 
.A1(n_3522),
.A2(n_3548),
.B(n_3573),
.Y(n_3640)
);

OAI21xp33_ASAP7_75t_L g3641 ( 
.A1(n_3548),
.A2(n_3595),
.B(n_3593),
.Y(n_3641)
);

INVx2_ASAP7_75t_SL g3642 ( 
.A(n_3594),
.Y(n_3642)
);

BUFx6f_ASAP7_75t_L g3643 ( 
.A(n_3557),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3588),
.B(n_3528),
.Y(n_3644)
);

NOR2xp33_ASAP7_75t_L g3645 ( 
.A(n_3518),
.B(n_3533),
.Y(n_3645)
);

INVx4_ASAP7_75t_L g3646 ( 
.A(n_3594),
.Y(n_3646)
);

HB1xp67_ASAP7_75t_L g3647 ( 
.A(n_3588),
.Y(n_3647)
);

OAI22xp33_ASAP7_75t_L g3648 ( 
.A1(n_3523),
.A2(n_3558),
.B1(n_3526),
.B2(n_3577),
.Y(n_3648)
);

OAI22xp33_ASAP7_75t_L g3649 ( 
.A1(n_3523),
.A2(n_3521),
.B1(n_3525),
.B2(n_3574),
.Y(n_3649)
);

AOI22xp33_ASAP7_75t_L g3650 ( 
.A1(n_3583),
.A2(n_3540),
.B1(n_3513),
.B2(n_3572),
.Y(n_3650)
);

AOI22xp33_ASAP7_75t_L g3651 ( 
.A1(n_3513),
.A2(n_3601),
.B1(n_3578),
.B2(n_3576),
.Y(n_3651)
);

OAI22xp5_ASAP7_75t_L g3652 ( 
.A1(n_3604),
.A2(n_3541),
.B1(n_3537),
.B2(n_3521),
.Y(n_3652)
);

OAI21xp5_ASAP7_75t_L g3653 ( 
.A1(n_3550),
.A2(n_3527),
.B(n_3524),
.Y(n_3653)
);

CKINVDCx20_ASAP7_75t_R g3654 ( 
.A(n_3597),
.Y(n_3654)
);

BUFx3_ASAP7_75t_L g3655 ( 
.A(n_3561),
.Y(n_3655)
);

OAI22xp5_ASAP7_75t_L g3656 ( 
.A1(n_3520),
.A2(n_3532),
.B1(n_3566),
.B2(n_3580),
.Y(n_3656)
);

OAI21xp33_ASAP7_75t_L g3657 ( 
.A1(n_3609),
.A2(n_3586),
.B(n_3535),
.Y(n_3657)
);

OAI21xp5_ASAP7_75t_SL g3658 ( 
.A1(n_3586),
.A2(n_3517),
.B(n_3551),
.Y(n_3658)
);

OAI21xp5_ASAP7_75t_SL g3659 ( 
.A1(n_3551),
.A2(n_3556),
.B(n_3591),
.Y(n_3659)
);

OAI21xp5_ASAP7_75t_SL g3660 ( 
.A1(n_3571),
.A2(n_3600),
.B(n_3606),
.Y(n_3660)
);

AOI22xp33_ASAP7_75t_L g3661 ( 
.A1(n_3529),
.A2(n_3552),
.B1(n_3563),
.B2(n_3596),
.Y(n_3661)
);

INVx4_ASAP7_75t_L g3662 ( 
.A(n_3596),
.Y(n_3662)
);

OAI21xp5_ASAP7_75t_SL g3663 ( 
.A1(n_3600),
.A2(n_3607),
.B(n_3575),
.Y(n_3663)
);

AOI22xp33_ASAP7_75t_L g3664 ( 
.A1(n_3530),
.A2(n_3567),
.B1(n_3564),
.B2(n_3536),
.Y(n_3664)
);

AOI22xp33_ASAP7_75t_SL g3665 ( 
.A1(n_3579),
.A2(n_3575),
.B1(n_3549),
.B2(n_3530),
.Y(n_3665)
);

OAI21xp5_ASAP7_75t_L g3666 ( 
.A1(n_3559),
.A2(n_3555),
.B(n_3582),
.Y(n_3666)
);

HB1xp67_ASAP7_75t_L g3667 ( 
.A(n_3544),
.Y(n_3667)
);

AOI22xp33_ASAP7_75t_SL g3668 ( 
.A1(n_3575),
.A2(n_3598),
.B1(n_3607),
.B2(n_3542),
.Y(n_3668)
);

INVx3_ASAP7_75t_L g3669 ( 
.A(n_3592),
.Y(n_3669)
);

OAI21xp5_ASAP7_75t_SL g3670 ( 
.A1(n_3542),
.A2(n_3581),
.B(n_3608),
.Y(n_3670)
);

OAI22xp5_ASAP7_75t_L g3671 ( 
.A1(n_3542),
.A2(n_3581),
.B1(n_3545),
.B2(n_3608),
.Y(n_3671)
);

AOI22xp33_ASAP7_75t_L g3672 ( 
.A1(n_3542),
.A2(n_3553),
.B1(n_3581),
.B2(n_3515),
.Y(n_3672)
);

NAND2xp33_ASAP7_75t_R g3673 ( 
.A(n_3584),
.B(n_1301),
.Y(n_3673)
);

OAI22xp5_ASAP7_75t_L g3674 ( 
.A1(n_3581),
.A2(n_3545),
.B1(n_3608),
.B2(n_3456),
.Y(n_3674)
);

OAI22xp5_ASAP7_75t_L g3675 ( 
.A1(n_3581),
.A2(n_3545),
.B1(n_3608),
.B2(n_3456),
.Y(n_3675)
);

NOR2xp33_ASAP7_75t_L g3676 ( 
.A(n_3569),
.B(n_3584),
.Y(n_3676)
);

AND2x2_ASAP7_75t_L g3677 ( 
.A(n_3602),
.B(n_3603),
.Y(n_3677)
);

OAI22xp5_ASAP7_75t_L g3678 ( 
.A1(n_3581),
.A2(n_3545),
.B1(n_3608),
.B2(n_3456),
.Y(n_3678)
);

AOI22xp33_ASAP7_75t_L g3679 ( 
.A1(n_3553),
.A2(n_3581),
.B1(n_3515),
.B2(n_3608),
.Y(n_3679)
);

AOI22xp33_ASAP7_75t_SL g3680 ( 
.A1(n_3553),
.A2(n_3516),
.B1(n_3445),
.B2(n_3546),
.Y(n_3680)
);

NAND2x1p5_ASAP7_75t_L g3681 ( 
.A(n_3565),
.B(n_3504),
.Y(n_3681)
);

AOI22xp33_ASAP7_75t_L g3682 ( 
.A1(n_3553),
.A2(n_3581),
.B1(n_3515),
.B2(n_3608),
.Y(n_3682)
);

AOI22xp33_ASAP7_75t_L g3683 ( 
.A1(n_3553),
.A2(n_3581),
.B1(n_3515),
.B2(n_3608),
.Y(n_3683)
);

INVx3_ASAP7_75t_L g3684 ( 
.A(n_3557),
.Y(n_3684)
);

OAI21xp33_ASAP7_75t_L g3685 ( 
.A1(n_3581),
.A2(n_3608),
.B(n_3545),
.Y(n_3685)
);

NOR2xp33_ASAP7_75t_L g3686 ( 
.A(n_3569),
.B(n_3584),
.Y(n_3686)
);

OAI21xp33_ASAP7_75t_L g3687 ( 
.A1(n_3581),
.A2(n_3608),
.B(n_3545),
.Y(n_3687)
);

AOI222xp33_ASAP7_75t_L g3688 ( 
.A1(n_3608),
.A2(n_3545),
.B1(n_3516),
.B2(n_3456),
.C1(n_3509),
.C2(n_3538),
.Y(n_3688)
);

AOI222xp33_ASAP7_75t_L g3689 ( 
.A1(n_3608),
.A2(n_3545),
.B1(n_3516),
.B2(n_3456),
.C1(n_3509),
.C2(n_3538),
.Y(n_3689)
);

AND2x2_ASAP7_75t_L g3690 ( 
.A(n_3677),
.B(n_3625),
.Y(n_3690)
);

INVxp67_ASAP7_75t_SL g3691 ( 
.A(n_3681),
.Y(n_3691)
);

AO21x2_ASAP7_75t_L g3692 ( 
.A1(n_3663),
.A2(n_3648),
.B(n_3653),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3647),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3647),
.Y(n_3694)
);

AO21x2_ASAP7_75t_L g3695 ( 
.A1(n_3648),
.A2(n_3670),
.B(n_3649),
.Y(n_3695)
);

AO21x2_ASAP7_75t_L g3696 ( 
.A1(n_3671),
.A2(n_3658),
.B(n_3623),
.Y(n_3696)
);

INVx2_ASAP7_75t_L g3697 ( 
.A(n_3646),
.Y(n_3697)
);

AND2x4_ASAP7_75t_L g3698 ( 
.A(n_3662),
.B(n_3646),
.Y(n_3698)
);

OAI21xp5_ASAP7_75t_L g3699 ( 
.A1(n_3685),
.A2(n_3687),
.B(n_3674),
.Y(n_3699)
);

INVx6_ASAP7_75t_L g3700 ( 
.A(n_3612),
.Y(n_3700)
);

OA21x2_ASAP7_75t_L g3701 ( 
.A1(n_3672),
.A2(n_3640),
.B(n_3683),
.Y(n_3701)
);

OR2x6_ASAP7_75t_L g3702 ( 
.A(n_3611),
.B(n_3627),
.Y(n_3702)
);

AND2x4_ASAP7_75t_L g3703 ( 
.A(n_3662),
.B(n_3669),
.Y(n_3703)
);

INVxp67_ASAP7_75t_SL g3704 ( 
.A(n_3642),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3680),
.B(n_3613),
.Y(n_3705)
);

OA21x2_ASAP7_75t_L g3706 ( 
.A1(n_3679),
.A2(n_3682),
.B(n_3650),
.Y(n_3706)
);

OAI21xp33_ASAP7_75t_L g3707 ( 
.A1(n_3680),
.A2(n_3675),
.B(n_3678),
.Y(n_3707)
);

OR2x2_ASAP7_75t_L g3708 ( 
.A(n_3644),
.B(n_3639),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_3616),
.Y(n_3709)
);

CKINVDCx20_ASAP7_75t_R g3710 ( 
.A(n_3635),
.Y(n_3710)
);

INVx2_ASAP7_75t_L g3711 ( 
.A(n_3616),
.Y(n_3711)
);

BUFx2_ASAP7_75t_L g3712 ( 
.A(n_3619),
.Y(n_3712)
);

HB1xp67_ASAP7_75t_L g3713 ( 
.A(n_3667),
.Y(n_3713)
);

AND2x2_ASAP7_75t_L g3714 ( 
.A(n_3620),
.B(n_3624),
.Y(n_3714)
);

OA21x2_ASAP7_75t_L g3715 ( 
.A1(n_3634),
.A2(n_3641),
.B(n_3637),
.Y(n_3715)
);

OR2x6_ASAP7_75t_L g3716 ( 
.A(n_3616),
.B(n_3614),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3667),
.Y(n_3717)
);

BUFx3_ASAP7_75t_L g3718 ( 
.A(n_3643),
.Y(n_3718)
);

INVx3_ASAP7_75t_L g3719 ( 
.A(n_3619),
.Y(n_3719)
);

INVx3_ASAP7_75t_L g3720 ( 
.A(n_3684),
.Y(n_3720)
);

INVx2_ASAP7_75t_SL g3721 ( 
.A(n_3643),
.Y(n_3721)
);

INVx2_ASAP7_75t_L g3722 ( 
.A(n_3655),
.Y(n_3722)
);

INVx3_ASAP7_75t_L g3723 ( 
.A(n_3684),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_L g3724 ( 
.A(n_3688),
.B(n_3689),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3618),
.B(n_3629),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3668),
.Y(n_3726)
);

INVx2_ASAP7_75t_SL g3727 ( 
.A(n_3643),
.Y(n_3727)
);

BUFx2_ASAP7_75t_L g3728 ( 
.A(n_3610),
.Y(n_3728)
);

INVx2_ASAP7_75t_L g3729 ( 
.A(n_3621),
.Y(n_3729)
);

HB1xp67_ASAP7_75t_L g3730 ( 
.A(n_3632),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3628),
.B(n_3615),
.Y(n_3731)
);

INVx2_ASAP7_75t_L g3732 ( 
.A(n_3626),
.Y(n_3732)
);

HB1xp67_ASAP7_75t_L g3733 ( 
.A(n_3652),
.Y(n_3733)
);

AO21x2_ASAP7_75t_L g3734 ( 
.A1(n_3666),
.A2(n_3617),
.B(n_3660),
.Y(n_3734)
);

HB1xp67_ASAP7_75t_L g3735 ( 
.A(n_3645),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3668),
.Y(n_3736)
);

HB1xp67_ASAP7_75t_L g3737 ( 
.A(n_3656),
.Y(n_3737)
);

OR2x2_ASAP7_75t_L g3738 ( 
.A(n_3638),
.B(n_3661),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3633),
.Y(n_3739)
);

AO21x2_ASAP7_75t_L g3740 ( 
.A1(n_3659),
.A2(n_3657),
.B(n_3636),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3628),
.Y(n_3741)
);

INVx3_ASAP7_75t_L g3742 ( 
.A(n_3665),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3665),
.Y(n_3743)
);

INVx2_ASAP7_75t_L g3744 ( 
.A(n_3654),
.Y(n_3744)
);

INVx3_ASAP7_75t_L g3745 ( 
.A(n_3622),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3676),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3664),
.Y(n_3747)
);

HB1xp67_ASAP7_75t_L g3748 ( 
.A(n_3630),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3686),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3651),
.Y(n_3750)
);

AND2x2_ASAP7_75t_L g3751 ( 
.A(n_3673),
.B(n_3677),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3647),
.Y(n_3752)
);

INVx3_ASAP7_75t_SL g3753 ( 
.A(n_3643),
.Y(n_3753)
);

INVxp67_ASAP7_75t_SL g3754 ( 
.A(n_3681),
.Y(n_3754)
);

HB1xp67_ASAP7_75t_L g3755 ( 
.A(n_3647),
.Y(n_3755)
);

AO21x2_ASAP7_75t_L g3756 ( 
.A1(n_3663),
.A2(n_3648),
.B(n_3653),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3647),
.Y(n_3757)
);

AND2x2_ASAP7_75t_L g3758 ( 
.A(n_3677),
.B(n_3625),
.Y(n_3758)
);

AND2x2_ASAP7_75t_L g3759 ( 
.A(n_3677),
.B(n_3625),
.Y(n_3759)
);

INVx3_ASAP7_75t_L g3760 ( 
.A(n_3646),
.Y(n_3760)
);

AND2x2_ASAP7_75t_L g3761 ( 
.A(n_3677),
.B(n_3625),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3647),
.Y(n_3762)
);

AND2x2_ASAP7_75t_L g3763 ( 
.A(n_3677),
.B(n_3625),
.Y(n_3763)
);

OR2x6_ASAP7_75t_L g3764 ( 
.A(n_3631),
.B(n_3640),
.Y(n_3764)
);

HB1xp67_ASAP7_75t_L g3765 ( 
.A(n_3647),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3647),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3713),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3755),
.Y(n_3768)
);

AND2x2_ASAP7_75t_L g3769 ( 
.A(n_3712),
.B(n_3716),
.Y(n_3769)
);

AND2x4_ASAP7_75t_L g3770 ( 
.A(n_3712),
.B(n_3719),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_3716),
.B(n_3728),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3765),
.Y(n_3772)
);

AO21x2_ASAP7_75t_L g3773 ( 
.A1(n_3726),
.A2(n_3736),
.B(n_3695),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3742),
.B(n_3735),
.Y(n_3774)
);

HB1xp67_ASAP7_75t_L g3775 ( 
.A(n_3693),
.Y(n_3775)
);

INVx3_ASAP7_75t_L g3776 ( 
.A(n_3700),
.Y(n_3776)
);

AND2x4_ASAP7_75t_L g3777 ( 
.A(n_3719),
.B(n_3720),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3694),
.Y(n_3778)
);

INVx4_ASAP7_75t_L g3779 ( 
.A(n_3753),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3742),
.B(n_3733),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3742),
.Y(n_3781)
);

INVx1_ASAP7_75t_L g3782 ( 
.A(n_3752),
.Y(n_3782)
);

BUFx2_ASAP7_75t_L g3783 ( 
.A(n_3728),
.Y(n_3783)
);

INVx5_ASAP7_75t_L g3784 ( 
.A(n_3700),
.Y(n_3784)
);

BUFx3_ASAP7_75t_L g3785 ( 
.A(n_3718),
.Y(n_3785)
);

INVx2_ASAP7_75t_L g3786 ( 
.A(n_3698),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3752),
.Y(n_3787)
);

OR2x2_ASAP7_75t_L g3788 ( 
.A(n_3726),
.B(n_3736),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3757),
.Y(n_3789)
);

OR2x2_ASAP7_75t_L g3790 ( 
.A(n_3708),
.B(n_3757),
.Y(n_3790)
);

BUFx3_ASAP7_75t_L g3791 ( 
.A(n_3718),
.Y(n_3791)
);

AND2x2_ASAP7_75t_L g3792 ( 
.A(n_3716),
.B(n_3719),
.Y(n_3792)
);

INVx2_ASAP7_75t_L g3793 ( 
.A(n_3698),
.Y(n_3793)
);

BUFx6f_ASAP7_75t_L g3794 ( 
.A(n_3753),
.Y(n_3794)
);

OA21x2_ASAP7_75t_L g3795 ( 
.A1(n_3743),
.A2(n_3705),
.B(n_3731),
.Y(n_3795)
);

INVx2_ASAP7_75t_SL g3796 ( 
.A(n_3700),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3762),
.Y(n_3797)
);

BUFx3_ASAP7_75t_L g3798 ( 
.A(n_3718),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_3701),
.B(n_3743),
.Y(n_3799)
);

INVx2_ASAP7_75t_L g3800 ( 
.A(n_3698),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3716),
.B(n_3720),
.Y(n_3801)
);

INVx2_ASAP7_75t_SL g3802 ( 
.A(n_3700),
.Y(n_3802)
);

AOI22xp33_ASAP7_75t_L g3803 ( 
.A1(n_3764),
.A2(n_3707),
.B1(n_3724),
.B2(n_3701),
.Y(n_3803)
);

INVx2_ASAP7_75t_L g3804 ( 
.A(n_3698),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_3703),
.Y(n_3805)
);

INVx2_ASAP7_75t_L g3806 ( 
.A(n_3703),
.Y(n_3806)
);

AND2x2_ASAP7_75t_L g3807 ( 
.A(n_3716),
.B(n_3720),
.Y(n_3807)
);

BUFx3_ASAP7_75t_L g3808 ( 
.A(n_3753),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3703),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3766),
.Y(n_3810)
);

HB1xp67_ASAP7_75t_L g3811 ( 
.A(n_3766),
.Y(n_3811)
);

INVx1_ASAP7_75t_SL g3812 ( 
.A(n_3751),
.Y(n_3812)
);

AND2x4_ASAP7_75t_L g3813 ( 
.A(n_3723),
.B(n_3760),
.Y(n_3813)
);

INVx3_ASAP7_75t_L g3814 ( 
.A(n_3703),
.Y(n_3814)
);

INVx2_ASAP7_75t_L g3815 ( 
.A(n_3721),
.Y(n_3815)
);

HB1xp67_ASAP7_75t_L g3816 ( 
.A(n_3717),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_3701),
.B(n_3751),
.Y(n_3817)
);

AND2x2_ASAP7_75t_L g3818 ( 
.A(n_3723),
.B(n_3690),
.Y(n_3818)
);

OAI22xp5_ASAP7_75t_L g3819 ( 
.A1(n_3702),
.A2(n_3764),
.B1(n_3741),
.B2(n_3730),
.Y(n_3819)
);

INVx2_ASAP7_75t_L g3820 ( 
.A(n_3721),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_3701),
.B(n_3737),
.Y(n_3821)
);

AND2x2_ASAP7_75t_L g3822 ( 
.A(n_3723),
.B(n_3690),
.Y(n_3822)
);

AND2x2_ASAP7_75t_L g3823 ( 
.A(n_3758),
.B(n_3759),
.Y(n_3823)
);

INVxp67_ASAP7_75t_L g3824 ( 
.A(n_3727),
.Y(n_3824)
);

INVx2_ASAP7_75t_L g3825 ( 
.A(n_3727),
.Y(n_3825)
);

AND2x2_ASAP7_75t_L g3826 ( 
.A(n_3758),
.B(n_3759),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3760),
.Y(n_3827)
);

AND2x2_ASAP7_75t_L g3828 ( 
.A(n_3761),
.B(n_3763),
.Y(n_3828)
);

HB1xp67_ASAP7_75t_L g3829 ( 
.A(n_3722),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3722),
.B(n_3750),
.Y(n_3830)
);

AND2x4_ASAP7_75t_L g3831 ( 
.A(n_3760),
.B(n_3729),
.Y(n_3831)
);

INVxp67_ASAP7_75t_SL g3832 ( 
.A(n_3744),
.Y(n_3832)
);

AOI222xp33_ASAP7_75t_L g3833 ( 
.A1(n_3707),
.A2(n_3699),
.B1(n_3725),
.B2(n_3741),
.C1(n_3750),
.C2(n_3748),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_L g3834 ( 
.A(n_3706),
.B(n_3704),
.Y(n_3834)
);

AO31x2_ASAP7_75t_L g3835 ( 
.A1(n_3747),
.A2(n_3711),
.A3(n_3709),
.B(n_3697),
.Y(n_3835)
);

AND2x2_ASAP7_75t_L g3836 ( 
.A(n_3761),
.B(n_3763),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3744),
.Y(n_3837)
);

INVx2_ASAP7_75t_L g3838 ( 
.A(n_3764),
.Y(n_3838)
);

INVx2_ASAP7_75t_L g3839 ( 
.A(n_3764),
.Y(n_3839)
);

AND2x2_ASAP7_75t_L g3840 ( 
.A(n_3783),
.B(n_3695),
.Y(n_3840)
);

INVx2_ASAP7_75t_L g3841 ( 
.A(n_3773),
.Y(n_3841)
);

AND2x2_ASAP7_75t_L g3842 ( 
.A(n_3783),
.B(n_3695),
.Y(n_3842)
);

INVx2_ASAP7_75t_L g3843 ( 
.A(n_3773),
.Y(n_3843)
);

AND2x2_ASAP7_75t_L g3844 ( 
.A(n_3771),
.B(n_3756),
.Y(n_3844)
);

AND2x2_ASAP7_75t_L g3845 ( 
.A(n_3771),
.B(n_3756),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3773),
.Y(n_3846)
);

INVx2_ASAP7_75t_L g3847 ( 
.A(n_3770),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3816),
.Y(n_3848)
);

AND2x2_ASAP7_75t_L g3849 ( 
.A(n_3769),
.B(n_3756),
.Y(n_3849)
);

AND2x2_ASAP7_75t_L g3850 ( 
.A(n_3769),
.B(n_3692),
.Y(n_3850)
);

HB1xp67_ASAP7_75t_L g3851 ( 
.A(n_3812),
.Y(n_3851)
);

OR2x2_ASAP7_75t_L g3852 ( 
.A(n_3795),
.B(n_3715),
.Y(n_3852)
);

INVx2_ASAP7_75t_L g3853 ( 
.A(n_3770),
.Y(n_3853)
);

AND2x2_ASAP7_75t_L g3854 ( 
.A(n_3818),
.B(n_3692),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3775),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_3795),
.B(n_3706),
.Y(n_3856)
);

OR2x2_ASAP7_75t_L g3857 ( 
.A(n_3795),
.B(n_3715),
.Y(n_3857)
);

INVx3_ASAP7_75t_L g3858 ( 
.A(n_3770),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3811),
.Y(n_3859)
);

OR2x2_ASAP7_75t_L g3860 ( 
.A(n_3795),
.B(n_3715),
.Y(n_3860)
);

AND2x4_ASAP7_75t_L g3861 ( 
.A(n_3777),
.B(n_3692),
.Y(n_3861)
);

AND2x2_ASAP7_75t_L g3862 ( 
.A(n_3818),
.B(n_3764),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3833),
.B(n_3706),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3790),
.Y(n_3864)
);

BUFx2_ASAP7_75t_L g3865 ( 
.A(n_3777),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3790),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3767),
.Y(n_3867)
);

BUFx3_ASAP7_75t_L g3868 ( 
.A(n_3794),
.Y(n_3868)
);

AND2x4_ASAP7_75t_L g3869 ( 
.A(n_3777),
.B(n_3691),
.Y(n_3869)
);

AND2x2_ASAP7_75t_L g3870 ( 
.A(n_3822),
.B(n_3740),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3767),
.Y(n_3871)
);

AND2x2_ASAP7_75t_L g3872 ( 
.A(n_3822),
.B(n_3740),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3794),
.Y(n_3873)
);

AND2x2_ASAP7_75t_L g3874 ( 
.A(n_3823),
.B(n_3740),
.Y(n_3874)
);

AND2x2_ASAP7_75t_L g3875 ( 
.A(n_3823),
.B(n_3734),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3768),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3768),
.Y(n_3877)
);

INVx2_ASAP7_75t_L g3878 ( 
.A(n_3794),
.Y(n_3878)
);

OR2x2_ASAP7_75t_L g3879 ( 
.A(n_3799),
.B(n_3715),
.Y(n_3879)
);

INVx2_ASAP7_75t_L g3880 ( 
.A(n_3794),
.Y(n_3880)
);

AND2x2_ASAP7_75t_L g3881 ( 
.A(n_3826),
.B(n_3734),
.Y(n_3881)
);

NOR2xp33_ASAP7_75t_L g3882 ( 
.A(n_3779),
.B(n_3732),
.Y(n_3882)
);

BUFx6f_ASAP7_75t_L g3883 ( 
.A(n_3794),
.Y(n_3883)
);

AND2x4_ASAP7_75t_L g3884 ( 
.A(n_3785),
.B(n_3754),
.Y(n_3884)
);

AND2x2_ASAP7_75t_L g3885 ( 
.A(n_3826),
.B(n_3734),
.Y(n_3885)
);

AND2x2_ASAP7_75t_L g3886 ( 
.A(n_3828),
.B(n_3702),
.Y(n_3886)
);

BUFx2_ASAP7_75t_L g3887 ( 
.A(n_3781),
.Y(n_3887)
);

AND2x2_ASAP7_75t_L g3888 ( 
.A(n_3828),
.B(n_3702),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3772),
.Y(n_3889)
);

AND2x2_ASAP7_75t_L g3890 ( 
.A(n_3836),
.B(n_3702),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_L g3891 ( 
.A(n_3781),
.B(n_3706),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_3803),
.B(n_3738),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3832),
.B(n_3738),
.Y(n_3893)
);

NOR2xp33_ASAP7_75t_L g3894 ( 
.A(n_3863),
.B(n_3779),
.Y(n_3894)
);

OA21x2_ASAP7_75t_L g3895 ( 
.A1(n_3841),
.A2(n_3821),
.B(n_3834),
.Y(n_3895)
);

AND2x2_ASAP7_75t_L g3896 ( 
.A(n_3858),
.B(n_3776),
.Y(n_3896)
);

INVx2_ASAP7_75t_L g3897 ( 
.A(n_3852),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3852),
.B(n_3837),
.Y(n_3898)
);

NOR2xp33_ASAP7_75t_L g3899 ( 
.A(n_3863),
.B(n_3779),
.Y(n_3899)
);

INVx2_ASAP7_75t_L g3900 ( 
.A(n_3852),
.Y(n_3900)
);

OR2x2_ASAP7_75t_L g3901 ( 
.A(n_3857),
.B(n_3788),
.Y(n_3901)
);

INVxp67_ASAP7_75t_SL g3902 ( 
.A(n_3857),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_SL g3903 ( 
.A(n_3857),
.B(n_3860),
.Y(n_3903)
);

AND2x2_ASAP7_75t_L g3904 ( 
.A(n_3858),
.B(n_3776),
.Y(n_3904)
);

OR2x2_ASAP7_75t_L g3905 ( 
.A(n_3860),
.B(n_3788),
.Y(n_3905)
);

BUFx3_ASAP7_75t_L g3906 ( 
.A(n_3841),
.Y(n_3906)
);

NOR2xp67_ASAP7_75t_L g3907 ( 
.A(n_3860),
.B(n_3784),
.Y(n_3907)
);

INVx2_ASAP7_75t_L g3908 ( 
.A(n_3841),
.Y(n_3908)
);

NAND3xp33_ASAP7_75t_L g3909 ( 
.A(n_3856),
.B(n_3817),
.C(n_3780),
.Y(n_3909)
);

INVx2_ASAP7_75t_L g3910 ( 
.A(n_3841),
.Y(n_3910)
);

INVxp67_ASAP7_75t_SL g3911 ( 
.A(n_3843),
.Y(n_3911)
);

NAND2xp5_ASAP7_75t_L g3912 ( 
.A(n_3856),
.B(n_3837),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3843),
.Y(n_3913)
);

BUFx3_ASAP7_75t_L g3914 ( 
.A(n_3843),
.Y(n_3914)
);

AOI22xp33_ASAP7_75t_L g3915 ( 
.A1(n_3892),
.A2(n_3702),
.B1(n_3696),
.B2(n_3747),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3843),
.Y(n_3916)
);

INVxp67_ASAP7_75t_L g3917 ( 
.A(n_3865),
.Y(n_3917)
);

AND2x2_ASAP7_75t_L g3918 ( 
.A(n_3858),
.B(n_3776),
.Y(n_3918)
);

HB1xp67_ASAP7_75t_L g3919 ( 
.A(n_3846),
.Y(n_3919)
);

AOI22xp33_ASAP7_75t_L g3920 ( 
.A1(n_3892),
.A2(n_3696),
.B1(n_3714),
.B2(n_3819),
.Y(n_3920)
);

AND2x4_ASAP7_75t_L g3921 ( 
.A(n_3858),
.B(n_3785),
.Y(n_3921)
);

AND2x2_ASAP7_75t_L g3922 ( 
.A(n_3858),
.B(n_3836),
.Y(n_3922)
);

INVx2_ASAP7_75t_L g3923 ( 
.A(n_3846),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3846),
.Y(n_3924)
);

AND2x2_ASAP7_75t_L g3925 ( 
.A(n_3865),
.B(n_3808),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3879),
.B(n_3772),
.Y(n_3926)
);

AND2x2_ASAP7_75t_L g3927 ( 
.A(n_3865),
.B(n_3808),
.Y(n_3927)
);

AND2x2_ASAP7_75t_L g3928 ( 
.A(n_3840),
.B(n_3792),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3879),
.B(n_3887),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3879),
.B(n_3829),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3846),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3840),
.B(n_3792),
.Y(n_3932)
);

INVx2_ASAP7_75t_L g3933 ( 
.A(n_3840),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3842),
.Y(n_3934)
);

AND2x2_ASAP7_75t_L g3935 ( 
.A(n_3842),
.B(n_3801),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3887),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3842),
.Y(n_3937)
);

AND2x2_ASAP7_75t_L g3938 ( 
.A(n_3847),
.B(n_3801),
.Y(n_3938)
);

HB1xp67_ASAP7_75t_L g3939 ( 
.A(n_3887),
.Y(n_3939)
);

BUFx2_ASAP7_75t_SL g3940 ( 
.A(n_3868),
.Y(n_3940)
);

OA211x2_ASAP7_75t_L g3941 ( 
.A1(n_3882),
.A2(n_3824),
.B(n_3774),
.C(n_3830),
.Y(n_3941)
);

INVx3_ASAP7_75t_L g3942 ( 
.A(n_3861),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3851),
.Y(n_3943)
);

AND2x2_ASAP7_75t_L g3944 ( 
.A(n_3847),
.B(n_3807),
.Y(n_3944)
);

AND2x2_ASAP7_75t_L g3945 ( 
.A(n_3847),
.B(n_3807),
.Y(n_3945)
);

AND2x2_ASAP7_75t_L g3946 ( 
.A(n_3928),
.B(n_3932),
.Y(n_3946)
);

AND2x2_ASAP7_75t_L g3947 ( 
.A(n_3928),
.B(n_3796),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3897),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3902),
.B(n_3851),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3939),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3939),
.Y(n_3951)
);

AND2x2_ASAP7_75t_L g3952 ( 
.A(n_3928),
.B(n_3796),
.Y(n_3952)
);

AND2x2_ASAP7_75t_L g3953 ( 
.A(n_3932),
.B(n_3802),
.Y(n_3953)
);

HB1xp67_ASAP7_75t_L g3954 ( 
.A(n_3903),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3902),
.B(n_3864),
.Y(n_3955)
);

INVx2_ASAP7_75t_SL g3956 ( 
.A(n_3903),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3897),
.Y(n_3957)
);

AOI221xp5_ASAP7_75t_L g3958 ( 
.A1(n_3920),
.A2(n_3893),
.B1(n_3891),
.B2(n_3855),
.C(n_3859),
.Y(n_3958)
);

BUFx2_ASAP7_75t_SL g3959 ( 
.A(n_3907),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3897),
.Y(n_3960)
);

AND2x2_ASAP7_75t_L g3961 ( 
.A(n_3932),
.B(n_3802),
.Y(n_3961)
);

INVx2_ASAP7_75t_L g3962 ( 
.A(n_3897),
.Y(n_3962)
);

AND2x2_ASAP7_75t_L g3963 ( 
.A(n_3935),
.B(n_3791),
.Y(n_3963)
);

INVx2_ASAP7_75t_L g3964 ( 
.A(n_3900),
.Y(n_3964)
);

OR2x2_ASAP7_75t_L g3965 ( 
.A(n_3900),
.B(n_3893),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3917),
.B(n_3864),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3900),
.Y(n_3967)
);

BUFx2_ASAP7_75t_L g3968 ( 
.A(n_3900),
.Y(n_3968)
);

INVxp67_ASAP7_75t_SL g3969 ( 
.A(n_3901),
.Y(n_3969)
);

INVx2_ASAP7_75t_L g3970 ( 
.A(n_3901),
.Y(n_3970)
);

AND2x2_ASAP7_75t_L g3971 ( 
.A(n_3935),
.B(n_3791),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_L g3972 ( 
.A(n_3917),
.B(n_3866),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3935),
.B(n_3798),
.Y(n_3973)
);

INVx2_ASAP7_75t_L g3974 ( 
.A(n_3901),
.Y(n_3974)
);

INVx2_ASAP7_75t_L g3975 ( 
.A(n_3905),
.Y(n_3975)
);

AND2x2_ASAP7_75t_L g3976 ( 
.A(n_3922),
.B(n_3798),
.Y(n_3976)
);

OAI33xp33_ASAP7_75t_L g3977 ( 
.A1(n_3909),
.A2(n_3905),
.A3(n_3926),
.B1(n_3929),
.B2(n_3912),
.B3(n_3898),
.Y(n_3977)
);

AND2x2_ASAP7_75t_L g3978 ( 
.A(n_3922),
.B(n_3847),
.Y(n_3978)
);

AND2x2_ASAP7_75t_L g3979 ( 
.A(n_3922),
.B(n_3925),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3925),
.B(n_3853),
.Y(n_3980)
);

HB1xp67_ASAP7_75t_L g3981 ( 
.A(n_3905),
.Y(n_3981)
);

AND2x2_ASAP7_75t_L g3982 ( 
.A(n_3925),
.B(n_3853),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3936),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3936),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3968),
.Y(n_3985)
);

INVx2_ASAP7_75t_SL g3986 ( 
.A(n_3979),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_3979),
.B(n_3927),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3968),
.Y(n_3988)
);

INVx1_ASAP7_75t_L g3989 ( 
.A(n_3968),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_L g3990 ( 
.A(n_3979),
.B(n_3927),
.Y(n_3990)
);

HB1xp67_ASAP7_75t_L g3991 ( 
.A(n_3954),
.Y(n_3991)
);

AND2x2_ASAP7_75t_L g3992 ( 
.A(n_3946),
.B(n_3862),
.Y(n_3992)
);

AND2x4_ASAP7_75t_SL g3993 ( 
.A(n_3976),
.B(n_3921),
.Y(n_3993)
);

INVx2_ASAP7_75t_L g3994 ( 
.A(n_3956),
.Y(n_3994)
);

AND2x2_ASAP7_75t_L g3995 ( 
.A(n_3946),
.B(n_3862),
.Y(n_3995)
);

AND2x2_ASAP7_75t_L g3996 ( 
.A(n_3946),
.B(n_3862),
.Y(n_3996)
);

INVx2_ASAP7_75t_L g3997 ( 
.A(n_3956),
.Y(n_3997)
);

NOR2x1p5_ASAP7_75t_L g3998 ( 
.A(n_3949),
.B(n_3943),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3954),
.Y(n_3999)
);

OA211x2_ASAP7_75t_L g4000 ( 
.A1(n_3958),
.A2(n_3882),
.B(n_3899),
.C(n_3894),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_3963),
.B(n_3927),
.Y(n_4001)
);

AND2x2_ASAP7_75t_L g4002 ( 
.A(n_3963),
.B(n_3784),
.Y(n_4002)
);

AND2x2_ASAP7_75t_L g4003 ( 
.A(n_3963),
.B(n_3784),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_L g4004 ( 
.A(n_3971),
.B(n_3938),
.Y(n_4004)
);

INVx2_ASAP7_75t_L g4005 ( 
.A(n_3956),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3981),
.Y(n_4006)
);

INVx2_ASAP7_75t_L g4007 ( 
.A(n_3981),
.Y(n_4007)
);

INVx2_ASAP7_75t_L g4008 ( 
.A(n_3970),
.Y(n_4008)
);

AND2x2_ASAP7_75t_L g4009 ( 
.A(n_3971),
.B(n_3784),
.Y(n_4009)
);

NOR2xp33_ASAP7_75t_L g4010 ( 
.A(n_3971),
.B(n_3784),
.Y(n_4010)
);

AND2x2_ASAP7_75t_L g4011 ( 
.A(n_3992),
.B(n_3745),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_L g4012 ( 
.A(n_4007),
.B(n_3969),
.Y(n_4012)
);

OR2x2_ASAP7_75t_L g4013 ( 
.A(n_4001),
.B(n_3987),
.Y(n_4013)
);

AND2x2_ASAP7_75t_L g4014 ( 
.A(n_3992),
.B(n_3745),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_L g4015 ( 
.A(n_4007),
.B(n_3969),
.Y(n_4015)
);

OR2x2_ASAP7_75t_L g4016 ( 
.A(n_3990),
.B(n_3949),
.Y(n_4016)
);

AND2x2_ASAP7_75t_L g4017 ( 
.A(n_3995),
.B(n_3996),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_L g4018 ( 
.A(n_3986),
.B(n_3970),
.Y(n_4018)
);

AND2x2_ASAP7_75t_L g4019 ( 
.A(n_3995),
.B(n_3745),
.Y(n_4019)
);

AND2x2_ASAP7_75t_L g4020 ( 
.A(n_3996),
.B(n_3973),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_3986),
.B(n_3970),
.Y(n_4021)
);

HB1xp67_ASAP7_75t_L g4022 ( 
.A(n_3985),
.Y(n_4022)
);

INVx2_ASAP7_75t_SL g4023 ( 
.A(n_3993),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3993),
.B(n_3973),
.Y(n_4024)
);

AND2x4_ASAP7_75t_L g4025 ( 
.A(n_3993),
.B(n_3980),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_L g4026 ( 
.A(n_4006),
.B(n_3974),
.Y(n_4026)
);

INVx2_ASAP7_75t_L g4027 ( 
.A(n_3985),
.Y(n_4027)
);

AND2x2_ASAP7_75t_L g4028 ( 
.A(n_4002),
.B(n_3973),
.Y(n_4028)
);

AND2x2_ASAP7_75t_L g4029 ( 
.A(n_4002),
.B(n_3976),
.Y(n_4029)
);

NAND2x1_ASAP7_75t_L g4030 ( 
.A(n_4003),
.B(n_3921),
.Y(n_4030)
);

INVxp67_ASAP7_75t_SL g4031 ( 
.A(n_4022),
.Y(n_4031)
);

HB1xp67_ASAP7_75t_L g4032 ( 
.A(n_4025),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_4020),
.B(n_3976),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_4025),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_4018),
.Y(n_4035)
);

NAND2x1_ASAP7_75t_L g4036 ( 
.A(n_4023),
.B(n_3921),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_4018),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_4021),
.Y(n_4038)
);

INVx2_ASAP7_75t_L g4039 ( 
.A(n_4030),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_4021),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_4017),
.B(n_3947),
.Y(n_4041)
);

INVx2_ASAP7_75t_L g4042 ( 
.A(n_4028),
.Y(n_4042)
);

INVx2_ASAP7_75t_L g4043 ( 
.A(n_4011),
.Y(n_4043)
);

AND2x2_ASAP7_75t_L g4044 ( 
.A(n_4014),
.B(n_4019),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_L g4045 ( 
.A(n_4029),
.B(n_3947),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_4012),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_4024),
.B(n_3947),
.Y(n_4047)
);

NOR2xp67_ASAP7_75t_SL g4048 ( 
.A(n_4032),
.B(n_3991),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_SL g4049 ( 
.A(n_4033),
.B(n_3884),
.Y(n_4049)
);

NOR2xp67_ASAP7_75t_L g4050 ( 
.A(n_4032),
.B(n_3943),
.Y(n_4050)
);

AOI22xp33_ASAP7_75t_L g4051 ( 
.A1(n_4042),
.A2(n_3696),
.B1(n_4000),
.B2(n_3920),
.Y(n_4051)
);

NOR2xp67_ASAP7_75t_SL g4052 ( 
.A(n_4043),
.B(n_4016),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_4031),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_L g4054 ( 
.A(n_4034),
.B(n_3952),
.Y(n_4054)
);

INVx2_ASAP7_75t_SL g4055 ( 
.A(n_4036),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_4031),
.Y(n_4056)
);

INVx1_ASAP7_75t_SL g4057 ( 
.A(n_4041),
.Y(n_4057)
);

NOR2x1_ASAP7_75t_L g4058 ( 
.A(n_4039),
.B(n_4006),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_4039),
.B(n_3952),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_4055),
.B(n_3980),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_4048),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_4050),
.Y(n_4062)
);

AOI32xp33_ASAP7_75t_L g4063 ( 
.A1(n_4051),
.A2(n_3915),
.A3(n_3958),
.B1(n_3899),
.B2(n_3894),
.Y(n_4063)
);

AND2x2_ASAP7_75t_L g4064 ( 
.A(n_4054),
.B(n_3952),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_4059),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_R g4066 ( 
.A(n_4052),
.B(n_4044),
.Y(n_4066)
);

AOI22xp33_ASAP7_75t_SL g4067 ( 
.A1(n_4057),
.A2(n_3844),
.B1(n_3845),
.B2(n_3849),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_4060),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_4067),
.B(n_3980),
.Y(n_4069)
);

NAND3xp33_ASAP7_75t_L g4070 ( 
.A(n_4063),
.B(n_3999),
.C(n_3997),
.Y(n_4070)
);

OAI21xp5_ASAP7_75t_SL g4071 ( 
.A1(n_4064),
.A2(n_4004),
.B(n_4045),
.Y(n_4071)
);

AOI222xp33_ASAP7_75t_L g4072 ( 
.A1(n_4061),
.A2(n_3915),
.B1(n_3977),
.B2(n_3909),
.C1(n_3999),
.C2(n_3844),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_4062),
.B(n_3982),
.Y(n_4073)
);

AOI221xp5_ASAP7_75t_L g4074 ( 
.A1(n_4065),
.A2(n_3977),
.B1(n_4005),
.B2(n_3997),
.C(n_3994),
.Y(n_4074)
);

AOI22xp5_ASAP7_75t_L g4075 ( 
.A1(n_4066),
.A2(n_3961),
.B1(n_3953),
.B2(n_4000),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_4060),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_L g4077 ( 
.A(n_4067),
.B(n_3982),
.Y(n_4077)
);

AOI222xp33_ASAP7_75t_L g4078 ( 
.A1(n_4061),
.A2(n_3844),
.B1(n_3845),
.B2(n_3850),
.C1(n_3849),
.C2(n_3891),
.Y(n_4078)
);

AOI221xp5_ASAP7_75t_L g4079 ( 
.A1(n_4063),
.A2(n_4005),
.B1(n_3994),
.B2(n_4010),
.C(n_3926),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_4060),
.Y(n_4080)
);

AOI21xp33_ASAP7_75t_L g4081 ( 
.A1(n_4072),
.A2(n_4015),
.B(n_4012),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_4078),
.B(n_4003),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_4075),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_4073),
.Y(n_4084)
);

INVx1_ASAP7_75t_L g4085 ( 
.A(n_4069),
.Y(n_4085)
);

INVx1_ASAP7_75t_SL g4086 ( 
.A(n_4077),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_4070),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_4068),
.Y(n_4088)
);

AOI21xp5_ASAP7_75t_L g4089 ( 
.A1(n_4071),
.A2(n_4015),
.B(n_4026),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_4076),
.Y(n_4090)
);

INVx2_ASAP7_75t_L g4091 ( 
.A(n_4080),
.Y(n_4091)
);

INVx2_ASAP7_75t_L g4092 ( 
.A(n_4079),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_4074),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_4078),
.B(n_4009),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_4078),
.B(n_4009),
.Y(n_4095)
);

NAND2xp33_ASAP7_75t_SL g4096 ( 
.A(n_4073),
.B(n_3883),
.Y(n_4096)
);

AOI22xp5_ASAP7_75t_L g4097 ( 
.A1(n_4075),
.A2(n_3953),
.B1(n_3961),
.B2(n_3921),
.Y(n_4097)
);

O2A1O1Ixp33_ASAP7_75t_L g4098 ( 
.A1(n_4072),
.A2(n_3988),
.B(n_3989),
.C(n_4026),
.Y(n_4098)
);

O2A1O1Ixp33_ASAP7_75t_SL g4099 ( 
.A1(n_4069),
.A2(n_3988),
.B(n_3989),
.C(n_3951),
.Y(n_4099)
);

INVxp67_ASAP7_75t_L g4100 ( 
.A(n_4073),
.Y(n_4100)
);

INVx2_ASAP7_75t_L g4101 ( 
.A(n_4073),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_4075),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_4097),
.Y(n_4103)
);

AOI22xp5_ASAP7_75t_L g4104 ( 
.A1(n_4083),
.A2(n_3953),
.B1(n_3961),
.B2(n_3921),
.Y(n_4104)
);

AOI22xp5_ASAP7_75t_L g4105 ( 
.A1(n_4102),
.A2(n_3978),
.B1(n_3982),
.B2(n_4047),
.Y(n_4105)
);

OAI221xp5_ASAP7_75t_L g4106 ( 
.A1(n_4081),
.A2(n_3955),
.B1(n_3868),
.B2(n_3966),
.C(n_3972),
.Y(n_4106)
);

AOI32xp33_ASAP7_75t_L g4107 ( 
.A1(n_4086),
.A2(n_3868),
.A3(n_4058),
.B1(n_3951),
.B2(n_3950),
.Y(n_4107)
);

AOI22xp33_ASAP7_75t_L g4108 ( 
.A1(n_4093),
.A2(n_3941),
.B1(n_3868),
.B2(n_3883),
.Y(n_4108)
);

OAI21xp5_ASAP7_75t_SL g4109 ( 
.A1(n_4086),
.A2(n_4013),
.B(n_3972),
.Y(n_4109)
);

OAI221xp5_ASAP7_75t_SL g4110 ( 
.A1(n_4087),
.A2(n_3965),
.B1(n_3966),
.B2(n_3955),
.C(n_3878),
.Y(n_4110)
);

OR2x2_ASAP7_75t_L g4111 ( 
.A(n_4082),
.B(n_3940),
.Y(n_4111)
);

OAI31xp33_ASAP7_75t_L g4112 ( 
.A1(n_4096),
.A2(n_3998),
.A3(n_3950),
.B(n_4053),
.Y(n_4112)
);

AOI221xp5_ASAP7_75t_L g4113 ( 
.A1(n_4081),
.A2(n_3940),
.B1(n_3880),
.B2(n_3878),
.C(n_3873),
.Y(n_4113)
);

O2A1O1Ixp33_ASAP7_75t_L g4114 ( 
.A1(n_4099),
.A2(n_4027),
.B(n_4056),
.C(n_4008),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_4098),
.Y(n_4115)
);

AOI211xp5_ASAP7_75t_L g4116 ( 
.A1(n_4089),
.A2(n_4049),
.B(n_4008),
.C(n_4046),
.Y(n_4116)
);

AOI21xp33_ASAP7_75t_L g4117 ( 
.A1(n_4094),
.A2(n_4037),
.B(n_4035),
.Y(n_4117)
);

INVx2_ASAP7_75t_L g4118 ( 
.A(n_4101),
.Y(n_4118)
);

OAI21xp5_ASAP7_75t_L g4119 ( 
.A1(n_4100),
.A2(n_4043),
.B(n_3878),
.Y(n_4119)
);

NOR2xp33_ASAP7_75t_L g4120 ( 
.A(n_4095),
.B(n_4038),
.Y(n_4120)
);

AOI21xp33_ASAP7_75t_L g4121 ( 
.A1(n_4085),
.A2(n_4040),
.B(n_3965),
.Y(n_4121)
);

NOR2xp33_ASAP7_75t_L g4122 ( 
.A(n_4092),
.B(n_3732),
.Y(n_4122)
);

AOI22xp5_ASAP7_75t_L g4123 ( 
.A1(n_4088),
.A2(n_3978),
.B1(n_3896),
.B2(n_3918),
.Y(n_4123)
);

OAI22xp5_ASAP7_75t_L g4124 ( 
.A1(n_4084),
.A2(n_3815),
.B1(n_3820),
.B2(n_3825),
.Y(n_4124)
);

OAI22xp5_ASAP7_75t_L g4125 ( 
.A1(n_4090),
.A2(n_3815),
.B1(n_3820),
.B2(n_3825),
.Y(n_4125)
);

AOI22xp33_ASAP7_75t_L g4126 ( 
.A1(n_4091),
.A2(n_3941),
.B1(n_3883),
.B2(n_3938),
.Y(n_4126)
);

NOR2xp33_ASAP7_75t_L g4127 ( 
.A(n_4097),
.B(n_3873),
.Y(n_4127)
);

AOI221xp5_ASAP7_75t_L g4128 ( 
.A1(n_4081),
.A2(n_3940),
.B1(n_3880),
.B2(n_3878),
.C(n_3873),
.Y(n_4128)
);

NOR2xp33_ASAP7_75t_L g4129 ( 
.A(n_4104),
.B(n_4106),
.Y(n_4129)
);

OAI221xp5_ASAP7_75t_L g4130 ( 
.A1(n_4126),
.A2(n_3959),
.B1(n_3965),
.B2(n_3880),
.C(n_3873),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_4123),
.Y(n_4131)
);

AOI21xp5_ASAP7_75t_L g4132 ( 
.A1(n_4114),
.A2(n_4112),
.B(n_4109),
.Y(n_4132)
);

O2A1O1Ixp33_ASAP7_75t_L g4133 ( 
.A1(n_4110),
.A2(n_3998),
.B(n_3984),
.C(n_3983),
.Y(n_4133)
);

AO21x1_ASAP7_75t_L g4134 ( 
.A1(n_4116),
.A2(n_3960),
.B(n_3957),
.Y(n_4134)
);

OAI21xp33_ASAP7_75t_L g4135 ( 
.A1(n_4122),
.A2(n_3978),
.B(n_3880),
.Y(n_4135)
);

AOI21xp33_ASAP7_75t_SL g4136 ( 
.A1(n_4107),
.A2(n_3984),
.B(n_3983),
.Y(n_4136)
);

NAND4xp25_ASAP7_75t_SL g4137 ( 
.A(n_4108),
.B(n_3975),
.C(n_3974),
.D(n_3960),
.Y(n_4137)
);

AOI21xp5_ASAP7_75t_L g4138 ( 
.A1(n_4121),
.A2(n_3962),
.B(n_3948),
.Y(n_4138)
);

AOI221xp5_ASAP7_75t_SL g4139 ( 
.A1(n_4125),
.A2(n_3957),
.B1(n_3959),
.B2(n_3967),
.C(n_3964),
.Y(n_4139)
);

AOI21xp5_ASAP7_75t_L g4140 ( 
.A1(n_4119),
.A2(n_3962),
.B(n_3948),
.Y(n_4140)
);

NOR2xp33_ASAP7_75t_L g4141 ( 
.A(n_4105),
.B(n_3883),
.Y(n_4141)
);

AOI221xp5_ASAP7_75t_L g4142 ( 
.A1(n_4124),
.A2(n_3883),
.B1(n_3975),
.B2(n_3974),
.C(n_3964),
.Y(n_4142)
);

AOI211xp5_ASAP7_75t_L g4143 ( 
.A1(n_4117),
.A2(n_3883),
.B(n_3967),
.C(n_3964),
.Y(n_4143)
);

OAI211xp5_ASAP7_75t_SL g4144 ( 
.A1(n_4103),
.A2(n_3912),
.B(n_3930),
.C(n_3929),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_4111),
.Y(n_4145)
);

NOR2xp33_ASAP7_75t_L g4146 ( 
.A(n_4127),
.B(n_3883),
.Y(n_4146)
);

AOI22xp5_ASAP7_75t_L g4147 ( 
.A1(n_4120),
.A2(n_3883),
.B1(n_3904),
.B2(n_3896),
.Y(n_4147)
);

AOI22xp5_ASAP7_75t_L g4148 ( 
.A1(n_4118),
.A2(n_3918),
.B1(n_3904),
.B2(n_3896),
.Y(n_4148)
);

O2A1O1Ixp33_ASAP7_75t_L g4149 ( 
.A1(n_4115),
.A2(n_3975),
.B(n_3967),
.C(n_3962),
.Y(n_4149)
);

OAI221xp5_ASAP7_75t_L g4150 ( 
.A1(n_4113),
.A2(n_3930),
.B1(n_3907),
.B2(n_3948),
.C(n_3898),
.Y(n_4150)
);

AOI221xp5_ASAP7_75t_L g4151 ( 
.A1(n_4128),
.A2(n_3911),
.B1(n_3918),
.B2(n_3904),
.C(n_3867),
.Y(n_4151)
);

NAND3xp33_ASAP7_75t_L g4152 ( 
.A(n_4107),
.B(n_3919),
.C(n_3859),
.Y(n_4152)
);

AOI211xp5_ASAP7_75t_L g4153 ( 
.A1(n_4130),
.A2(n_3855),
.B(n_3911),
.C(n_3877),
.Y(n_4153)
);

AOI211xp5_ASAP7_75t_SL g4154 ( 
.A1(n_4132),
.A2(n_3945),
.B(n_3944),
.C(n_3938),
.Y(n_4154)
);

OAI211xp5_ASAP7_75t_L g4155 ( 
.A1(n_4135),
.A2(n_3919),
.B(n_3942),
.C(n_3876),
.Y(n_4155)
);

AOI221x1_ASAP7_75t_L g4156 ( 
.A1(n_4138),
.A2(n_3916),
.B1(n_3931),
.B2(n_3913),
.C(n_3942),
.Y(n_4156)
);

O2A1O1Ixp33_ASAP7_75t_L g4157 ( 
.A1(n_4136),
.A2(n_3895),
.B(n_3933),
.C(n_3934),
.Y(n_4157)
);

INVxp67_ASAP7_75t_SL g4158 ( 
.A(n_4149),
.Y(n_4158)
);

AOI22xp5_ASAP7_75t_L g4159 ( 
.A1(n_4144),
.A2(n_3945),
.B1(n_3944),
.B2(n_3839),
.Y(n_4159)
);

A2O1A1Ixp33_ASAP7_75t_SL g4160 ( 
.A1(n_4129),
.A2(n_3942),
.B(n_3910),
.C(n_3908),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_SL g4161 ( 
.A(n_4148),
.B(n_3942),
.Y(n_4161)
);

INVx2_ASAP7_75t_L g4162 ( 
.A(n_4150),
.Y(n_4162)
);

AOI221xp5_ASAP7_75t_L g4163 ( 
.A1(n_4133),
.A2(n_3906),
.B1(n_3914),
.B2(n_3942),
.C(n_3913),
.Y(n_4163)
);

AOI222xp33_ASAP7_75t_L g4164 ( 
.A1(n_4151),
.A2(n_3914),
.B1(n_3906),
.B2(n_3937),
.C1(n_3934),
.C2(n_3933),
.Y(n_4164)
);

OAI211xp5_ASAP7_75t_SL g4165 ( 
.A1(n_4131),
.A2(n_3931),
.B(n_3916),
.C(n_3910),
.Y(n_4165)
);

AOI22xp5_ASAP7_75t_L g4166 ( 
.A1(n_4145),
.A2(n_3945),
.B1(n_3944),
.B2(n_3838),
.Y(n_4166)
);

O2A1O1Ixp33_ASAP7_75t_L g4167 ( 
.A1(n_4143),
.A2(n_3895),
.B(n_3934),
.C(n_3933),
.Y(n_4167)
);

O2A1O1Ixp5_ASAP7_75t_SL g4168 ( 
.A1(n_4134),
.A2(n_3867),
.B(n_3871),
.C(n_3876),
.Y(n_4168)
);

OAI211xp5_ASAP7_75t_L g4169 ( 
.A1(n_4147),
.A2(n_4142),
.B(n_4141),
.C(n_4152),
.Y(n_4169)
);

NAND3xp33_ASAP7_75t_L g4170 ( 
.A(n_4154),
.B(n_4146),
.C(n_4140),
.Y(n_4170)
);

OR2x2_ASAP7_75t_L g4171 ( 
.A(n_4159),
.B(n_3838),
.Y(n_4171)
);

NAND4xp25_ASAP7_75t_SL g4172 ( 
.A(n_4166),
.B(n_4139),
.C(n_3867),
.D(n_3877),
.Y(n_4172)
);

INVxp67_ASAP7_75t_L g4173 ( 
.A(n_4161),
.Y(n_4173)
);

NAND3xp33_ASAP7_75t_SL g4174 ( 
.A(n_4168),
.B(n_3848),
.C(n_3937),
.Y(n_4174)
);

NOR4xp75_ASAP7_75t_L g4175 ( 
.A(n_4169),
.B(n_4137),
.C(n_3845),
.D(n_3850),
.Y(n_4175)
);

AOI221xp5_ASAP7_75t_L g4176 ( 
.A1(n_4163),
.A2(n_3906),
.B1(n_3914),
.B2(n_3923),
.C(n_3924),
.Y(n_4176)
);

NAND3xp33_ASAP7_75t_L g4177 ( 
.A(n_4162),
.B(n_3871),
.C(n_3889),
.Y(n_4177)
);

INVxp67_ASAP7_75t_L g4178 ( 
.A(n_4158),
.Y(n_4178)
);

NAND4xp25_ASAP7_75t_L g4179 ( 
.A(n_4153),
.B(n_3906),
.C(n_3914),
.D(n_3923),
.Y(n_4179)
);

NOR2x1_ASAP7_75t_L g4180 ( 
.A(n_4165),
.B(n_3933),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_L g4181 ( 
.A(n_4164),
.B(n_3839),
.Y(n_4181)
);

NAND3xp33_ASAP7_75t_SL g4182 ( 
.A(n_4157),
.B(n_3848),
.C(n_3934),
.Y(n_4182)
);

NAND3xp33_ASAP7_75t_SL g4183 ( 
.A(n_4160),
.B(n_3937),
.C(n_3889),
.Y(n_4183)
);

OAI322xp33_ASAP7_75t_L g4184 ( 
.A1(n_4167),
.A2(n_3924),
.A3(n_3923),
.B1(n_3910),
.B2(n_3908),
.C1(n_3937),
.C2(n_3853),
.Y(n_4184)
);

NAND4xp25_ASAP7_75t_L g4185 ( 
.A(n_4177),
.B(n_4156),
.C(n_4155),
.D(n_3924),
.Y(n_4185)
);

AOI221x1_ASAP7_75t_L g4186 ( 
.A1(n_4170),
.A2(n_3924),
.B1(n_3923),
.B2(n_3910),
.C(n_3908),
.Y(n_4186)
);

NAND4xp25_ASAP7_75t_L g4187 ( 
.A(n_4176),
.B(n_3908),
.C(n_3853),
.D(n_3850),
.Y(n_4187)
);

NAND3xp33_ASAP7_75t_L g4188 ( 
.A(n_4178),
.B(n_3895),
.C(n_3866),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_4183),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_L g4190 ( 
.A(n_4173),
.B(n_3739),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_4171),
.B(n_3739),
.Y(n_4191)
);

AOI22xp5_ASAP7_75t_L g4192 ( 
.A1(n_4172),
.A2(n_3884),
.B1(n_3895),
.B2(n_3869),
.Y(n_4192)
);

OAI221xp5_ASAP7_75t_L g4193 ( 
.A1(n_4179),
.A2(n_3895),
.B1(n_3849),
.B2(n_3870),
.C(n_3872),
.Y(n_4193)
);

NOR2xp33_ASAP7_75t_L g4194 ( 
.A(n_4181),
.B(n_3895),
.Y(n_4194)
);

OAI211xp5_ASAP7_75t_L g4195 ( 
.A1(n_4180),
.A2(n_3854),
.B(n_3870),
.C(n_3872),
.Y(n_4195)
);

NAND2xp5_ASAP7_75t_L g4196 ( 
.A(n_4182),
.B(n_3746),
.Y(n_4196)
);

OAI21xp5_ASAP7_75t_L g4197 ( 
.A1(n_4174),
.A2(n_3854),
.B(n_3874),
.Y(n_4197)
);

NAND4xp25_ASAP7_75t_L g4198 ( 
.A(n_4175),
.B(n_3854),
.C(n_3888),
.D(n_3886),
.Y(n_4198)
);

NAND3xp33_ASAP7_75t_SL g4199 ( 
.A(n_4184),
.B(n_3874),
.C(n_3870),
.Y(n_4199)
);

NAND4xp25_ASAP7_75t_L g4200 ( 
.A(n_4177),
.B(n_3890),
.C(n_3888),
.D(n_3886),
.Y(n_4200)
);

OAI211xp5_ASAP7_75t_SL g4201 ( 
.A1(n_4178),
.A2(n_3746),
.B(n_3749),
.C(n_3793),
.Y(n_4201)
);

OAI21xp33_ASAP7_75t_L g4202 ( 
.A1(n_4181),
.A2(n_3890),
.B(n_3888),
.Y(n_4202)
);

OAI21xp33_ASAP7_75t_SL g4203 ( 
.A1(n_4192),
.A2(n_3872),
.B(n_3874),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4202),
.Y(n_4204)
);

CKINVDCx5p33_ASAP7_75t_R g4205 ( 
.A(n_4190),
.Y(n_4205)
);

NOR2x1_ASAP7_75t_L g4206 ( 
.A(n_4185),
.B(n_3884),
.Y(n_4206)
);

NOR2x1_ASAP7_75t_L g4207 ( 
.A(n_4188),
.B(n_3884),
.Y(n_4207)
);

BUFx6f_ASAP7_75t_L g4208 ( 
.A(n_4189),
.Y(n_4208)
);

NOR2xp33_ASAP7_75t_SL g4209 ( 
.A(n_4194),
.B(n_3884),
.Y(n_4209)
);

INVx2_ASAP7_75t_L g4210 ( 
.A(n_4191),
.Y(n_4210)
);

INVxp33_ASAP7_75t_SL g4211 ( 
.A(n_4196),
.Y(n_4211)
);

NOR2xp67_ASAP7_75t_L g4212 ( 
.A(n_4187),
.B(n_3749),
.Y(n_4212)
);

NOR2x1_ASAP7_75t_L g4213 ( 
.A(n_4199),
.B(n_3861),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_4197),
.Y(n_4214)
);

NOR2x1_ASAP7_75t_L g4215 ( 
.A(n_4195),
.B(n_3861),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_4201),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_4200),
.Y(n_4217)
);

NOR2x1_ASAP7_75t_L g4218 ( 
.A(n_4198),
.B(n_3861),
.Y(n_4218)
);

INVxp33_ASAP7_75t_SL g4219 ( 
.A(n_4186),
.Y(n_4219)
);

NAND5xp2_ASAP7_75t_L g4220 ( 
.A(n_4209),
.B(n_4193),
.C(n_3875),
.D(n_3885),
.E(n_3881),
.Y(n_4220)
);

NOR2x1_ASAP7_75t_L g4221 ( 
.A(n_4206),
.B(n_3861),
.Y(n_4221)
);

NAND4xp75_ASAP7_75t_L g4222 ( 
.A(n_4204),
.B(n_3885),
.C(n_3881),
.D(n_3875),
.Y(n_4222)
);

AND2x4_ASAP7_75t_L g4223 ( 
.A(n_4212),
.B(n_3831),
.Y(n_4223)
);

AOI31xp33_ASAP7_75t_L g4224 ( 
.A1(n_4216),
.A2(n_3885),
.A3(n_3881),
.B(n_3875),
.Y(n_4224)
);

NAND4xp25_ASAP7_75t_L g4225 ( 
.A(n_4217),
.B(n_4218),
.C(n_4213),
.D(n_4207),
.Y(n_4225)
);

NOR2x1_ASAP7_75t_L g4226 ( 
.A(n_4215),
.B(n_3813),
.Y(n_4226)
);

INVx2_ASAP7_75t_L g4227 ( 
.A(n_4208),
.Y(n_4227)
);

NAND2x1p5_ASAP7_75t_L g4228 ( 
.A(n_4208),
.B(n_3813),
.Y(n_4228)
);

NAND2x1p5_ASAP7_75t_L g4229 ( 
.A(n_4210),
.B(n_3813),
.Y(n_4229)
);

NAND4xp75_ASAP7_75t_L g4230 ( 
.A(n_4214),
.B(n_3890),
.C(n_3886),
.D(n_3786),
.Y(n_4230)
);

AOI211xp5_ASAP7_75t_L g4231 ( 
.A1(n_4225),
.A2(n_4203),
.B(n_4205),
.C(n_4219),
.Y(n_4231)
);

OAI211xp5_ASAP7_75t_SL g4232 ( 
.A1(n_4227),
.A2(n_4211),
.B(n_3786),
.C(n_3793),
.Y(n_4232)
);

AND2x4_ASAP7_75t_L g4233 ( 
.A(n_4223),
.B(n_3831),
.Y(n_4233)
);

XNOR2xp5_ASAP7_75t_L g4234 ( 
.A(n_4228),
.B(n_3710),
.Y(n_4234)
);

NAND3xp33_ASAP7_75t_SL g4235 ( 
.A(n_4229),
.B(n_3804),
.C(n_3800),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_4226),
.Y(n_4236)
);

OR2x2_ASAP7_75t_L g4237 ( 
.A(n_4235),
.B(n_4224),
.Y(n_4237)
);

AOI22xp33_ASAP7_75t_L g4238 ( 
.A1(n_4233),
.A2(n_4220),
.B1(n_4221),
.B2(n_4230),
.Y(n_4238)
);

AND2x4_ASAP7_75t_L g4239 ( 
.A(n_4236),
.B(n_3831),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4239),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_4237),
.Y(n_4241)
);

AOI21x1_ASAP7_75t_L g4242 ( 
.A1(n_4240),
.A2(n_4234),
.B(n_4231),
.Y(n_4242)
);

BUFx3_ASAP7_75t_L g4243 ( 
.A(n_4242),
.Y(n_4243)
);

INVx2_ASAP7_75t_L g4244 ( 
.A(n_4243),
.Y(n_4244)
);

INVxp67_ASAP7_75t_SL g4245 ( 
.A(n_4244),
.Y(n_4245)
);

OAI21xp5_ASAP7_75t_L g4246 ( 
.A1(n_4245),
.A2(n_4241),
.B(n_4238),
.Y(n_4246)
);

XOR2xp5_ASAP7_75t_L g4247 ( 
.A(n_4246),
.B(n_4222),
.Y(n_4247)
);

AOI22xp5_ASAP7_75t_L g4248 ( 
.A1(n_4247),
.A2(n_4232),
.B1(n_3869),
.B2(n_3800),
.Y(n_4248)
);

INVxp67_ASAP7_75t_L g4249 ( 
.A(n_4248),
.Y(n_4249)
);

OAI21xp33_ASAP7_75t_L g4250 ( 
.A1(n_4249),
.A2(n_3869),
.B(n_3804),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4250),
.Y(n_4251)
);

AO221x2_ASAP7_75t_L g4252 ( 
.A1(n_4251),
.A2(n_3827),
.B1(n_3809),
.B2(n_3805),
.C(n_3806),
.Y(n_4252)
);

XNOR2x1_ASAP7_75t_L g4253 ( 
.A(n_4251),
.B(n_3869),
.Y(n_4253)
);

OAI221xp5_ASAP7_75t_R g4254 ( 
.A1(n_4253),
.A2(n_3835),
.B1(n_3869),
.B2(n_3814),
.C(n_3827),
.Y(n_4254)
);

AOI221xp5_ASAP7_75t_L g4255 ( 
.A1(n_4252),
.A2(n_3810),
.B1(n_3789),
.B2(n_3787),
.C(n_3782),
.Y(n_4255)
);

AOI22xp33_ASAP7_75t_L g4256 ( 
.A1(n_4255),
.A2(n_3814),
.B1(n_3805),
.B2(n_3809),
.Y(n_4256)
);

AOI211xp5_ASAP7_75t_L g4257 ( 
.A1(n_4256),
.A2(n_4254),
.B(n_3797),
.C(n_3778),
.Y(n_4257)
);


endmodule