module fake_jpeg_972_n_503 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_503);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_503;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_54),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_56),
.B(n_84),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_57),
.Y(n_171)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_60),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_61),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_63),
.B(n_70),
.Y(n_135)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_64),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_66),
.Y(n_172)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_67),
.Y(n_176)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_69),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_37),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_71),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_72),
.Y(n_189)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_73),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_37),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_74),
.B(n_79),
.Y(n_144)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_76),
.Y(n_178)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_78),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_82),
.Y(n_193)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_83),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_38),
.B(n_17),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_85),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_44),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_89),
.B(n_93),
.Y(n_168)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_90),
.Y(n_199)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

BUFx8_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

BUFx4f_ASAP7_75t_SL g93 ( 
.A(n_20),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_17),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_104),
.Y(n_140)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_49),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_101),
.B(n_114),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_19),
.B(n_27),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_43),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_105),
.B(n_118),
.Y(n_156)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_106),
.Y(n_175)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

BUFx4f_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_108),
.Y(n_184)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_109),
.Y(n_191)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_110),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_24),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_45),
.B(n_15),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_116),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_41),
.Y(n_113)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_113),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_41),
.B(n_16),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g115 ( 
.A(n_45),
.Y(n_115)
);

BUFx2_ASAP7_75t_R g150 ( 
.A(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_19),
.B(n_14),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_21),
.Y(n_117)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_21),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_47),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_119),
.B(n_93),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_23),
.Y(n_120)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_92),
.A2(n_47),
.B1(n_46),
.B2(n_39),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g205 ( 
.A1(n_125),
.A2(n_131),
.B1(n_162),
.B2(n_174),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_62),
.A2(n_46),
.B1(n_39),
.B2(n_52),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_128),
.A2(n_155),
.B1(n_173),
.B2(n_179),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_114),
.B(n_23),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_129),
.B(n_152),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_69),
.A2(n_24),
.B1(n_50),
.B2(n_42),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_132),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_61),
.B(n_52),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_136),
.B(n_159),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_118),
.B(n_35),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_65),
.A2(n_50),
.B1(n_42),
.B2(n_40),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_73),
.A2(n_94),
.B1(n_83),
.B2(n_66),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_157),
.A2(n_181),
.B1(n_185),
.B2(n_143),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_76),
.A2(n_40),
.B1(n_35),
.B2(n_34),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_61),
.A2(n_34),
.B1(n_33),
.B2(n_27),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_111),
.B(n_33),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_156),
.Y(n_214)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_169),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_72),
.A2(n_25),
.B1(n_2),
.B2(n_3),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_91),
.A2(n_25),
.B1(n_3),
.B2(n_5),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_86),
.A2(n_13),
.B1(n_3),
.B2(n_5),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_113),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_82),
.A2(n_1),
.B1(n_6),
.B2(n_7),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_182),
.A2(n_200),
.B1(n_146),
.B2(n_143),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_102),
.A2(n_111),
.B1(n_60),
.B2(n_59),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_96),
.Y(n_186)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_186),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_71),
.A2(n_13),
.B1(n_6),
.B2(n_9),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_187),
.A2(n_75),
.B1(n_78),
.B2(n_107),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_196),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_98),
.B(n_1),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_136),
.Y(n_224)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_57),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_109),
.A2(n_6),
.B(n_9),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_198),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_82),
.A2(n_10),
.B1(n_11),
.B2(n_110),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_203),
.A2(n_226),
.B1(n_229),
.B2(n_259),
.Y(n_283)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_204),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_206),
.Y(n_307)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_207),
.Y(n_296)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_208),
.Y(n_320)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_133),
.B(n_10),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_212),
.B(n_234),
.C(n_256),
.Y(n_271)
);

OR2x4_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_11),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_L g300 ( 
.A1(n_213),
.A2(n_214),
.B(n_244),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_135),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_215),
.B(n_224),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_126),
.Y(n_217)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_217),
.Y(n_274)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_158),
.Y(n_218)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_218),
.Y(n_303)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_219),
.Y(n_305)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_221),
.Y(n_281)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_222),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_223),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_168),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_225),
.B(n_228),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_200),
.B1(n_131),
.B2(n_162),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_121),
.B(n_140),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_233),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_142),
.B(n_144),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_134),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_230),
.Y(n_311)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_231),
.Y(n_294)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_232),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_122),
.B(n_123),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_130),
.B(n_163),
.C(n_153),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_141),
.Y(n_235)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_235),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_134),
.Y(n_236)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_236),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_132),
.B(n_167),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_238),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_145),
.B(n_126),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_160),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_239),
.B(n_248),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_180),
.Y(n_240)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_240),
.Y(n_312)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_166),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_241),
.B(n_242),
.Y(n_290)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_146),
.A2(n_147),
.B1(n_199),
.B2(n_171),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_243),
.A2(n_247),
.B1(n_252),
.B2(n_260),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_154),
.B(n_176),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_180),
.Y(n_246)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_246),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_146),
.A2(n_147),
.B1(n_171),
.B2(n_175),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_150),
.B(n_183),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_124),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_249),
.B(n_253),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_181),
.B(n_137),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_258),
.Y(n_277)
);

OR2x4_ASAP7_75t_L g251 ( 
.A(n_155),
.B(n_125),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_251),
.A2(n_205),
.B(n_216),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_178),
.A2(n_188),
.B1(n_177),
.B2(n_192),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_139),
.B(n_148),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_160),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_254),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_149),
.B(n_178),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_138),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_257),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_138),
.Y(n_258)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_193),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_191),
.B(n_127),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_262),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_128),
.B(n_173),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_161),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_263),
.A2(n_264),
.B1(n_269),
.B2(n_217),
.Y(n_295)
);

BUFx12f_ASAP7_75t_L g264 ( 
.A(n_161),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_172),
.B(n_189),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_266),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_127),
.B(n_172),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_189),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_267),
.B(n_270),
.Y(n_304)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_127),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_182),
.B(n_174),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_250),
.A2(n_164),
.B1(n_255),
.B2(n_229),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_272),
.A2(n_276),
.B1(n_284),
.B2(n_287),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_255),
.A2(n_164),
.B1(n_262),
.B2(n_251),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_214),
.A2(n_209),
.B(n_270),
.Y(n_279)
);

OA21x2_ASAP7_75t_L g325 ( 
.A1(n_279),
.A2(n_221),
.B(n_264),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_234),
.B(n_220),
.C(n_233),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_280),
.B(n_301),
.C(n_318),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_283),
.A2(n_309),
.B1(n_310),
.B2(n_314),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_209),
.A2(n_212),
.B1(n_226),
.B2(n_205),
.Y(n_284)
);

OAI32xp33_ASAP7_75t_L g286 ( 
.A1(n_227),
.A2(n_213),
.A3(n_210),
.B1(n_212),
.B2(n_205),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_286),
.B(n_317),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_205),
.A2(n_203),
.B1(n_232),
.B2(n_231),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_292),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_295),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_245),
.B(n_256),
.C(n_268),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_219),
.A2(n_222),
.B1(n_211),
.B2(n_242),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_263),
.A2(n_208),
.B1(n_207),
.B2(n_204),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_256),
.A2(n_218),
.B1(n_241),
.B2(n_206),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_235),
.A2(n_249),
.B1(n_264),
.B2(n_240),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_315),
.A2(n_308),
.B1(n_287),
.B2(n_284),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_260),
.B(n_230),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_236),
.B(n_246),
.C(n_269),
.Y(n_318)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_290),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_322),
.B(n_330),
.Y(n_366)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_294),
.Y(n_323)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_323),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_324),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_325),
.A2(n_281),
.B(n_299),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_273),
.B(n_221),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g361 ( 
.A(n_326),
.Y(n_361)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_294),
.Y(n_327)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_327),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_275),
.B(n_280),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_328),
.B(n_336),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_290),
.Y(n_330)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_335),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_278),
.B(n_285),
.Y(n_337)
);

BUFx24_ASAP7_75t_SL g363 ( 
.A(n_337),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_283),
.A2(n_289),
.B1(n_304),
.B2(n_277),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_338),
.A2(n_351),
.B1(n_357),
.B2(n_318),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_297),
.B(n_275),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_340),
.A2(n_334),
.B1(n_333),
.B2(n_325),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_308),
.A2(n_276),
.B1(n_272),
.B2(n_304),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_341),
.A2(n_356),
.B1(n_315),
.B2(n_299),
.Y(n_376)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_298),
.Y(n_342)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_342),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_279),
.B(n_302),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_345),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_290),
.Y(n_344)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_289),
.B(n_286),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_305),
.Y(n_346)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_346),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_311),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_347),
.B(n_349),
.Y(n_375)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_306),
.Y(n_348)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_348),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_277),
.B(n_292),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_350),
.B(n_352),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_302),
.A2(n_319),
.B1(n_282),
.B2(n_271),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_314),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_271),
.B(n_301),
.Y(n_353)
);

NOR2x1_ASAP7_75t_L g365 ( 
.A(n_353),
.B(n_281),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_311),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_355),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_274),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_307),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_300),
.A2(n_316),
.B1(n_288),
.B2(n_313),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_274),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_355),
.Y(n_385)
);

AOI221xp5_ASAP7_75t_L g390 ( 
.A1(n_359),
.A2(n_343),
.B1(n_338),
.B2(n_357),
.C(n_321),
.Y(n_390)
);

OAI21xp33_ASAP7_75t_L g410 ( 
.A1(n_365),
.A2(n_386),
.B(n_389),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_293),
.C(n_296),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_367),
.B(n_379),
.C(n_330),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_344),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_329),
.A2(n_313),
.B1(n_312),
.B2(n_320),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_372),
.A2(n_383),
.B1(n_384),
.B2(n_388),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_374),
.A2(n_324),
.B(n_356),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_376),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_336),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_329),
.A2(n_312),
.B1(n_320),
.B2(n_296),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_349),
.A2(n_291),
.B1(n_293),
.B2(n_332),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_385),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_333),
.A2(n_291),
.B(n_325),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_345),
.A2(n_332),
.B(n_351),
.Y(n_389)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_390),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_384),
.Y(n_391)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_400),
.C(n_379),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_394),
.B(n_389),
.Y(n_419)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_362),
.Y(n_395)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_395),
.Y(n_425)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_362),
.Y(n_397)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_397),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_371),
.B(n_354),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_399),
.Y(n_423)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_375),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_347),
.C(n_350),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_371),
.B(n_348),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_401),
.B(n_406),
.Y(n_436)
);

BUFx24_ASAP7_75t_SL g402 ( 
.A(n_363),
.Y(n_402)
);

BUFx24_ASAP7_75t_SL g428 ( 
.A(n_402),
.Y(n_428)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_378),
.Y(n_403)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_403),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_359),
.A2(n_352),
.B1(n_334),
.B2(n_331),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_404),
.A2(n_408),
.B1(n_409),
.B2(n_411),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_378),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_412),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_364),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_365),
.B(n_323),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_407),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_375),
.A2(n_360),
.B1(n_372),
.B2(n_383),
.Y(n_408)
);

OAI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_361),
.A2(n_358),
.B1(n_327),
.B2(n_342),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_369),
.A2(n_346),
.B1(n_335),
.B2(n_324),
.Y(n_411)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_382),
.Y(n_414)
);

BUFx4f_ASAP7_75t_SL g434 ( 
.A(n_414),
.Y(n_434)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_415),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_417),
.B(n_404),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_407),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_418),
.B(n_364),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_419),
.B(n_421),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_400),
.B(n_367),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_394),
.B(n_369),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_427),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_393),
.B(n_366),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_396),
.B(n_381),
.C(n_386),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_433),
.B(n_419),
.C(n_417),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_410),
.B(n_381),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_435),
.B(n_437),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_364),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_440),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_416),
.A2(n_413),
.B(n_396),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_439),
.B(n_445),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_422),
.A2(n_392),
.B1(n_406),
.B2(n_413),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_441),
.A2(n_448),
.B1(n_449),
.B2(n_432),
.Y(n_460)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_423),
.Y(n_442)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_442),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_433),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_443),
.B(n_446),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_420),
.A2(n_374),
.B(n_412),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_380),
.C(n_392),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_447),
.B(n_440),
.C(n_443),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_432),
.A2(n_436),
.B1(n_424),
.B2(n_435),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_422),
.A2(n_408),
.B1(n_405),
.B2(n_395),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_380),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_451),
.B(n_453),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_377),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_426),
.B(n_387),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_454),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_456),
.B(n_457),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_450),
.B(n_437),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_380),
.C(n_432),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_459),
.B(n_464),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_460),
.A2(n_434),
.B1(n_397),
.B2(n_414),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_434),
.Y(n_463)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_463),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_441),
.A2(n_385),
.B(n_431),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_385),
.C(n_405),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_465),
.B(n_452),
.C(n_444),
.Y(n_473)
);

OAI22xp33_ASAP7_75t_L g468 ( 
.A1(n_463),
.A2(n_448),
.B1(n_425),
.B2(n_430),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_468),
.B(n_469),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_461),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_467),
.B(n_447),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_475),
.C(n_459),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_474),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_452),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_444),
.C(n_403),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_476),
.B(n_478),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_458),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_477),
.B(n_475),
.C(n_456),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_482),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_467),
.Y(n_483)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_483),
.Y(n_488)
);

MAJx2_ASAP7_75t_L g485 ( 
.A(n_473),
.B(n_457),
.C(n_458),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_485),
.B(n_474),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_466),
.Y(n_486)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_486),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_489),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_479),
.B(n_434),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_484),
.A2(n_468),
.B(n_465),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_490),
.A2(n_464),
.B(n_460),
.Y(n_493)
);

AO21x1_ASAP7_75t_L g498 ( 
.A1(n_493),
.A2(n_496),
.B(n_489),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_492),
.B(n_481),
.Y(n_495)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_495),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_488),
.B(n_491),
.Y(n_496)
);

AOI321xp33_ASAP7_75t_L g499 ( 
.A1(n_498),
.A2(n_494),
.A3(n_485),
.B1(n_480),
.B2(n_415),
.C(n_387),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_499),
.A2(n_497),
.B1(n_373),
.B2(n_370),
.Y(n_500)
);

OA21x2_ASAP7_75t_SL g501 ( 
.A1(n_500),
.A2(n_373),
.B(n_370),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_501),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_502),
.A2(n_356),
.B(n_428),
.Y(n_503)
);


endmodule