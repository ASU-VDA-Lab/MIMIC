module fake_jpeg_16156_n_150 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_150);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_30),
.A2(n_35),
.B(n_23),
.Y(n_44)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_19),
.B(n_2),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_2),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_15),
.B1(n_14),
.B2(n_25),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_41),
.B1(n_48),
.B2(n_49),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_16),
.B1(n_25),
.B2(n_17),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_26),
.C(n_14),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_2),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_23),
.B1(n_16),
.B2(n_17),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_32),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_27),
.B1(n_22),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_31),
.A2(n_24),
.B1(n_20),
.B2(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_52),
.B(n_62),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_57),
.B1(n_3),
.B2(n_20),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_65),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_64),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_3),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_33),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_34),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_37),
.B1(n_40),
.B2(n_39),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_67),
.A2(n_74),
.B1(n_75),
.B2(n_58),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_57),
.B(n_53),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_82),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_40),
.B1(n_37),
.B2(n_38),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_34),
.B1(n_26),
.B2(n_47),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_79),
.Y(n_92)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_47),
.C(n_34),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_83),
.B(n_67),
.Y(n_102)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_71),
.B(n_57),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_79),
.B(n_70),
.Y(n_100)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_78),
.A2(n_53),
.B(n_60),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_96),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_76),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_95),
.B(n_68),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_99),
.B(n_107),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_104),
.C(n_83),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_80),
.B(n_75),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_101),
.Y(n_114)
);

OAI322xp33_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_91),
.A3(n_93),
.B1(n_85),
.B2(n_84),
.C1(n_94),
.C2(n_87),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_21),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_5),
.B(n_6),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_89),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_116),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_98),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_120),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_116),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_88),
.C(n_85),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_96),
.C(n_86),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_128),
.C(n_110),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_117),
.Y(n_129)
);

XOR2x2_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_114),
.C(n_118),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

NAND2x1p5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_103),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_132),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_130),
.C(n_126),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_125),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_142),
.C(n_143),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_141),
.A2(n_138),
.B1(n_137),
.B2(n_97),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_90),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_86),
.C(n_89),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_147),
.C(n_10),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_9),
.C(n_10),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_11),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_12),
.Y(n_150)
);


endmodule