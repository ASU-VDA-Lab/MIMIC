module fake_netlist_6_4830_n_1661 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1661);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1661;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_17),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_65),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_50),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_28),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_118),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_37),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_74),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_67),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_31),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_43),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_36),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_108),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_69),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_39),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_78),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_113),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_88),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_143),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_10),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_95),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_102),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_144),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_2),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_155),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_75),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_98),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_112),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_21),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_131),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_18),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_9),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_129),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_52),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_63),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_15),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_61),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g198 ( 
.A(n_3),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_29),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_5),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_140),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_28),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_56),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_62),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_120),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_76),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_115),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_64),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_4),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_142),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_14),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_41),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_101),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_146),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_111),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_82),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_57),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_77),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_123),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_110),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_56),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_133),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_128),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_91),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_71),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_89),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_154),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_60),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_157),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_106),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_39),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_16),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_58),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_43),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_24),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_19),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_8),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_35),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_26),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_68),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_34),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_125),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_148),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_86),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_19),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_130),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_47),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_23),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_11),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_83),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_35),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_85),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_26),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_134),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_79),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_150),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_15),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_46),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_12),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_107),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_17),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_31),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_8),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_0),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_117),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_94),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_32),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_50),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_59),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_52),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_149),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_137),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_66),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_48),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_11),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_27),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_153),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_124),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_109),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_141),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_13),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_1),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_114),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_14),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_47),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_96),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_36),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_41),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_21),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_44),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_104),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_48),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_22),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_37),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_45),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_16),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_38),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_135),
.Y(n_299)
);

BUFx5_ASAP7_75t_L g300 ( 
.A(n_46),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_99),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_105),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_13),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_100),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_72),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_44),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_27),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_80),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_0),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_145),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_32),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_33),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_20),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_84),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_192),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_272),
.B(n_1),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_300),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_194),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_202),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_159),
.B(n_2),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_200),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_3),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_205),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_300),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_244),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_300),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_300),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_196),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_206),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_208),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_300),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_300),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_263),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_203),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_L g335 ( 
.A(n_168),
.B(n_4),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_300),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_211),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_214),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_158),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_238),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_158),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_215),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_216),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_158),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_158),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_158),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_219),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_R g348 ( 
.A(n_165),
.B(n_138),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_307),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_307),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_280),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_176),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_221),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_307),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_184),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_223),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_160),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_307),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_218),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_159),
.B(n_5),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_311),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_R g363 ( 
.A(n_163),
.B(n_6),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_226),
.B(n_6),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_225),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_228),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_L g367 ( 
.A(n_173),
.B(n_7),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_311),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_311),
.Y(n_369)
);

INVxp33_ASAP7_75t_L g370 ( 
.A(n_191),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_226),
.B(n_7),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_311),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_230),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_311),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_201),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_234),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_238),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_210),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_255),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_196),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_212),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_243),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_222),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_251),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_232),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_237),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_246),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_253),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_227),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_248),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_353),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_328),
.B(n_247),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_315),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_324),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_339),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_320),
.B(n_247),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_358),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_324),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_339),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_L g400 ( 
.A(n_348),
.B(n_160),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_356),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_317),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_317),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_341),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_341),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_318),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_319),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_326),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_326),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_361),
.B(n_163),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_360),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_333),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g413 ( 
.A(n_327),
.B(n_162),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_323),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_329),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_327),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_371),
.B(n_171),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_330),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_R g420 ( 
.A(n_382),
.B(n_257),
.Y(n_420)
);

CKINVDCx6p67_ASAP7_75t_R g421 ( 
.A(n_325),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_331),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_344),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_345),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_379),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_R g426 ( 
.A(n_384),
.B(n_267),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_331),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_345),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_337),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_338),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_332),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_342),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_343),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_346),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_346),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_389),
.B(n_238),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_349),
.B(n_171),
.Y(n_437)
);

NAND2xp33_ASAP7_75t_R g438 ( 
.A(n_347),
.B(n_172),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_349),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_380),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_350),
.Y(n_441)
);

INVxp33_ASAP7_75t_SL g442 ( 
.A(n_354),
.Y(n_442)
);

AND3x2_ASAP7_75t_L g443 ( 
.A(n_316),
.B(n_287),
.C(n_166),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_332),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_357),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_350),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_380),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_336),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_365),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_377),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_336),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_R g452 ( 
.A(n_366),
.B(n_273),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_351),
.B(n_172),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_351),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_355),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_340),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_355),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_359),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_359),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_362),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_362),
.B(n_174),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_373),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_402),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_394),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_410),
.A2(n_364),
.B1(n_352),
.B2(n_389),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_420),
.Y(n_466)
);

AND2x6_ASAP7_75t_L g467 ( 
.A(n_427),
.B(n_166),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_392),
.B(n_368),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_412),
.B(n_321),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_440),
.Y(n_470)
);

INVx6_ASAP7_75t_L g471 ( 
.A(n_417),
.Y(n_471)
);

AND2x2_ASAP7_75t_SL g472 ( 
.A(n_396),
.B(n_287),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_396),
.B(n_376),
.Y(n_473)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_413),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_456),
.B(n_388),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_394),
.Y(n_476)
);

INVx6_ASAP7_75t_L g477 ( 
.A(n_417),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_392),
.B(n_368),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_402),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_456),
.B(n_321),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_394),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_442),
.B(n_340),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_412),
.B(n_334),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_417),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_398),
.Y(n_485)
);

AND3x2_ASAP7_75t_L g486 ( 
.A(n_436),
.B(n_305),
.C(n_304),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_447),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_410),
.A2(n_322),
.B1(n_367),
.B2(n_335),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_402),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_417),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_418),
.B(n_369),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_417),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_418),
.B(n_369),
.Y(n_493)
);

BUFx6f_ASAP7_75t_SL g494 ( 
.A(n_447),
.Y(n_494)
);

NAND3xp33_ASAP7_75t_L g495 ( 
.A(n_397),
.B(n_363),
.C(n_370),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_L g496 ( 
.A(n_413),
.B(n_162),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_447),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_436),
.B(n_227),
.Y(n_498)
);

INVx4_ASAP7_75t_L g499 ( 
.A(n_417),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_398),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_458),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_458),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_393),
.B(n_217),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_403),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_458),
.Y(n_505)
);

AND2x6_ASAP7_75t_L g506 ( 
.A(n_427),
.B(n_304),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_391),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_403),
.Y(n_508)
);

BUFx6f_ASAP7_75t_SL g509 ( 
.A(n_421),
.Y(n_509)
);

BUFx4f_ASAP7_75t_L g510 ( 
.A(n_413),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_403),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_423),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_452),
.B(n_227),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_426),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_427),
.A2(n_298),
.B1(n_293),
.B2(n_254),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_440),
.B(n_372),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_408),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_427),
.B(n_372),
.Y(n_518)
);

INVx4_ASAP7_75t_SL g519 ( 
.A(n_413),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_444),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_408),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_408),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_443),
.B(n_199),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_444),
.B(n_374),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_406),
.B(n_174),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_437),
.B(n_453),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_423),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_401),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_407),
.B(n_175),
.Y(n_529)
);

INVx6_ASAP7_75t_L g530 ( 
.A(n_423),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_444),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_414),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_438),
.A2(n_187),
.B1(n_186),
.B2(n_183),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_409),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_SL g535 ( 
.A1(n_450),
.A2(n_239),
.B1(n_252),
.B2(n_250),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_421),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_413),
.Y(n_537)
);

INVx5_ASAP7_75t_L g538 ( 
.A(n_413),
.Y(n_538)
);

BUFx10_ASAP7_75t_L g539 ( 
.A(n_415),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_462),
.B(n_261),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_409),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_409),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_443),
.B(n_199),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_444),
.B(n_374),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_416),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_419),
.B(n_175),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_450),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_416),
.Y(n_548)
);

BUFx4f_ASAP7_75t_L g549 ( 
.A(n_413),
.Y(n_549)
);

AO22x2_ASAP7_75t_L g550 ( 
.A1(n_397),
.A2(n_306),
.B1(n_198),
.B2(n_305),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_429),
.B(n_177),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_416),
.A2(n_269),
.B1(n_259),
.B2(n_260),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_430),
.B(n_261),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_432),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_433),
.B(n_177),
.Y(n_555)
);

INVxp33_ASAP7_75t_L g556 ( 
.A(n_437),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_422),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_445),
.B(n_261),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_453),
.B(n_375),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_422),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_461),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_422),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_411),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_461),
.B(n_421),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_449),
.B(n_179),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_431),
.B(n_301),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_431),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_460),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_423),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_431),
.B(n_270),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_448),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_448),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_448),
.B(n_270),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_395),
.B(n_375),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_395),
.B(n_301),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_399),
.B(n_378),
.Y(n_576)
);

BUFx4f_ASAP7_75t_L g577 ( 
.A(n_413),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_451),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_451),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_425),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_451),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_399),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_404),
.B(n_274),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_423),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_400),
.B(n_179),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_404),
.B(n_378),
.Y(n_586)
);

BUFx8_ASAP7_75t_SL g587 ( 
.A(n_423),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_405),
.B(n_278),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_405),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_424),
.B(n_270),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_424),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_413),
.A2(n_303),
.B1(n_262),
.B2(n_265),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_441),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_428),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_428),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_434),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_434),
.A2(n_180),
.B1(n_292),
.B2(n_187),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_435),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_435),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_441),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_441),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_441),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_441),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_439),
.B(n_180),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_441),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_439),
.B(n_446),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_446),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_454),
.B(n_381),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_454),
.B(n_181),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_455),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_455),
.B(n_181),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_457),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_561),
.A2(n_207),
.B1(n_170),
.B2(n_185),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_516),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_472),
.A2(n_285),
.B1(n_291),
.B2(n_313),
.Y(n_615)
);

OAI22xp33_ASAP7_75t_L g616 ( 
.A1(n_561),
.A2(n_297),
.B1(n_195),
.B2(n_295),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_472),
.B(n_526),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_526),
.B(n_457),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_556),
.B(n_183),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_472),
.B(n_162),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_574),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_559),
.B(n_468),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_550),
.A2(n_282),
.B1(n_162),
.B2(n_241),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_516),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_520),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_559),
.B(n_459),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_473),
.B(n_186),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_495),
.B(n_292),
.Y(n_628)
);

AOI221xp5_ASAP7_75t_L g629 ( 
.A1(n_550),
.A2(n_535),
.B1(n_465),
.B2(n_498),
.C(n_182),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_482),
.B(n_299),
.Y(n_630)
);

BUFx5_ASAP7_75t_L g631 ( 
.A(n_467),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_469),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_468),
.B(n_459),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_510),
.B(n_162),
.Y(n_634)
);

AND2x6_ASAP7_75t_SL g635 ( 
.A(n_503),
.B(n_381),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_478),
.B(n_460),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_547),
.B(n_250),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_478),
.B(n_189),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_487),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_576),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_547),
.B(n_250),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_576),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_491),
.B(n_493),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_469),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_591),
.B(n_299),
.Y(n_645)
);

BUFx5_ASAP7_75t_L g646 ( 
.A(n_467),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_586),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_591),
.B(n_302),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_568),
.B(n_197),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_585),
.B(n_302),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_464),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_520),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_488),
.A2(n_279),
.B1(n_281),
.B2(n_314),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_586),
.Y(n_654)
);

OR2x6_ASAP7_75t_L g655 ( 
.A(n_483),
.B(n_383),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_487),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_510),
.B(n_241),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_610),
.B(n_209),
.Y(n_658)
);

NOR2xp67_ASAP7_75t_L g659 ( 
.A(n_466),
.B(n_308),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_564),
.B(n_308),
.Y(n_660)
);

OR2x6_ASAP7_75t_L g661 ( 
.A(n_483),
.B(n_383),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_610),
.B(n_582),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_470),
.B(n_310),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_582),
.B(n_220),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_594),
.B(n_595),
.Y(n_665)
);

BUFx6f_ASAP7_75t_SL g666 ( 
.A(n_532),
.Y(n_666)
);

O2A1O1Ixp5_ASAP7_75t_L g667 ( 
.A1(n_594),
.A2(n_229),
.B(n_256),
.C(n_245),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_595),
.B(n_224),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_464),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_608),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_598),
.B(n_231),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_564),
.B(n_310),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_598),
.B(n_266),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_L g674 ( 
.A(n_467),
.B(n_241),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_533),
.B(n_188),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_497),
.Y(n_676)
);

AND2x6_ASAP7_75t_L g677 ( 
.A(n_523),
.B(n_241),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_466),
.B(n_284),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_514),
.B(n_241),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_475),
.A2(n_390),
.B1(n_387),
.B2(n_386),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_531),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_476),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_SL g683 ( 
.A1(n_550),
.A2(n_161),
.B1(n_164),
.B2(n_167),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_549),
.B(n_190),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_599),
.B(n_385),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_476),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_549),
.B(n_193),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_523),
.A2(n_390),
.B1(n_387),
.B2(n_386),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_589),
.B(n_385),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_497),
.B(n_70),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_599),
.B(n_204),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_549),
.B(n_213),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_514),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_481),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_612),
.B(n_233),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_589),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_608),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_523),
.A2(n_268),
.B1(n_236),
.B2(n_240),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_577),
.B(n_271),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_612),
.B(n_275),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_485),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_525),
.B(n_264),
.Y(n_702)
);

BUFx6f_ASAP7_75t_SL g703 ( 
.A(n_532),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_529),
.B(n_276),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_606),
.B(n_258),
.Y(n_705)
);

INVxp67_ASAP7_75t_SL g706 ( 
.A(n_606),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_583),
.B(n_277),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_588),
.B(n_249),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_596),
.B(n_283),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_596),
.B(n_242),
.Y(n_710)
);

O2A1O1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_566),
.A2(n_312),
.B(n_309),
.C(n_296),
.Y(n_711)
);

OAI221xp5_ASAP7_75t_L g712 ( 
.A1(n_552),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.C(n_294),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_607),
.B(n_312),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_607),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_532),
.Y(n_715)
);

NOR2xp67_ASAP7_75t_L g716 ( 
.A(n_546),
.B(n_92),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_575),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_575),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_518),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_543),
.A2(n_290),
.B1(n_235),
.B2(n_182),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_463),
.B(n_479),
.Y(n_721)
);

NOR2xp67_ASAP7_75t_SL g722 ( 
.A(n_474),
.B(n_290),
.Y(n_722)
);

NAND2xp33_ASAP7_75t_L g723 ( 
.A(n_467),
.B(n_235),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_577),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_543),
.A2(n_178),
.B1(n_169),
.B2(n_167),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_463),
.B(n_178),
.Y(n_726)
);

BUFx12f_ASAP7_75t_L g727 ( 
.A(n_539),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_551),
.B(n_169),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_524),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_555),
.B(n_164),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_479),
.B(n_161),
.Y(n_731)
);

NOR2xp67_ASAP7_75t_L g732 ( 
.A(n_565),
.B(n_136),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_544),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_539),
.B(n_9),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_467),
.B(n_132),
.Y(n_735)
);

OAI22xp33_ASAP7_75t_L g736 ( 
.A1(n_597),
.A2(n_10),
.B1(n_12),
.B2(n_18),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_501),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_486),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_489),
.B(n_127),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_504),
.B(n_126),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_513),
.B(n_539),
.Y(n_741)
);

AND2x6_ASAP7_75t_L g742 ( 
.A(n_504),
.B(n_511),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_550),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_500),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_501),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_511),
.B(n_122),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_494),
.A2(n_121),
.B1(n_119),
.B2(n_116),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_577),
.B(n_103),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_467),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_570),
.B(n_97),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_517),
.B(n_93),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_SL g752 ( 
.A(n_536),
.B(n_24),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_521),
.B(n_90),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_584),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_540),
.B(n_25),
.Y(n_755)
);

AND2x6_ASAP7_75t_L g756 ( 
.A(n_521),
.B(n_87),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_534),
.B(n_81),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_554),
.B(n_25),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_508),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_508),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_515),
.A2(n_73),
.B1(n_33),
.B2(n_34),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_507),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_534),
.B(n_30),
.Y(n_763)
);

INVx8_ASAP7_75t_L g764 ( 
.A(n_509),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_L g765 ( 
.A(n_604),
.B(n_30),
.C(n_38),
.Y(n_765)
);

O2A1O1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_609),
.A2(n_40),
.B(n_42),
.C(n_45),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_553),
.B(n_40),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_558),
.B(n_42),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_554),
.B(n_49),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_522),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_480),
.B(n_49),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_522),
.Y(n_772)
);

AOI21x1_ASAP7_75t_L g773 ( 
.A1(n_620),
.A2(n_541),
.B(n_557),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_728),
.B(n_580),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_622),
.A2(n_542),
.B(n_545),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_706),
.B(n_579),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_706),
.A2(n_542),
.B(n_545),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_617),
.A2(n_571),
.B(n_548),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_617),
.A2(n_494),
.B1(n_592),
.B2(n_573),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_643),
.B(n_560),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_618),
.A2(n_571),
.B(n_572),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_652),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_637),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_626),
.B(n_557),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_652),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_702),
.B(n_554),
.Y(n_786)
);

AOI21x1_ASAP7_75t_L g787 ( 
.A1(n_620),
.A2(n_567),
.B(n_541),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_702),
.B(n_579),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_728),
.A2(n_590),
.B(n_611),
.C(n_567),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_L g790 ( 
.A1(n_719),
.A2(n_560),
.B(n_548),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_704),
.B(n_536),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_662),
.A2(n_581),
.B(n_578),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_615),
.A2(n_494),
.B1(n_581),
.B2(n_562),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_633),
.A2(n_578),
.B(n_572),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_704),
.B(n_562),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_621),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_696),
.B(n_528),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_651),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_743),
.A2(n_614),
.B(n_624),
.C(n_705),
.Y(n_799)
);

INVx4_ASAP7_75t_L g800 ( 
.A(n_652),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_724),
.A2(n_600),
.B(n_499),
.Y(n_801)
);

O2A1O1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_743),
.A2(n_496),
.B(n_505),
.C(n_502),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_729),
.A2(n_506),
.B(n_467),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_652),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_675),
.A2(n_527),
.B(n_603),
.C(n_602),
.Y(n_805)
);

AOI21x1_ASAP7_75t_L g806 ( 
.A1(n_634),
.A2(n_502),
.B(n_505),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_733),
.B(n_492),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_696),
.B(n_563),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_762),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_639),
.B(n_519),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_754),
.A2(n_537),
.B(n_538),
.Y(n_811)
);

XOR2xp5_ASAP7_75t_L g812 ( 
.A(n_693),
.B(n_509),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_754),
.A2(n_537),
.B(n_538),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_634),
.A2(n_506),
.B(n_603),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_675),
.A2(n_506),
.B1(n_603),
.B2(n_602),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_640),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_636),
.A2(n_537),
.B(n_474),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_625),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_615),
.A2(n_527),
.B1(n_602),
.B2(n_601),
.Y(n_819)
);

NAND3xp33_ASAP7_75t_L g820 ( 
.A(n_619),
.B(n_496),
.C(n_601),
.Y(n_820)
);

NOR3xp33_ASAP7_75t_L g821 ( 
.A(n_629),
.B(n_601),
.C(n_569),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_669),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_665),
.A2(n_537),
.B(n_538),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_628),
.A2(n_527),
.B(n_492),
.C(n_569),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_682),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_628),
.A2(n_569),
.B(n_492),
.C(n_587),
.Y(n_826)
);

O2A1O1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_638),
.A2(n_506),
.B(n_53),
.C(n_54),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_642),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_686),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_641),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_647),
.B(n_506),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_715),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_SL g833 ( 
.A(n_727),
.B(n_509),
.Y(n_833)
);

AND2x2_ASAP7_75t_SL g834 ( 
.A(n_752),
.B(n_490),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_721),
.A2(n_657),
.B(n_674),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_623),
.A2(n_471),
.B1(n_477),
.B2(n_530),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_R g837 ( 
.A(n_764),
.B(n_506),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_619),
.B(n_490),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_666),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_654),
.B(n_506),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_657),
.A2(n_538),
.B(n_474),
.Y(n_841)
);

A2O1A1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_755),
.A2(n_538),
.B(n_474),
.C(n_484),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_623),
.A2(n_530),
.B1(n_471),
.B2(n_477),
.Y(n_843)
);

AO32x1_ASAP7_75t_L g844 ( 
.A1(n_613),
.A2(n_51),
.A3(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_681),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_670),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_666),
.Y(n_847)
);

O2A1O1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_697),
.A2(n_51),
.B(n_55),
.C(n_519),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_694),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_644),
.B(n_512),
.Y(n_850)
);

INVx4_ASAP7_75t_L g851 ( 
.A(n_676),
.Y(n_851)
);

A2O1A1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_755),
.A2(n_512),
.B(n_593),
.C(n_484),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_689),
.B(n_519),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_645),
.B(n_490),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_681),
.B(n_490),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_655),
.B(n_471),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_707),
.B(n_708),
.Y(n_857)
);

BUFx12f_ASAP7_75t_L g858 ( 
.A(n_655),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_749),
.A2(n_471),
.B1(n_477),
.B2(n_530),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_SL g860 ( 
.A1(n_684),
.A2(n_477),
.B(n_530),
.C(n_512),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_663),
.B(n_512),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_658),
.A2(n_605),
.B(n_709),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_684),
.A2(n_605),
.B(n_687),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_701),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_710),
.A2(n_605),
.B(n_735),
.Y(n_865)
);

AO32x1_ASAP7_75t_L g866 ( 
.A1(n_761),
.A2(n_745),
.A3(n_737),
.B1(n_760),
.B2(n_759),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_664),
.A2(n_671),
.B(n_668),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_673),
.A2(n_699),
.B(n_692),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_766),
.A2(n_726),
.B(n_731),
.C(n_763),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_749),
.A2(n_718),
.B1(n_717),
.B2(n_690),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_656),
.Y(n_871)
);

BUFx4f_ASAP7_75t_L g872 ( 
.A(n_764),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_687),
.A2(n_699),
.B(n_692),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_750),
.B(n_690),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_742),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_663),
.B(n_649),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_691),
.B(n_695),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_750),
.B(n_659),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_742),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_770),
.A2(n_772),
.B(n_700),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_656),
.B(n_716),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_742),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_732),
.B(n_685),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_650),
.B(n_713),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_744),
.A2(n_757),
.B(n_753),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_742),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_627),
.B(n_738),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_739),
.A2(n_746),
.B(n_751),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_740),
.A2(n_723),
.B(n_672),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_767),
.B(n_768),
.Y(n_890)
);

OAI21x1_ASAP7_75t_L g891 ( 
.A1(n_667),
.A2(n_679),
.B(n_747),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_660),
.A2(n_630),
.B(n_730),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_741),
.A2(n_648),
.B(n_678),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_631),
.A2(n_646),
.B(n_667),
.Y(n_894)
);

NAND3xp33_ASAP7_75t_L g895 ( 
.A(n_771),
.B(n_768),
.C(n_767),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_632),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_742),
.B(n_771),
.Y(n_897)
);

AOI21x1_ASAP7_75t_L g898 ( 
.A1(n_722),
.A2(n_661),
.B(n_655),
.Y(n_898)
);

OAI321xp33_ASAP7_75t_L g899 ( 
.A1(n_736),
.A2(n_616),
.A3(n_765),
.B1(n_712),
.B2(n_720),
.C(n_725),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_631),
.A2(n_646),
.B(n_661),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_653),
.B(n_698),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_683),
.A2(n_661),
.B1(n_756),
.B2(n_677),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_711),
.A2(n_688),
.B(n_680),
.Y(n_903)
);

NOR2x1_ASAP7_75t_SL g904 ( 
.A(n_734),
.B(n_758),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_631),
.A2(n_646),
.B(n_736),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_677),
.B(n_683),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_756),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_756),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_756),
.A2(n_677),
.B1(n_616),
.B2(n_769),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_631),
.A2(n_646),
.B(n_677),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_677),
.A2(n_756),
.B(n_646),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_764),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_635),
.B(n_703),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_L g914 ( 
.A(n_703),
.B(n_503),
.C(n_702),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_631),
.B(n_639),
.Y(n_915)
);

INVx1_ASAP7_75t_SL g916 ( 
.A(n_762),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_706),
.B(n_526),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_689),
.B(n_412),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_728),
.A2(n_622),
.B(n_704),
.C(n_702),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_706),
.B(n_526),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_SL g921 ( 
.A1(n_620),
.A2(n_634),
.B(n_657),
.C(n_748),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_724),
.A2(n_622),
.B(n_754),
.Y(n_922)
);

OAI321xp33_ASAP7_75t_L g923 ( 
.A1(n_736),
.A2(n_629),
.A3(n_616),
.B1(n_768),
.B2(n_767),
.C(n_755),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_617),
.A2(n_622),
.B(n_706),
.C(n_743),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_706),
.B(n_526),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_652),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_728),
.B(n_556),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_620),
.A2(n_617),
.B(n_622),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_622),
.A2(n_706),
.B(n_617),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_706),
.B(n_526),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_706),
.B(n_526),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_622),
.A2(n_706),
.B(n_617),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_714),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_706),
.B(n_526),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_706),
.B(n_526),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_617),
.A2(n_472),
.B1(n_615),
.B2(n_620),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_721),
.A2(n_665),
.B(n_759),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_622),
.A2(n_706),
.B(n_617),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_622),
.A2(n_706),
.B(n_617),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_728),
.B(n_556),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_SL g941 ( 
.A1(n_620),
.A2(n_634),
.B(n_657),
.C(n_748),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_706),
.A2(n_617),
.B1(n_622),
.B2(n_643),
.Y(n_942)
);

BUFx2_ASAP7_75t_L g943 ( 
.A(n_762),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_622),
.A2(n_706),
.B(n_617),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_622),
.A2(n_706),
.B(n_617),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_622),
.A2(n_706),
.B(n_617),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_SL g947 ( 
.A1(n_834),
.A2(n_895),
.B1(n_940),
.B2(n_927),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_917),
.B(n_920),
.Y(n_948)
);

AOI21xp33_ASAP7_75t_L g949 ( 
.A1(n_919),
.A2(n_774),
.B(n_890),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_916),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_923),
.B(n_857),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_785),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_929),
.A2(n_938),
.B(n_932),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_921),
.A2(n_941),
.B(n_868),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_918),
.B(n_809),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_778),
.A2(n_806),
.B(n_775),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_778),
.A2(n_775),
.B(n_781),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_912),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_796),
.Y(n_959)
);

OAI21x1_ASAP7_75t_L g960 ( 
.A1(n_781),
.A2(n_894),
.B(n_794),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_794),
.A2(n_792),
.B(n_937),
.Y(n_961)
);

AOI221xp5_ASAP7_75t_L g962 ( 
.A1(n_899),
.A2(n_901),
.B1(n_925),
.B2(n_935),
.C(n_934),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_868),
.A2(n_942),
.B(n_922),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_930),
.B(n_931),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_SL g965 ( 
.A1(n_911),
.A2(n_908),
.B(n_910),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_783),
.B(n_830),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_943),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_835),
.A2(n_780),
.B(n_873),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_832),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_912),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_835),
.A2(n_932),
.B(n_929),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_874),
.A2(n_914),
.B1(n_878),
.B2(n_877),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_876),
.B(n_938),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_856),
.B(n_851),
.Y(n_974)
);

AO31x2_ASAP7_75t_L g975 ( 
.A1(n_852),
.A2(n_805),
.A3(n_824),
.B(n_939),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_880),
.A2(n_777),
.B(n_801),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_939),
.A2(n_945),
.B(n_944),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_773),
.A2(n_787),
.B(n_885),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_944),
.A2(n_946),
.B(n_945),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_797),
.B(n_896),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_839),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_946),
.B(n_788),
.Y(n_982)
);

OAI21x1_ASAP7_75t_L g983 ( 
.A1(n_865),
.A2(n_855),
.B(n_862),
.Y(n_983)
);

AO31x2_ASAP7_75t_L g984 ( 
.A1(n_870),
.A2(n_842),
.A3(n_905),
.B(n_789),
.Y(n_984)
);

AO21x1_ASAP7_75t_L g985 ( 
.A1(n_928),
.A2(n_924),
.B(n_869),
.Y(n_985)
);

AOI221xp5_ASAP7_75t_L g986 ( 
.A1(n_936),
.A2(n_816),
.B1(n_846),
.B2(n_828),
.C(n_892),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_867),
.A2(n_883),
.B(n_861),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_853),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_884),
.B(n_776),
.Y(n_989)
);

AOI21xp33_ASAP7_75t_L g990 ( 
.A1(n_799),
.A2(n_906),
.B(n_887),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_867),
.A2(n_795),
.B(n_838),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_889),
.A2(n_905),
.B(n_784),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_897),
.A2(n_909),
.B1(n_902),
.B2(n_907),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_900),
.A2(n_840),
.B(n_831),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_785),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_863),
.A2(n_888),
.B(n_790),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_R g997 ( 
.A(n_847),
.B(n_872),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_858),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_820),
.A2(n_803),
.B(n_807),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_850),
.B(n_904),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_903),
.A2(n_893),
.B(n_854),
.C(n_891),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_SL g1002 ( 
.A1(n_908),
.A2(n_915),
.B(n_881),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_814),
.A2(n_819),
.B(n_898),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_802),
.A2(n_821),
.B(n_815),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_851),
.B(n_791),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_859),
.A2(n_843),
.B(n_836),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_860),
.A2(n_793),
.B(n_866),
.Y(n_1007)
);

AO21x2_ASAP7_75t_L g1008 ( 
.A1(n_826),
.A2(n_786),
.B(n_903),
.Y(n_1008)
);

HAxp5_ASAP7_75t_L g1009 ( 
.A(n_812),
.B(n_913),
.CON(n_1009),
.SN(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_808),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_785),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_811),
.A2(n_813),
.B(n_875),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_779),
.A2(n_933),
.B(n_827),
.C(n_879),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_866),
.A2(n_817),
.B(n_845),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_818),
.B(n_845),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_798),
.B(n_864),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_866),
.A2(n_818),
.B(n_823),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_822),
.Y(n_1018)
);

NAND2x1p5_ASAP7_75t_L g1019 ( 
.A(n_915),
.B(n_908),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_782),
.B(n_829),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_825),
.A2(n_849),
.B(n_841),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_782),
.B(n_871),
.Y(n_1022)
);

NAND3x1_ASAP7_75t_L g1023 ( 
.A(n_833),
.B(n_872),
.C(n_844),
.Y(n_1023)
);

BUFx2_ASAP7_75t_SL g1024 ( 
.A(n_912),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_882),
.A2(n_886),
.B(n_841),
.Y(n_1025)
);

OA21x2_ASAP7_75t_L g1026 ( 
.A1(n_810),
.A2(n_844),
.B(n_848),
.Y(n_1026)
);

AO31x2_ASAP7_75t_L g1027 ( 
.A1(n_800),
.A2(n_844),
.A3(n_871),
.B(n_886),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_804),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_810),
.B(n_800),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_804),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_926),
.Y(n_1031)
);

AO21x1_ASAP7_75t_L g1032 ( 
.A1(n_926),
.A2(n_890),
.B(n_942),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_SL g1033 ( 
.A1(n_837),
.A2(n_774),
.B(n_927),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_778),
.A2(n_806),
.B(n_775),
.Y(n_1034)
);

INVxp67_ASAP7_75t_SL g1035 ( 
.A(n_917),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_778),
.A2(n_806),
.B(n_775),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_919),
.A2(n_895),
.B(n_923),
.C(n_890),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_856),
.B(n_639),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_927),
.B(n_940),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_917),
.B(n_920),
.Y(n_1040)
);

AOI21xp33_ASAP7_75t_L g1041 ( 
.A1(n_927),
.A2(n_940),
.B(n_895),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_809),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_778),
.A2(n_806),
.B(n_775),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_SL g1044 ( 
.A(n_916),
.B(n_693),
.Y(n_1044)
);

AOI21xp33_ASAP7_75t_L g1045 ( 
.A1(n_927),
.A2(n_940),
.B(n_895),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_809),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_917),
.B(n_920),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_918),
.B(n_927),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_921),
.A2(n_941),
.B(n_868),
.Y(n_1049)
);

AND3x2_ASAP7_75t_L g1050 ( 
.A(n_833),
.B(n_752),
.C(n_436),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_SL g1051 ( 
.A1(n_904),
.A2(n_900),
.B(n_905),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_919),
.A2(n_920),
.B1(n_925),
.B2(n_917),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_796),
.Y(n_1053)
);

NAND2xp33_ASAP7_75t_L g1054 ( 
.A(n_919),
.B(n_917),
.Y(n_1054)
);

OAI21xp33_ASAP7_75t_L g1055 ( 
.A1(n_927),
.A2(n_412),
.B(n_728),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_919),
.A2(n_932),
.B(n_929),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_834),
.B(n_927),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_SL g1058 ( 
.A1(n_904),
.A2(n_900),
.B(n_905),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_918),
.B(n_927),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_785),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_921),
.A2(n_941),
.B(n_868),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_809),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_921),
.A2(n_941),
.B(n_868),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_921),
.A2(n_941),
.B(n_868),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_919),
.A2(n_895),
.B(n_923),
.C(n_890),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_921),
.A2(n_941),
.B(n_868),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_785),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_921),
.A2(n_941),
.B(n_868),
.Y(n_1068)
);

AO31x2_ASAP7_75t_L g1069 ( 
.A1(n_852),
.A2(n_942),
.A3(n_805),
.B(n_824),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_919),
.A2(n_895),
.B(n_923),
.C(n_890),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_917),
.B(n_920),
.Y(n_1071)
);

NOR2x1_ASAP7_75t_SL g1072 ( 
.A(n_908),
.B(n_724),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_921),
.A2(n_941),
.B(n_868),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_778),
.A2(n_806),
.B(n_775),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_921),
.A2(n_941),
.B(n_868),
.Y(n_1075)
);

AO31x2_ASAP7_75t_L g1076 ( 
.A1(n_852),
.A2(n_805),
.A3(n_824),
.B(n_942),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_778),
.A2(n_806),
.B(n_775),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_834),
.B(n_927),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_SL g1079 ( 
.A(n_916),
.B(n_693),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_917),
.B(n_920),
.Y(n_1080)
);

AOI21x1_ASAP7_75t_L g1081 ( 
.A1(n_773),
.A2(n_787),
.B(n_861),
.Y(n_1081)
);

AO31x2_ASAP7_75t_L g1082 ( 
.A1(n_852),
.A2(n_805),
.A3(n_824),
.B(n_942),
.Y(n_1082)
);

OR2x6_ASAP7_75t_L g1083 ( 
.A(n_1024),
.B(n_1002),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_951),
.A2(n_1039),
.B1(n_1055),
.B2(n_949),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_969),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1035),
.B(n_1048),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1035),
.B(n_1059),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_980),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_1029),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_974),
.B(n_1038),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_959),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_SL g1092 ( 
.A1(n_1032),
.A2(n_1058),
.B(n_1051),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1037),
.A2(n_1065),
.B1(n_1070),
.B2(n_948),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_947),
.A2(n_1057),
.B1(n_1078),
.B2(n_1041),
.Y(n_1094)
);

CKINVDCx9p33_ASAP7_75t_R g1095 ( 
.A(n_1046),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_SL g1096 ( 
.A1(n_1056),
.A2(n_953),
.B(n_1004),
.C(n_999),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_996),
.A2(n_982),
.B(n_991),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_964),
.A2(n_1040),
.B1(n_1071),
.B2(n_1047),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_947),
.B(n_955),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1053),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1016),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_989),
.B(n_1080),
.Y(n_1102)
);

INVx3_ASAP7_75t_SL g1103 ( 
.A(n_950),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_996),
.A2(n_991),
.B(n_1054),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1045),
.B(n_1038),
.Y(n_1105)
);

OR2x2_ASAP7_75t_L g1106 ( 
.A(n_1042),
.B(n_1062),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_962),
.B(n_973),
.Y(n_1107)
);

O2A1O1Ixp5_ASAP7_75t_SL g1108 ( 
.A1(n_990),
.A2(n_1052),
.B(n_993),
.C(n_1000),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_987),
.A2(n_992),
.B(n_965),
.Y(n_1109)
);

INVx3_ASAP7_75t_SL g1110 ( 
.A(n_981),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_962),
.B(n_1033),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_1029),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_1019),
.Y(n_1113)
);

AO22x1_ASAP7_75t_L g1114 ( 
.A1(n_1005),
.A2(n_974),
.B1(n_1010),
.B2(n_966),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_967),
.B(n_972),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_987),
.A2(n_992),
.B(n_968),
.Y(n_1116)
);

INVx3_ASAP7_75t_SL g1117 ( 
.A(n_958),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_986),
.A2(n_988),
.B1(n_1013),
.B2(n_1001),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1018),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_967),
.B(n_1044),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1079),
.B(n_988),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_970),
.B(n_1031),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_952),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1009),
.B(n_995),
.Y(n_1124)
);

CKINVDCx8_ASAP7_75t_R g1125 ( 
.A(n_998),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1020),
.Y(n_1126)
);

NAND2x1p5_ASAP7_75t_L g1127 ( 
.A(n_952),
.B(n_1060),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_986),
.A2(n_985),
.B1(n_1008),
.B2(n_1050),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_995),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1023),
.A2(n_968),
.B1(n_1026),
.B2(n_1007),
.Y(n_1130)
);

INVx6_ASAP7_75t_L g1131 ( 
.A(n_997),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_963),
.A2(n_954),
.B(n_1075),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_1015),
.B(n_1022),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1050),
.B(n_979),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_1011),
.B(n_1030),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1011),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_963),
.A2(n_954),
.B(n_1075),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_1028),
.B(n_1067),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1008),
.A2(n_1006),
.B1(n_1026),
.B2(n_977),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_1060),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1049),
.A2(n_1068),
.B(n_1061),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_1027),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_SL g1144 ( 
.A1(n_1061),
.A2(n_1066),
.B1(n_1073),
.B2(n_1063),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_984),
.B(n_971),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1021),
.B(n_984),
.Y(n_1146)
);

NAND3xp33_ASAP7_75t_L g1147 ( 
.A(n_1063),
.B(n_1064),
.C(n_1073),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_1027),
.Y(n_1148)
);

AO32x1_ASAP7_75t_L g1149 ( 
.A1(n_1007),
.A2(n_1014),
.A3(n_1017),
.B1(n_975),
.B2(n_984),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_984),
.B(n_971),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1064),
.A2(n_1066),
.B1(n_994),
.B2(n_1025),
.Y(n_1151)
);

NAND3xp33_ASAP7_75t_L g1152 ( 
.A(n_1025),
.B(n_1082),
.C(n_1076),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1027),
.Y(n_1153)
);

NOR2xp67_ASAP7_75t_L g1154 ( 
.A(n_1081),
.B(n_1003),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1069),
.B(n_1082),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1027),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_976),
.A2(n_957),
.B1(n_983),
.B2(n_960),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1069),
.B(n_1082),
.Y(n_1158)
);

BUFx4f_ASAP7_75t_SL g1159 ( 
.A(n_1069),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_SL g1160 ( 
.A(n_1012),
.Y(n_1160)
);

INVx4_ASAP7_75t_L g1161 ( 
.A(n_975),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_978),
.A2(n_956),
.B(n_1034),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1076),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_1036),
.B(n_1043),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1074),
.B(n_1077),
.Y(n_1165)
);

NOR2xp67_ASAP7_75t_SL g1166 ( 
.A(n_1024),
.B(n_727),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1048),
.B(n_1059),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_996),
.A2(n_982),
.B(n_991),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_996),
.A2(n_982),
.B(n_991),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1042),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_1042),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_951),
.B(n_917),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_955),
.B(n_1048),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1029),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1016),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_996),
.A2(n_982),
.B(n_991),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1016),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_974),
.B(n_1038),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_951),
.A2(n_1039),
.B1(n_895),
.B2(n_1055),
.Y(n_1179)
);

AOI21xp33_ASAP7_75t_SL g1180 ( 
.A1(n_1055),
.A2(n_412),
.B(n_774),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_996),
.A2(n_982),
.B(n_991),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_958),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_996),
.A2(n_982),
.B(n_991),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_969),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_1046),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_974),
.B(n_1038),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_996),
.A2(n_982),
.B(n_991),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1039),
.B(n_927),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1046),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_1042),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_1042),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_959),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1046),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1016),
.Y(n_1194)
);

AOI21xp33_ASAP7_75t_SL g1195 ( 
.A1(n_1055),
.A2(n_412),
.B(n_774),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_958),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_951),
.A2(n_1039),
.B1(n_895),
.B2(n_1055),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1042),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1037),
.A2(n_919),
.B(n_1065),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1037),
.A2(n_919),
.B(n_1065),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_974),
.B(n_1038),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_974),
.B(n_1038),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_959),
.Y(n_1203)
);

BUFx4_ASAP7_75t_SL g1204 ( 
.A(n_981),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_958),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_955),
.B(n_1048),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1046),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1016),
.Y(n_1208)
);

AOI221xp5_ASAP7_75t_L g1209 ( 
.A1(n_1055),
.A2(n_923),
.B1(n_951),
.B2(n_616),
.C(n_1039),
.Y(n_1209)
);

OAI21xp33_ASAP7_75t_L g1210 ( 
.A1(n_1055),
.A2(n_951),
.B(n_940),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_996),
.A2(n_982),
.B(n_991),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_996),
.A2(n_982),
.B(n_991),
.Y(n_1212)
);

NOR2xp67_ASAP7_75t_L g1213 ( 
.A(n_972),
.B(n_877),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_951),
.A2(n_917),
.B1(n_925),
.B2(n_920),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1209),
.A2(n_1188),
.B1(n_1210),
.B2(n_1084),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1163),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1210),
.A2(n_1197),
.B1(n_1179),
.B2(n_1105),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1091),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1113),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1134),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1142),
.A2(n_1109),
.B(n_1132),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1213),
.A2(n_1179),
.B1(n_1197),
.B2(n_1094),
.Y(n_1222)
);

OA21x2_ASAP7_75t_L g1223 ( 
.A1(n_1116),
.A2(n_1137),
.B(n_1104),
.Y(n_1223)
);

BUFx2_ASAP7_75t_R g1224 ( 
.A(n_1110),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1092),
.A2(n_1164),
.B(n_1165),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1213),
.A2(n_1111),
.B1(n_1200),
.B2(n_1199),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1100),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1099),
.B(n_1172),
.Y(n_1228)
);

AO21x2_ASAP7_75t_L g1229 ( 
.A1(n_1147),
.A2(n_1212),
.B(n_1169),
.Y(n_1229)
);

AO21x1_ASAP7_75t_SL g1230 ( 
.A1(n_1199),
.A2(n_1200),
.B(n_1128),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_1184),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1097),
.A2(n_1176),
.B(n_1168),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1167),
.B(n_1173),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1204),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1159),
.A2(n_1124),
.B1(n_1093),
.B2(n_1115),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_1117),
.Y(n_1236)
);

BUFx8_ASAP7_75t_SL g1237 ( 
.A(n_1085),
.Y(n_1237)
);

OAI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1180),
.A2(n_1195),
.B1(n_1086),
.B2(n_1087),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1103),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1131),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1131),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_1185),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1102),
.A2(n_1098),
.B1(n_1088),
.B2(n_1172),
.Y(n_1243)
);

OAI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1206),
.A2(n_1098),
.B1(n_1107),
.B2(n_1128),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1155),
.Y(n_1245)
);

OAI22xp33_ASAP7_75t_SL g1246 ( 
.A1(n_1093),
.A2(n_1118),
.B1(n_1083),
.B2(n_1214),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1108),
.A2(n_1214),
.B(n_1096),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_SL g1248 ( 
.A1(n_1121),
.A2(n_1120),
.B1(n_1118),
.B2(n_1083),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1164),
.A2(n_1157),
.B(n_1183),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1146),
.A2(n_1177),
.B1(n_1194),
.B2(n_1101),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1192),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1203),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1170),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1114),
.B(n_1083),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1189),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1119),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1095),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1126),
.B(n_1175),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1193),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1198),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1146),
.A2(n_1208),
.B1(n_1207),
.B2(n_1161),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1161),
.A2(n_1178),
.B1(n_1090),
.B2(n_1201),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1158),
.B(n_1136),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1181),
.A2(n_1211),
.B(n_1187),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1125),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1135),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1141),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1106),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1145),
.B(n_1150),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1090),
.A2(n_1202),
.B1(n_1201),
.B2(n_1178),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1147),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1186),
.A2(n_1202),
.B1(n_1133),
.B2(n_1152),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1152),
.B(n_1130),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1129),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1186),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_SL g1276 ( 
.A1(n_1151),
.A2(n_1130),
.B1(n_1191),
.B2(n_1190),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1143),
.B(n_1148),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1153),
.Y(n_1278)
);

OAI21xp33_ASAP7_75t_L g1279 ( 
.A1(n_1139),
.A2(n_1144),
.B(n_1166),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1156),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1149),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1089),
.A2(n_1112),
.B1(n_1174),
.B2(n_1171),
.Y(n_1282)
);

NAND2x1p5_ASAP7_75t_L g1283 ( 
.A(n_1154),
.B(n_1139),
.Y(n_1283)
);

AO21x1_ASAP7_75t_L g1284 ( 
.A1(n_1141),
.A2(n_1149),
.B(n_1127),
.Y(n_1284)
);

OAI22xp33_ASAP7_75t_SL g1285 ( 
.A1(n_1140),
.A2(n_1112),
.B1(n_1174),
.B2(n_1127),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1160),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1123),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1149),
.A2(n_1138),
.B(n_1122),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1122),
.A2(n_1196),
.B1(n_1182),
.B2(n_1205),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1083),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_1184),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1111),
.B(n_951),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1091),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1091),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1188),
.B(n_1039),
.Y(n_1295)
);

OAI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1179),
.A2(n_436),
.B1(n_752),
.B2(n_1197),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1188),
.A2(n_436),
.B1(n_752),
.B2(n_834),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1134),
.Y(n_1298)
);

NOR2xp67_ASAP7_75t_L g1299 ( 
.A(n_1088),
.B(n_851),
.Y(n_1299)
);

CKINVDCx11_ASAP7_75t_R g1300 ( 
.A(n_1110),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1213),
.A2(n_919),
.B(n_895),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1188),
.B(n_1039),
.Y(n_1302)
);

OAI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1179),
.A2(n_436),
.B1(n_752),
.B2(n_1197),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1145),
.B(n_1150),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1091),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1185),
.Y(n_1306)
);

CKINVDCx14_ASAP7_75t_R g1307 ( 
.A(n_1184),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1131),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1162),
.A2(n_961),
.B(n_976),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1103),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1091),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1188),
.A2(n_436),
.B1(n_752),
.B2(n_834),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1188),
.A2(n_436),
.B1(n_752),
.B2(n_834),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1188),
.A2(n_1084),
.B1(n_1039),
.B2(n_1179),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1209),
.A2(n_951),
.B1(n_1188),
.B2(n_895),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1228),
.B(n_1230),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1216),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1314),
.A2(n_1301),
.B(n_1215),
.Y(n_1318)
);

INVx3_ASAP7_75t_SL g1319 ( 
.A(n_1234),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1247),
.A2(n_1232),
.B(n_1221),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1295),
.B(n_1302),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1315),
.A2(n_1303),
.B(n_1296),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1266),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1290),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1228),
.B(n_1230),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1290),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1266),
.Y(n_1327)
);

NAND2x1p5_ASAP7_75t_L g1328 ( 
.A(n_1286),
.B(n_1290),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1237),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1263),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_1268),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1278),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1280),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1280),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1290),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1245),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1245),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1263),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1274),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1269),
.B(n_1304),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1222),
.A2(n_1217),
.B(n_1238),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1220),
.B(n_1298),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1274),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_R g1344 ( 
.A(n_1234),
.B(n_1231),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1292),
.B(n_1243),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1220),
.B(n_1298),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1273),
.Y(n_1347)
);

INVx4_ASAP7_75t_SL g1348 ( 
.A(n_1254),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1273),
.B(n_1277),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1271),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1288),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1233),
.B(n_1310),
.Y(n_1352)
);

INVx5_ASAP7_75t_L g1353 ( 
.A(n_1254),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1292),
.B(n_1251),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1252),
.B(n_1226),
.Y(n_1355)
);

INVx5_ASAP7_75t_L g1356 ( 
.A(n_1254),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1288),
.Y(n_1357)
);

BUFx4f_ASAP7_75t_SL g1358 ( 
.A(n_1231),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1218),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1284),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1258),
.B(n_1244),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1281),
.B(n_1261),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1242),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1227),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1283),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1281),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1284),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1258),
.B(n_1255),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1297),
.A2(n_1313),
.B(n_1312),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1229),
.B(n_1235),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1259),
.B(n_1306),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1293),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1254),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1276),
.B(n_1294),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1250),
.B(n_1256),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1317),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1340),
.B(n_1246),
.Y(n_1377)
);

INVxp67_ASAP7_75t_L g1378 ( 
.A(n_1327),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1366),
.B(n_1229),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1366),
.B(n_1229),
.Y(n_1380)
);

OAI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1318),
.A2(n_1257),
.B1(n_1311),
.B2(n_1305),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1342),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1347),
.B(n_1223),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1344),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1329),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1342),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1349),
.B(n_1357),
.Y(n_1387)
);

INVx2_ASAP7_75t_R g1388 ( 
.A(n_1357),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1322),
.A2(n_1248),
.B1(n_1279),
.B2(n_1300),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1349),
.B(n_1264),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1351),
.B(n_1249),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1348),
.B(n_1225),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1373),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1353),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1340),
.B(n_1309),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1345),
.B(n_1285),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1367),
.B(n_1267),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1348),
.B(n_1219),
.Y(n_1398)
);

AND2x4_ASAP7_75t_SL g1399 ( 
.A(n_1324),
.B(n_1272),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1360),
.B(n_1362),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1346),
.B(n_1287),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1362),
.B(n_1282),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1376),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1382),
.B(n_1330),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1389),
.A2(n_1341),
.B(n_1381),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1395),
.B(n_1316),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1382),
.B(n_1346),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1396),
.A2(n_1369),
.B1(n_1353),
.B2(n_1356),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1389),
.A2(n_1381),
.B1(n_1361),
.B2(n_1321),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1386),
.B(n_1323),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1386),
.B(n_1323),
.Y(n_1411)
);

NAND3xp33_ASAP7_75t_L g1412 ( 
.A(n_1396),
.B(n_1352),
.C(n_1375),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1397),
.B(n_1325),
.Y(n_1413)
);

NAND3xp33_ASAP7_75t_L g1414 ( 
.A(n_1377),
.B(n_1331),
.C(n_1374),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1377),
.B(n_1338),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1376),
.Y(n_1416)
);

OAI221xp5_ASAP7_75t_SL g1417 ( 
.A1(n_1400),
.A2(n_1370),
.B1(n_1374),
.B2(n_1363),
.C(n_1371),
.Y(n_1417)
);

AOI221xp5_ASAP7_75t_L g1418 ( 
.A1(n_1378),
.A2(n_1339),
.B1(n_1343),
.B2(n_1368),
.C(n_1354),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1400),
.A2(n_1257),
.B1(n_1370),
.B2(n_1262),
.Y(n_1419)
);

OAI21xp33_ASAP7_75t_L g1420 ( 
.A1(n_1400),
.A2(n_1355),
.B(n_1364),
.Y(n_1420)
);

AND2x2_ASAP7_75t_SL g1421 ( 
.A(n_1392),
.B(n_1365),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1379),
.B(n_1365),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_SL g1423 ( 
.A1(n_1399),
.A2(n_1270),
.B(n_1307),
.Y(n_1423)
);

OAI21xp5_ASAP7_75t_SL g1424 ( 
.A1(n_1399),
.A2(n_1289),
.B(n_1328),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1384),
.B(n_1358),
.Y(n_1425)
);

AOI221x1_ASAP7_75t_SL g1426 ( 
.A1(n_1401),
.A2(n_1372),
.B1(n_1299),
.B2(n_1337),
.C(n_1336),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1399),
.A2(n_1356),
.B1(n_1353),
.B2(n_1326),
.Y(n_1427)
);

OAI21xp5_ASAP7_75t_SL g1428 ( 
.A1(n_1399),
.A2(n_1328),
.B(n_1335),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1379),
.B(n_1332),
.Y(n_1429)
);

NAND3xp33_ASAP7_75t_L g1430 ( 
.A(n_1378),
.B(n_1320),
.C(n_1372),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1401),
.B(n_1402),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1380),
.B(n_1350),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1380),
.B(n_1333),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1402),
.B(n_1359),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1402),
.B(n_1359),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1391),
.B(n_1334),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1398),
.B(n_1353),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1393),
.A2(n_1356),
.B1(n_1275),
.B2(n_1348),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1431),
.B(n_1387),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1429),
.B(n_1383),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1403),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1404),
.B(n_1390),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1437),
.B(n_1392),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1403),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1421),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1416),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1416),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1406),
.B(n_1388),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1421),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1433),
.Y(n_1450)
);

INVx4_ASAP7_75t_L g1451 ( 
.A(n_1421),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1412),
.B(n_1356),
.Y(n_1452)
);

AND2x2_ASAP7_75t_SL g1453 ( 
.A(n_1438),
.B(n_1392),
.Y(n_1453)
);

AND2x4_ASAP7_75t_SL g1454 ( 
.A(n_1413),
.B(n_1398),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1436),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1404),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1432),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1434),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1435),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1405),
.A2(n_1356),
.B1(n_1393),
.B2(n_1348),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_1414),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1442),
.B(n_1410),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1461),
.B(n_1426),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1444),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1442),
.B(n_1411),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1448),
.B(n_1422),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1444),
.Y(n_1467)
);

NAND2x1p5_ASAP7_75t_L g1468 ( 
.A(n_1451),
.B(n_1394),
.Y(n_1468)
);

INVxp67_ASAP7_75t_L g1469 ( 
.A(n_1461),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1456),
.B(n_1426),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1446),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1441),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1451),
.B(n_1392),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1441),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1447),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1451),
.B(n_1392),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1440),
.B(n_1415),
.Y(n_1477)
);

AND2x4_ASAP7_75t_SL g1478 ( 
.A(n_1451),
.B(n_1398),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1440),
.B(n_1407),
.Y(n_1479)
);

NOR2x1p5_ASAP7_75t_L g1480 ( 
.A(n_1443),
.B(n_1414),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1452),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1450),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1450),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1455),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1445),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1445),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1443),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1464),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1486),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1469),
.B(n_1456),
.Y(n_1490)
);

NAND2xp33_ASAP7_75t_SL g1491 ( 
.A(n_1480),
.B(n_1449),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1464),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1469),
.B(n_1439),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1463),
.B(n_1412),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1472),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1463),
.B(n_1458),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1485),
.Y(n_1497)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1498 ( 
.A1(n_1470),
.A2(n_1405),
.B(n_1409),
.C(n_1420),
.D(n_1419),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1467),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1470),
.B(n_1458),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1486),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1487),
.B(n_1449),
.Y(n_1502)
);

INVxp67_ASAP7_75t_L g1503 ( 
.A(n_1486),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1472),
.Y(n_1504)
);

INVx2_ASAP7_75t_SL g1505 ( 
.A(n_1478),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1472),
.Y(n_1506)
);

INVxp33_ASAP7_75t_SL g1507 ( 
.A(n_1485),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1474),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1471),
.Y(n_1509)
);

OAI21xp33_ASAP7_75t_L g1510 ( 
.A1(n_1481),
.A2(n_1409),
.B(n_1417),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1482),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1481),
.A2(n_1453),
.B(n_1423),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1477),
.B(n_1459),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1482),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1487),
.B(n_1454),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1471),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1477),
.B(n_1459),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1479),
.B(n_1385),
.Y(n_1518)
);

BUFx3_ASAP7_75t_L g1519 ( 
.A(n_1468),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1475),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1462),
.B(n_1439),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1475),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1483),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1480),
.B(n_1457),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1487),
.B(n_1454),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1479),
.B(n_1457),
.Y(n_1526)
);

OAI21xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1468),
.A2(n_1408),
.B(n_1423),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1519),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1489),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1494),
.B(n_1462),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1511),
.Y(n_1531)
);

AND2x4_ASAP7_75t_SL g1532 ( 
.A(n_1501),
.B(n_1487),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_1507),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1507),
.A2(n_1453),
.B1(n_1460),
.B2(n_1468),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1496),
.B(n_1465),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1512),
.A2(n_1468),
.B(n_1474),
.Y(n_1536)
);

NOR2x1_ASAP7_75t_L g1537 ( 
.A(n_1489),
.B(n_1291),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1495),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1514),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1500),
.B(n_1465),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1510),
.B(n_1466),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1488),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1510),
.B(n_1466),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1518),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1497),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1519),
.B(n_1473),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1503),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1495),
.Y(n_1548)
);

INVx1_ASAP7_75t_SL g1549 ( 
.A(n_1491),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1505),
.B(n_1473),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1493),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1493),
.B(n_1521),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1521),
.B(n_1484),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1488),
.Y(n_1554)
);

CKINVDCx20_ASAP7_75t_R g1555 ( 
.A(n_1524),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1490),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1504),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1505),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1492),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1515),
.B(n_1525),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1504),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1515),
.B(n_1473),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1526),
.B(n_1484),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1532),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1537),
.A2(n_1533),
.B1(n_1549),
.B2(n_1555),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1529),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1542),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1542),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1532),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1554),
.Y(n_1570)
);

AOI221xp5_ASAP7_75t_L g1571 ( 
.A1(n_1533),
.A2(n_1527),
.B1(n_1498),
.B2(n_1517),
.C(n_1513),
.Y(n_1571)
);

INVxp67_ASAP7_75t_L g1572 ( 
.A(n_1537),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1549),
.B(n_1502),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1554),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1545),
.B(n_1502),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1547),
.B(n_1556),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1529),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1559),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1534),
.B(n_1551),
.Y(n_1579)
);

INVxp67_ASAP7_75t_L g1580 ( 
.A(n_1529),
.Y(n_1580)
);

OAI221xp5_ASAP7_75t_SL g1581 ( 
.A1(n_1541),
.A2(n_1498),
.B1(n_1424),
.B2(n_1420),
.C(n_1418),
.Y(n_1581)
);

OAI322xp33_ASAP7_75t_L g1582 ( 
.A1(n_1543),
.A2(n_1520),
.A3(n_1522),
.B1(n_1523),
.B2(n_1499),
.C1(n_1516),
.C2(n_1509),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1530),
.A2(n_1419),
.B1(n_1453),
.B2(n_1430),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1552),
.B(n_1492),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1544),
.A2(n_1329),
.B(n_1425),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1551),
.B(n_1466),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1559),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1552),
.B(n_1499),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1531),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1575),
.B(n_1540),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1566),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1573),
.B(n_1560),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1565),
.B(n_1535),
.Y(n_1593)
);

BUFx12f_ASAP7_75t_L g1594 ( 
.A(n_1569),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1576),
.B(n_1558),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1572),
.B(n_1573),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1571),
.B(n_1558),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1583),
.A2(n_1560),
.B1(n_1550),
.B2(n_1546),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1566),
.Y(n_1599)
);

OAI221xp5_ASAP7_75t_L g1600 ( 
.A1(n_1579),
.A2(n_1531),
.B1(n_1539),
.B2(n_1528),
.C(n_1546),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1569),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1564),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1577),
.B(n_1539),
.Y(n_1603)
);

OR2x6_ASAP7_75t_L g1604 ( 
.A(n_1585),
.B(n_1236),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1580),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1564),
.B(n_1589),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1579),
.B(n_1528),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1584),
.B(n_1560),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1595),
.B(n_1581),
.Y(n_1609)
);

AOI221xp5_ASAP7_75t_L g1610 ( 
.A1(n_1600),
.A2(n_1582),
.B1(n_1583),
.B2(n_1567),
.C(n_1587),
.Y(n_1610)
);

AOI222xp33_ASAP7_75t_L g1611 ( 
.A1(n_1593),
.A2(n_1586),
.B1(n_1574),
.B2(n_1568),
.C1(n_1578),
.C2(n_1570),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1597),
.A2(n_1588),
.B(n_1536),
.Y(n_1612)
);

OAI211xp5_ASAP7_75t_L g1613 ( 
.A1(n_1607),
.A2(n_1528),
.B(n_1536),
.C(n_1550),
.Y(n_1613)
);

OAI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1596),
.A2(n_1528),
.B(n_1560),
.Y(n_1614)
);

NAND5xp2_ASAP7_75t_L g1615 ( 
.A(n_1592),
.B(n_1562),
.C(n_1424),
.D(n_1428),
.E(n_1427),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1598),
.A2(n_1532),
.B1(n_1473),
.B2(n_1476),
.Y(n_1616)
);

AOI221xp5_ASAP7_75t_L g1617 ( 
.A1(n_1605),
.A2(n_1601),
.B1(n_1603),
.B2(n_1602),
.C(n_1599),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_R g1618 ( 
.A(n_1594),
.B(n_1239),
.Y(n_1618)
);

AOI221xp5_ASAP7_75t_L g1619 ( 
.A1(n_1602),
.A2(n_1538),
.B1(n_1561),
.B2(n_1557),
.C(n_1548),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1609),
.B(n_1606),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1616),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1617),
.Y(n_1622)
);

NAND3xp33_ASAP7_75t_SL g1623 ( 
.A(n_1611),
.B(n_1610),
.C(n_1612),
.Y(n_1623)
);

NOR2x1_ASAP7_75t_L g1624 ( 
.A(n_1614),
.B(n_1591),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1619),
.Y(n_1625)
);

OA22x2_ASAP7_75t_L g1626 ( 
.A1(n_1613),
.A2(n_1608),
.B1(n_1604),
.B2(n_1562),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1618),
.B(n_1608),
.Y(n_1627)
);

OAI21xp33_ASAP7_75t_L g1628 ( 
.A1(n_1615),
.A2(n_1590),
.B(n_1604),
.Y(n_1628)
);

NOR2x1_ASAP7_75t_L g1629 ( 
.A(n_1614),
.B(n_1604),
.Y(n_1629)
);

NAND4xp75_ASAP7_75t_L g1630 ( 
.A(n_1617),
.B(n_1548),
.C(n_1557),
.D(n_1538),
.Y(n_1630)
);

AOI221xp5_ASAP7_75t_L g1631 ( 
.A1(n_1623),
.A2(n_1548),
.B1(n_1561),
.B2(n_1557),
.C(n_1538),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1624),
.B(n_1563),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1627),
.B(n_1237),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1630),
.Y(n_1634)
);

NAND4xp75_ASAP7_75t_L g1635 ( 
.A(n_1622),
.B(n_1561),
.C(n_1522),
.D(n_1520),
.Y(n_1635)
);

AND3x4_ASAP7_75t_L g1636 ( 
.A(n_1633),
.B(n_1621),
.C(n_1629),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1634),
.B(n_1620),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1632),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1635),
.Y(n_1639)
);

INVxp67_ASAP7_75t_L g1640 ( 
.A(n_1631),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1632),
.Y(n_1641)
);

NAND3xp33_ASAP7_75t_SL g1642 ( 
.A(n_1638),
.B(n_1625),
.C(n_1628),
.Y(n_1642)
);

NAND3xp33_ASAP7_75t_SL g1643 ( 
.A(n_1636),
.B(n_1625),
.C(n_1641),
.Y(n_1643)
);

AND4x2_ASAP7_75t_L g1644 ( 
.A(n_1640),
.B(n_1626),
.C(n_1639),
.D(n_1637),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1638),
.B(n_1319),
.Y(n_1645)
);

CKINVDCx16_ASAP7_75t_R g1646 ( 
.A(n_1638),
.Y(n_1646)
);

NAND3x1_ASAP7_75t_L g1647 ( 
.A(n_1645),
.B(n_1239),
.C(n_1265),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1646),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1644),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1648),
.A2(n_1642),
.B1(n_1643),
.B2(n_1291),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1650),
.Y(n_1651)
);

AOI31xp33_ASAP7_75t_L g1652 ( 
.A1(n_1651),
.A2(n_1649),
.A3(n_1265),
.B(n_1647),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1651),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1653),
.Y(n_1654)
);

OAI21x1_ASAP7_75t_L g1655 ( 
.A1(n_1652),
.A2(n_1553),
.B(n_1563),
.Y(n_1655)
);

AOI21x1_ASAP7_75t_L g1656 ( 
.A1(n_1654),
.A2(n_1508),
.B(n_1506),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1655),
.A2(n_1553),
.B(n_1260),
.Y(n_1657)
);

NAND3xp33_ASAP7_75t_L g1658 ( 
.A(n_1657),
.B(n_1655),
.C(n_1260),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1658),
.A2(n_1656),
.B(n_1253),
.Y(n_1659)
);

OAI221xp5_ASAP7_75t_R g1660 ( 
.A1(n_1659),
.A2(n_1319),
.B1(n_1224),
.B2(n_1253),
.C(n_1308),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1660),
.A2(n_1319),
.B1(n_1240),
.B2(n_1241),
.Y(n_1661)
);


endmodule