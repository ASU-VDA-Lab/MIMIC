module fake_jpeg_8907_n_79 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_79);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_79;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVxp67_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_44),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_12),
.B1(n_28),
.B2(n_27),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_46),
.B1(n_31),
.B2(n_11),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_5),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_1),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_1),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_48),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_2),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_9),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_56),
.Y(n_66)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_57),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_39),
.B1(n_5),
.B2(n_6),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_61),
.B1(n_62),
.B2(n_24),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_4),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_7),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_8),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_58),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_52),
.Y(n_64)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_10),
.B1(n_13),
.B2(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_18),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_68),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_SL g71 ( 
.A(n_67),
.B(n_51),
.C(n_54),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_51),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_65),
.C(n_69),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_70),
.C(n_64),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_63),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_76),
.A2(n_53),
.B1(n_61),
.B2(n_66),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_25),
.Y(n_79)
);


endmodule