module real_jpeg_15021_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_0),
.A2(n_29),
.B1(n_32),
.B2(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_0),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_89),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_0),
.A2(n_68),
.B1(n_69),
.B2(n_89),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_0),
.A2(n_57),
.B1(n_63),
.B2(n_89),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_1),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_1),
.A2(n_29),
.B1(n_32),
.B2(n_81),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_1),
.A2(n_68),
.B1(n_69),
.B2(n_81),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_1),
.A2(n_57),
.B1(n_63),
.B2(n_81),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_2),
.A2(n_42),
.B1(n_68),
.B2(n_69),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_2),
.A2(n_29),
.B1(n_32),
.B2(n_42),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_2),
.A2(n_42),
.B1(n_57),
.B2(n_63),
.Y(n_126)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_5),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_5),
.A2(n_34),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_5),
.B(n_37),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_5),
.B(n_32),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_L g261 ( 
.A1(n_5),
.A2(n_68),
.B1(n_69),
.B2(n_190),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_5),
.A2(n_69),
.B(n_72),
.C(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_5),
.B(n_97),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_5),
.B(n_61),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_5),
.B(n_76),
.Y(n_288)
);

AOI21xp33_ASAP7_75t_L g297 ( 
.A1(n_5),
.A2(n_32),
.B(n_247),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_6),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_6),
.A2(n_29),
.B1(n_32),
.B2(n_79),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_6),
.A2(n_68),
.B1(n_69),
.B2(n_79),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_6),
.A2(n_57),
.B1(n_63),
.B2(n_79),
.Y(n_250)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_8),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_8),
.A2(n_29),
.B1(n_32),
.B2(n_67),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_67),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_8),
.A2(n_57),
.B1(n_63),
.B2(n_67),
.Y(n_162)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_10),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_10),
.A2(n_29),
.B1(n_32),
.B2(n_198),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_10),
.A2(n_68),
.B1(n_69),
.B2(n_198),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_10),
.A2(n_57),
.B1(n_63),
.B2(n_198),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_11),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_11),
.A2(n_29),
.B1(n_32),
.B2(n_135),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_11),
.A2(n_68),
.B1(n_69),
.B2(n_135),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_11),
.A2(n_57),
.B1(n_63),
.B2(n_135),
.Y(n_271)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_12),
.Y(n_340)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_14),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_17),
.A2(n_34),
.B1(n_35),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_17),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_17),
.A2(n_29),
.B1(n_32),
.B2(n_171),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_17),
.A2(n_68),
.B1(n_69),
.B2(n_171),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_17),
.A2(n_57),
.B1(n_63),
.B2(n_171),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_21),
.B(n_339),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_18),
.B(n_340),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_19),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_19),
.A2(n_39),
.B1(n_57),
.B2(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_19),
.A2(n_39),
.B1(n_68),
.B2(n_69),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_19),
.A2(n_29),
.B1(n_32),
.B2(n_39),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_45),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_43),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_37),
.B(n_38),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_26),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_26),
.A2(n_37),
.B1(n_196),
.B2(n_199),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_26),
.A2(n_37),
.B1(n_41),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_27),
.A2(n_28),
.B1(n_78),
.B2(n_80),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_27),
.A2(n_28),
.B1(n_80),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_27),
.A2(n_28),
.B1(n_78),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_27),
.A2(n_28),
.B1(n_101),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_27),
.A2(n_28),
.B1(n_134),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_27),
.A2(n_28),
.B1(n_197),
.B2(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_28)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_29),
.A2(n_32),
.B1(n_93),
.B2(n_94),
.Y(n_95)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_29),
.A2(n_31),
.A3(n_34),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_30),
.B(n_32),
.Y(n_188)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI32xp33_ASAP7_75t_L g245 ( 
.A1(n_32),
.A2(n_68),
.A3(n_94),
.B1(n_246),
.B2(n_248),
.Y(n_245)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_35),
.B(n_190),
.Y(n_189)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_40),
.B(n_335),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_44),
.B(n_338),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_334),
.B(n_336),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_322),
.B(n_333),
.Y(n_46)
);

AO21x1_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_149),
.B(n_319),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_136),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_112),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_50),
.B(n_112),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_82),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_51),
.B(n_98),
.C(n_110),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_55),
.B(n_77),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_52),
.A2(n_53),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_64),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_54),
.A2(n_55),
.B1(n_77),
.B2(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_54),
.A2(n_55),
.B1(n_64),
.B2(n_65),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_61),
.B(n_62),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_56),
.A2(n_61),
.B1(n_62),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_56),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_56),
.A2(n_61),
.B1(n_162),
.B2(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_56),
.A2(n_61),
.B1(n_186),
.B2(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_56),
.A2(n_61),
.B1(n_226),
.B2(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_56),
.A2(n_61),
.B1(n_250),
.B2(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_56),
.A2(n_61),
.B1(n_190),
.B2(n_283),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_56),
.A2(n_61),
.B1(n_276),
.B2(n_283),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_63),
.B1(n_72),
.B2(n_73),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_57),
.B(n_285),
.Y(n_284)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_60),
.A2(n_126),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_60),
.A2(n_160),
.B1(n_275),
.B2(n_277),
.Y(n_274)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g264 ( 
.A1(n_63),
.A2(n_73),
.B(n_190),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_66),
.A2(n_70),
.B1(n_76),
.B2(n_129),
.Y(n_128)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_69),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_69),
.B(n_93),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_75),
.B1(n_76),
.B2(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_70),
.A2(n_76),
.B(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_70),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_70),
.A2(n_76),
.B1(n_165),
.B2(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_70),
.A2(n_76),
.B1(n_214),
.B2(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_70),
.A2(n_76),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_70),
.A2(n_76),
.B1(n_262),
.B2(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_74),
.A2(n_130),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_74),
.A2(n_166),
.B1(n_241),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_98),
.B1(n_110),
.B2(n_111),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_83),
.A2(n_84),
.B(n_86),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_90),
.B1(n_96),
.B2(n_97),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_88),
.A2(n_91),
.B1(n_92),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_96),
.B1(n_97),
.B2(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_90),
.A2(n_97),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_90),
.A2(n_97),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_90),
.A2(n_97),
.B(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_91),
.A2(n_92),
.B1(n_108),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_91),
.A2(n_92),
.B1(n_132),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_91),
.A2(n_92),
.B1(n_193),
.B2(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_91),
.A2(n_92),
.B1(n_222),
.B2(n_297),
.Y(n_296)
);

NAND2x1_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_92),
.Y(n_97)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_99),
.A2(n_100),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_104),
.C(n_106),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_100),
.B(n_139),
.C(n_142),
.Y(n_323)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_109),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_104),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_109),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_104),
.B(n_145),
.C(n_147),
.Y(n_332)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.C(n_120),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_119),
.Y(n_173)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_120),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_131),
.C(n_133),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_122),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_133),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_136),
.A2(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_137),
.B(n_138),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_146),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_148),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_174),
.B(n_318),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_172),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_151),
.B(n_172),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_156),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_167),
.C(n_169),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_158),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_159),
.B(n_163),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_169),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_202),
.B(n_317),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_200),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_176),
.B(n_200),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.C(n_182),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_177),
.A2(n_178),
.B1(n_181),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_181),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_182),
.B(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_191),
.C(n_195),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_183),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_189),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_195),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_233),
.B(n_311),
.C(n_316),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_227),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_204),
.B(n_227),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_217),
.C(n_219),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_205),
.A2(n_206),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_211),
.C(n_216),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_219),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.C(n_225),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_220),
.B(n_238),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_225),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_229),
.B(n_230),
.C(n_231),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_310),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_254),
.B(n_309),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_251),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_236),
.B(n_251),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.C(n_242),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_237),
.B(n_306),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_239),
.A2(n_242),
.B1(n_243),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_239),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_249),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_244),
.A2(n_245),
.B1(n_249),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_249),
.Y(n_301)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_252),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_303),
.B(n_308),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_292),
.B(n_302),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_272),
.B(n_291),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_265),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_258),
.B(n_265),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_263),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_259),
.A2(n_260),
.B1(n_263),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_270),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_268),
.C(n_270),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_271),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_280),
.B(n_290),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_278),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_274),
.B(n_278),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_286),
.B(n_289),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_287),
.B(n_288),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_293),
.B(n_294),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_300),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_298),
.C(n_300),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_313),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_324),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_332),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_328),
.B1(n_330),
.B2(n_331),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_328),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_330),
.C(n_332),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_335),
.Y(n_338)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);


endmodule