module fake_jpeg_25064_n_25 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_25);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_25;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_9),
.Y(n_10)
);

OAI22xp5_ASAP7_75t_L g11 ( 
.A1(n_8),
.A2(n_4),
.B1(n_2),
.B2(n_1),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_10),
.B(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_16),
.C(n_13),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_1),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_12),
.B1(n_11),
.B2(n_13),
.Y(n_18)
);

INVxp33_ASAP7_75t_SL g20 ( 
.A(n_18),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_17),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_23),
.B(n_2),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_7),
.B(n_3),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_19),
.B(n_3),
.C(n_4),
.Y(n_25)
);


endmodule