module fake_jpeg_26313_n_100 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_100);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_9),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_12),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_27),
.Y(n_32)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_21),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_25),
.A2(n_16),
.B1(n_23),
.B2(n_14),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_18),
.B1(n_17),
.B2(n_24),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_23),
.B1(n_20),
.B2(n_16),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_38),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_1),
.B(n_2),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_21),
.B(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_51),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_25),
.C(n_29),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_52),
.C(n_54),
.Y(n_59)
);

AO21x1_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_28),
.B(n_15),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_47),
.B(n_49),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_27),
.B1(n_29),
.B2(n_28),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_56),
.B1(n_34),
.B2(n_30),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_29),
.B(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_2),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_64),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_54),
.B1(n_55),
.B2(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_67),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_30),
.B1(n_18),
.B2(n_17),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_30),
.B1(n_43),
.B2(n_10),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_30),
.B1(n_24),
.B2(n_3),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_4),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_68),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_75),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_53),
.C(n_44),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_65),
.C(n_61),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_64),
.B1(n_63),
.B2(n_66),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_47),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_57),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_57),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_80),
.C(n_81),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_76),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_72),
.B1(n_60),
.B2(n_77),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_71),
.B1(n_30),
.B2(n_11),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_70),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_78),
.C(n_73),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_88),
.C(n_87),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_97),
.C(n_94),
.Y(n_99)
);

AOI221xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_92),
.B1(n_8),
.B2(n_11),
.C(n_6),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_99),
.Y(n_100)
);


endmodule