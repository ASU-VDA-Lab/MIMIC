module fake_jpeg_31569_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_64),
.Y(n_65)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_39),
.B(n_18),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_2),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_0),
.B(n_1),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_0),
.B(n_1),
.Y(n_72)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_44),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_15),
.Y(n_64)
);

AND2x6_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_76),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_72),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_44),
.B1(n_52),
.B2(n_63),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_55),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_75),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_73),
.B(n_77),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_48),
.B1(n_46),
.B2(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_3),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_53),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

AO22x1_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_54),
.B1(n_49),
.B2(n_47),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_23),
.B1(n_37),
.B2(n_36),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_92),
.Y(n_99)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_2),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_89),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_91),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_48),
.C(n_22),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_96),
.C(n_102),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_21),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_101),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_20),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_104),
.A2(n_13),
.B1(n_33),
.B2(n_31),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_92),
.B(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_4),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_14),
.C(n_35),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_38),
.C(n_29),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_91),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_27),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_112),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_114),
.C(n_9),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_4),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_117),
.C(n_111),
.Y(n_120)
);

XNOR2x1_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_5),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_103),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_119),
.B(n_120),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_126),
.B1(n_110),
.B2(n_121),
.Y(n_127)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_110),
.B(n_96),
.C(n_115),
.D(n_98),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_124),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_11),
.B(n_24),
.Y(n_131)
);

AOI221xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_108),
.B1(n_9),
.B2(n_100),
.C(n_94),
.Y(n_132)
);


endmodule