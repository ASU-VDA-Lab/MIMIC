module fake_aes_2024_n_1214 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_1214);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1214;
wire n_1173;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_1198;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_1202;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_1196;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_1211;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_1175;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_1177;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_1185;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1197;
wire n_1163;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_1200;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_360;
wire n_345;
wire n_1090;
wire n_1201;
wire n_1191;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_1194;
wire n_694;
wire n_301;
wire n_1179;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1174;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1078;
wire n_1097;
wire n_572;
wire n_1017;
wire n_324;
wire n_1024;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_1169;
wire n_1204;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_1042;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_1183;
wire n_567;
wire n_809;
wire n_888;
wire n_1188;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1011;
wire n_1025;
wire n_1159;
wire n_880;
wire n_1101;
wire n_1132;
wire n_630;
wire n_1155;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_1180;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_1160;
wire n_1184;
wire n_274;
wire n_1018;
wire n_1195;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_1138;
wire n_506;
wire n_533;
wire n_490;
wire n_393;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_1171;
wire n_665;
wire n_571;
wire n_1154;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_1212;
wire n_771;
wire n_735;
wire n_696;
wire n_1091;
wire n_1203;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_1046;
wire n_460;
wire n_950;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_805;
wire n_699;
wire n_729;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_1167;
wire n_864;
wire n_1186;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_1106;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_1206;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_1178;
wire n_1209;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1210;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_875;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_1176;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_285;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_1181;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_1157;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_1199;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_363;
wire n_315;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_1170;
wire n_419;
wire n_1193;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_1125;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_1208;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_912;
wire n_620;
wire n_841;
wire n_924;
wire n_947;
wire n_1043;
wire n_1141;
wire n_378;
wire n_582;
wire n_1213;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_1189;
wire n_923;
wire n_1205;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_1172;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1007;
wire n_859;
wire n_1117;
wire n_1040;
wire n_1165;
wire n_994;
wire n_930;
wire n_1182;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_1207;
wire n_867;
wire n_1070;
wire n_1168;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_901;
wire n_834;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1164;
wire n_1038;
wire n_341;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_1104;
wire n_1187;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_1190;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_1146;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_1192;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_1166;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_1127;
wire n_269;
INVx1_ASAP7_75t_L g261 ( .A(n_99), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_228), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_201), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_184), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_29), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_178), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_129), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_174), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_246), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_46), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_195), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_170), .Y(n_272) );
INVxp67_ASAP7_75t_SL g273 ( .A(n_107), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_37), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_238), .Y(n_275) );
BUFx3_ASAP7_75t_L g276 ( .A(n_142), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_82), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_4), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_133), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_109), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_141), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_101), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_8), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_233), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_250), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_197), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_223), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_177), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_179), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_245), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_62), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_256), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_37), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_27), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_231), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_124), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_68), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_128), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_237), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_176), .Y(n_300) );
INVxp33_ASAP7_75t_L g301 ( .A(n_92), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_12), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_11), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_224), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_97), .Y(n_305) );
INVxp33_ASAP7_75t_SL g306 ( .A(n_182), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_24), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_167), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_255), .Y(n_309) );
CKINVDCx14_ASAP7_75t_R g310 ( .A(n_172), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_85), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_254), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_218), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_242), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_94), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_215), .Y(n_316) );
NOR2xp67_ASAP7_75t_L g317 ( .A(n_51), .B(n_110), .Y(n_317) );
CKINVDCx16_ASAP7_75t_R g318 ( .A(n_76), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_78), .Y(n_319) );
INVxp67_ASAP7_75t_L g320 ( .A(n_23), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_118), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_48), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_8), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_78), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_193), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_21), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_131), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_260), .Y(n_328) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_136), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_88), .Y(n_330) );
INVxp67_ASAP7_75t_L g331 ( .A(n_81), .Y(n_331) );
BUFx2_ASAP7_75t_L g332 ( .A(n_71), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_104), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_116), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_93), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_227), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_13), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_207), .Y(n_338) );
INVx1_ASAP7_75t_SL g339 ( .A(n_190), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_52), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_134), .Y(n_341) );
CKINVDCx16_ASAP7_75t_R g342 ( .A(n_158), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_150), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_77), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_196), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_257), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_157), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_50), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_9), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_2), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_241), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_60), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_66), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_236), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_206), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_36), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_181), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_185), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_56), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_90), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_200), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_243), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_70), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_41), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_27), .Y(n_365) );
INVxp67_ASAP7_75t_SL g366 ( .A(n_248), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_21), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_219), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_192), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_210), .Y(n_370) );
BUFx2_ASAP7_75t_L g371 ( .A(n_49), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_19), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_17), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_59), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_55), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_188), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_155), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_2), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_0), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_249), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_171), .Y(n_381) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_135), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_30), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_214), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_198), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_180), .Y(n_386) );
INVxp33_ASAP7_75t_SL g387 ( .A(n_162), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_117), .Y(n_388) );
CKINVDCx16_ASAP7_75t_R g389 ( .A(n_145), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_222), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_211), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_20), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_161), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_102), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_183), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_26), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_83), .Y(n_397) );
BUFx5_ASAP7_75t_L g398 ( .A(n_96), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_82), .Y(n_399) );
INVx1_ASAP7_75t_SL g400 ( .A(n_91), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_121), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_229), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_57), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_235), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_0), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_111), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_234), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_132), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_45), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_147), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_175), .Y(n_411) );
INVxp67_ASAP7_75t_L g412 ( .A(n_45), .Y(n_412) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_263), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_291), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_398), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_291), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_398), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_398), .Y(n_418) );
OAI22xp5_ASAP7_75t_SL g419 ( .A1(n_297), .A2(n_4), .B1(n_1), .B2(n_3), .Y(n_419) );
OAI22xp5_ASAP7_75t_SL g420 ( .A1(n_297), .A2(n_5), .B1(n_1), .B2(n_3), .Y(n_420) );
INVxp67_ASAP7_75t_L g421 ( .A(n_332), .Y(n_421) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_263), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_293), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_337), .B(n_5), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_398), .Y(n_425) );
CKINVDCx8_ASAP7_75t_R g426 ( .A(n_342), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_398), .Y(n_427) );
OAI22xp5_ASAP7_75t_SL g428 ( .A1(n_311), .A2(n_9), .B1(n_6), .B2(n_7), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_398), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_293), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_371), .B(n_7), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_375), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_375), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_398), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_364), .Y(n_435) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_263), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_344), .Y(n_437) );
AND2x6_ASAP7_75t_L g438 ( .A(n_276), .B(n_89), .Y(n_438) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_263), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_355), .B(n_10), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_343), .B(n_10), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_364), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_318), .A2(n_13), .B1(n_11), .B2(n_12), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_383), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_272), .B(n_14), .Y(n_445) );
AND2x2_ASAP7_75t_SL g446 ( .A(n_351), .B(n_259), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_289), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_383), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_415), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_413), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_413), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_415), .Y(n_452) );
OAI22xp33_ASAP7_75t_L g453 ( .A1(n_443), .A2(n_344), .B1(n_374), .B2(n_372), .Y(n_453) );
BUFx10_ASAP7_75t_L g454 ( .A(n_438), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_446), .B(n_389), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_417), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_417), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_421), .B(n_301), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_435), .B(n_265), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_418), .Y(n_460) );
NAND2x1p5_ASAP7_75t_L g461 ( .A(n_446), .B(n_261), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_437), .B(n_301), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_418), .Y(n_463) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_413), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_425), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_446), .A2(n_274), .B1(n_277), .B2(n_270), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_426), .B(n_264), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_442), .B(n_310), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_425), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_442), .B(n_310), .Y(n_470) );
INVx2_ASAP7_75t_SL g471 ( .A(n_438), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_427), .Y(n_472) );
INVx6_ASAP7_75t_L g473 ( .A(n_438), .Y(n_473) );
BUFx4f_ASAP7_75t_L g474 ( .A(n_438), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_427), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_429), .Y(n_476) );
BUFx3_ASAP7_75t_L g477 ( .A(n_438), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_444), .B(n_403), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_448), .B(n_278), .Y(n_479) );
INVx4_ASAP7_75t_SL g480 ( .A(n_438), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_424), .B(n_403), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_426), .B(n_264), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_413), .Y(n_483) );
INVx4_ASAP7_75t_L g484 ( .A(n_438), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_429), .Y(n_485) );
INVxp67_ASAP7_75t_SL g486 ( .A(n_431), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_448), .B(n_284), .Y(n_487) );
OR2x6_ASAP7_75t_L g488 ( .A(n_419), .B(n_283), .Y(n_488) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_441), .Y(n_489) );
NAND2xp33_ASAP7_75t_SL g490 ( .A(n_440), .B(n_275), .Y(n_490) );
INVx4_ASAP7_75t_SL g491 ( .A(n_413), .Y(n_491) );
OR2x6_ASAP7_75t_L g492 ( .A(n_419), .B(n_294), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_455), .A2(n_331), .B(n_356), .C(n_320), .Y(n_493) );
INVx2_ASAP7_75t_SL g494 ( .A(n_481), .Y(n_494) );
INVxp67_ASAP7_75t_L g495 ( .A(n_458), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_466), .A2(n_443), .B1(n_275), .B2(n_370), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_461), .A2(n_370), .B1(n_386), .B2(n_305), .Y(n_497) );
O2A1O1Ixp5_ASAP7_75t_L g498 ( .A1(n_474), .A2(n_445), .B(n_329), .C(n_366), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_461), .A2(n_386), .B1(n_305), .B2(n_420), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_457), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_489), .B(n_414), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_459), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_484), .B(n_434), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_457), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_484), .B(n_434), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_458), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_490), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_486), .B(n_288), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_460), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_468), .B(n_290), .Y(n_510) );
INVx3_ASAP7_75t_L g511 ( .A(n_484), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_468), .B(n_290), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_481), .B(n_303), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_461), .A2(n_306), .B1(n_387), .B2(n_307), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_470), .B(n_295), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_462), .A2(n_420), .B1(n_428), .B2(n_340), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_474), .B(n_262), .Y(n_517) );
INVx5_ASAP7_75t_L g518 ( .A(n_473), .Y(n_518) );
INVx3_ASAP7_75t_L g519 ( .A(n_459), .Y(n_519) );
INVx3_ASAP7_75t_L g520 ( .A(n_459), .Y(n_520) );
BUFx12f_ASAP7_75t_L g521 ( .A(n_488), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_460), .Y(n_522) );
BUFx2_ASAP7_75t_L g523 ( .A(n_470), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_477), .B(n_267), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_477), .B(n_268), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_459), .Y(n_526) );
NOR2x1p5_ASAP7_75t_L g527 ( .A(n_453), .B(n_296), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_487), .B(n_296), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_475), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_477), .B(n_269), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_479), .A2(n_319), .B1(n_322), .B2(n_302), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_467), .B(n_312), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_478), .B(n_412), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_475), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_476), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_482), .B(n_312), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_471), .A2(n_447), .B(n_338), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_479), .Y(n_538) );
NAND2x1p5_ASAP7_75t_L g539 ( .A(n_479), .B(n_323), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_488), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_449), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_452), .Y(n_542) );
OR2x6_ASAP7_75t_L g543 ( .A(n_488), .B(n_324), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_480), .B(n_416), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_480), .B(n_271), .Y(n_545) );
INVx3_ASAP7_75t_L g546 ( .A(n_454), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_492), .A2(n_365), .B1(n_326), .B2(n_349), .Y(n_547) );
INVx3_ASAP7_75t_L g548 ( .A(n_454), .Y(n_548) );
AND3x2_ASAP7_75t_SL g549 ( .A(n_488), .B(n_409), .C(n_311), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_488), .B(n_409), .Y(n_550) );
NAND3xp33_ASAP7_75t_SL g551 ( .A(n_452), .B(n_354), .C(n_346), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_473), .B(n_346), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_492), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_476), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_456), .B(n_354), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_492), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_480), .B(n_279), .Y(n_557) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_454), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_456), .Y(n_559) );
O2A1O1Ixp33_ASAP7_75t_L g560 ( .A1(n_492), .A2(n_423), .B(n_430), .C(n_416), .Y(n_560) );
INVx3_ASAP7_75t_L g561 ( .A(n_454), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_463), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_463), .A2(n_350), .B1(n_352), .B2(n_348), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_465), .B(n_360), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_492), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_469), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_469), .B(n_361), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_473), .A2(n_359), .B1(n_363), .B2(n_353), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_472), .B(n_361), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_472), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_485), .A2(n_373), .B1(n_378), .B2(n_367), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_473), .A2(n_392), .B1(n_396), .B2(n_379), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_485), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_480), .A2(n_399), .B1(n_405), .B2(n_397), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_491), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_450), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_450), .B(n_280), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_450), .B(n_281), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_451), .B(n_282), .Y(n_579) );
INVx8_ASAP7_75t_L g580 ( .A(n_543), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_539), .A2(n_376), .B1(n_369), .B2(n_273), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_519), .Y(n_582) );
BUFx2_ASAP7_75t_L g583 ( .A(n_539), .Y(n_583) );
NOR2xp33_ASAP7_75t_R g584 ( .A(n_540), .B(n_376), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_501), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_508), .B(n_266), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_501), .B(n_432), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_543), .A2(n_286), .B1(n_287), .B2(n_285), .Y(n_588) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_558), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_519), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_523), .B(n_433), .Y(n_591) );
INVx2_ASAP7_75t_SL g592 ( .A(n_513), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_506), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_495), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_520), .A2(n_292), .B1(n_299), .B2(n_298), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_520), .A2(n_300), .B1(n_308), .B2(n_304), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_497), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_526), .B(n_314), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_526), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_526), .B(n_339), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_510), .B(n_400), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_570), .Y(n_602) );
INVx2_ASAP7_75t_SL g603 ( .A(n_543), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_570), .Y(n_604) );
NOR3xp33_ASAP7_75t_SL g605 ( .A(n_553), .B(n_313), .C(n_309), .Y(n_605) );
A2O1A1Ixp33_ASAP7_75t_L g606 ( .A1(n_560), .A2(n_317), .B(n_315), .C(n_316), .Y(n_606) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_558), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_503), .A2(n_325), .B(n_321), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_550), .B(n_14), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g610 ( .A1(n_493), .A2(n_328), .B(n_330), .C(n_327), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_503), .A2(n_334), .B(n_333), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_505), .A2(n_341), .B(n_335), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_512), .B(n_345), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_573), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_L g615 ( .A1(n_515), .A2(n_357), .B(n_358), .C(n_347), .Y(n_615) );
AND2x4_ASAP7_75t_L g616 ( .A(n_543), .B(n_362), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g617 ( .A1(n_505), .A2(n_377), .B(n_368), .Y(n_617) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_558), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_502), .A2(n_381), .B1(n_384), .B2(n_380), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_544), .B(n_385), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_556), .A2(n_393), .B1(n_394), .B2(n_390), .Y(n_621) );
AND2x4_ASAP7_75t_L g622 ( .A(n_565), .B(n_395), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_538), .A2(n_402), .B1(n_404), .B2(n_401), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_573), .Y(n_624) );
AOI222xp33_ASAP7_75t_L g625 ( .A1(n_521), .A2(n_410), .B1(n_406), .B2(n_407), .C1(n_411), .C2(n_408), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_499), .Y(n_626) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_558), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_533), .B(n_276), .Y(n_628) );
INVx5_ASAP7_75t_L g629 ( .A(n_544), .Y(n_629) );
OR2x6_ASAP7_75t_SL g630 ( .A(n_507), .B(n_391), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_541), .Y(n_631) );
BUFx2_ASAP7_75t_L g632 ( .A(n_521), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_531), .B(n_15), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_537), .A2(n_483), .B(n_464), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_517), .A2(n_483), .B(n_464), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_517), .A2(n_483), .B(n_464), .Y(n_636) );
CKINVDCx8_ASAP7_75t_R g637 ( .A(n_549), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g638 ( .A1(n_563), .A2(n_382), .B(n_336), .Y(n_638) );
A2O1A1Ixp33_ASAP7_75t_L g639 ( .A1(n_542), .A2(n_382), .B(n_388), .C(n_336), .Y(n_639) );
A2O1A1Ixp33_ASAP7_75t_L g640 ( .A1(n_559), .A2(n_382), .B(n_388), .C(n_336), .Y(n_640) );
AND2x4_ASAP7_75t_L g641 ( .A(n_527), .B(n_568), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_562), .A2(n_388), .B1(n_382), .B2(n_422), .Y(n_642) );
INVx3_ASAP7_75t_L g643 ( .A(n_511), .Y(n_643) );
NOR3xp33_ASAP7_75t_SL g644 ( .A(n_551), .B(n_15), .C(n_16), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_524), .A2(n_464), .B(n_388), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_555), .B(n_422), .Y(n_646) );
XNOR2xp5_ASAP7_75t_L g647 ( .A(n_496), .B(n_16), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_566), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_524), .A2(n_530), .B(n_525), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_564), .B(n_422), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_500), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_514), .A2(n_436), .B1(n_439), .B2(n_422), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g653 ( .A1(n_498), .A2(n_436), .B(n_439), .C(n_422), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_525), .A2(n_530), .B(n_528), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_572), .A2(n_436), .B1(n_439), .B2(n_22), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_532), .B(n_18), .Y(n_656) );
NOR3xp33_ASAP7_75t_L g657 ( .A(n_516), .B(n_20), .C(n_22), .Y(n_657) );
A2O1A1Ixp33_ASAP7_75t_L g658 ( .A1(n_504), .A2(n_436), .B(n_439), .C(n_464), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_509), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_547), .B(n_23), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_571), .A2(n_574), .B1(n_569), .B2(n_567), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_536), .B(n_25), .Y(n_662) );
CKINVDCx8_ASAP7_75t_R g663 ( .A(n_549), .Y(n_663) );
A2O1A1Ixp33_ASAP7_75t_L g664 ( .A1(n_509), .A2(n_436), .B(n_439), .C(n_464), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_522), .B(n_26), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_529), .B(n_28), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_529), .B(n_28), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_552), .B(n_30), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_534), .A2(n_31), .B1(n_32), .B2(n_33), .Y(n_669) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_518), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_535), .Y(n_671) );
NOR3xp33_ASAP7_75t_SL g672 ( .A(n_577), .B(n_32), .C(n_33), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_535), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_554), .Y(n_674) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_554), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_578), .B(n_34), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_518), .B(n_35), .Y(n_677) );
O2A1O1Ixp33_ASAP7_75t_SL g678 ( .A1(n_545), .A2(n_557), .B(n_579), .C(n_575), .Y(n_678) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_518), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_518), .B(n_546), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_546), .B(n_35), .Y(n_681) );
BUFx2_ASAP7_75t_L g682 ( .A(n_548), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_548), .A2(n_36), .B1(n_38), .B2(n_39), .Y(n_683) );
CKINVDCx14_ASAP7_75t_R g684 ( .A(n_561), .Y(n_684) );
INVx3_ASAP7_75t_L g685 ( .A(n_576), .Y(n_685) );
OAI22x1_ASAP7_75t_L g686 ( .A1(n_499), .A2(n_40), .B1(n_41), .B2(n_42), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_543), .A2(n_40), .B1(n_42), .B2(n_43), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_501), .B(n_43), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_494), .B(n_44), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_501), .B(n_44), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_539), .A2(n_46), .B1(n_47), .B2(n_48), .Y(n_691) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_560), .A2(n_47), .B(n_49), .C(n_50), .Y(n_692) );
O2A1O1Ixp33_ASAP7_75t_L g693 ( .A1(n_606), .A2(n_51), .B(n_52), .C(n_53), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_688), .Y(n_694) );
OAI21xp5_ASAP7_75t_L g695 ( .A1(n_654), .A2(n_98), .B(n_95), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_597), .A2(n_54), .B1(n_55), .B2(n_56), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_591), .A2(n_54), .B1(n_57), .B2(n_58), .C(n_59), .Y(n_697) );
BUFx3_ASAP7_75t_L g698 ( .A(n_583), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_674), .Y(n_699) );
NAND2xp33_ASAP7_75t_R g700 ( .A(n_584), .B(n_58), .Y(n_700) );
OAI22x1_ASAP7_75t_L g701 ( .A1(n_687), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_592), .B(n_61), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_641), .B(n_63), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_641), .B(n_63), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_615), .A2(n_64), .B(n_65), .C(n_66), .Y(n_705) );
OAI21x1_ASAP7_75t_L g706 ( .A1(n_634), .A2(n_103), .B(n_100), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_594), .B(n_64), .Y(n_707) );
BUFx6f_ASAP7_75t_L g708 ( .A(n_589), .Y(n_708) );
AND2x4_ASAP7_75t_L g709 ( .A(n_603), .B(n_65), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_626), .A2(n_67), .B1(n_68), .B2(n_69), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_602), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_588), .A2(n_67), .B1(n_69), .B2(n_70), .Y(n_712) );
CKINVDCx5p33_ASAP7_75t_R g713 ( .A(n_637), .Y(n_713) );
NOR2xp33_ASAP7_75t_SL g714 ( .A(n_580), .B(n_663), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_585), .B(n_71), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_646), .A2(n_164), .B(n_253), .Y(n_716) );
O2A1O1Ixp33_ASAP7_75t_SL g717 ( .A1(n_653), .A2(n_163), .B(n_252), .C(n_251), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_588), .A2(n_72), .B1(n_73), .B2(n_74), .Y(n_718) );
AO32x2_ASAP7_75t_L g719 ( .A1(n_683), .A2(n_72), .A3(n_73), .B1(n_74), .B2(n_75), .Y(n_719) );
OAI221xp5_ASAP7_75t_L g720 ( .A1(n_647), .A2(n_75), .B1(n_76), .B2(n_77), .C(n_79), .Y(n_720) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_630), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_650), .A2(n_165), .B(n_247), .Y(n_722) );
NAND3xp33_ASAP7_75t_L g723 ( .A(n_605), .B(n_79), .C(n_80), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g724 ( .A1(n_656), .A2(n_80), .B(n_81), .C(n_83), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_661), .A2(n_168), .B(n_244), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g726 ( .A1(n_662), .A2(n_84), .B(n_85), .C(n_86), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_593), .A2(n_84), .B1(n_86), .B2(n_87), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g728 ( .A1(n_649), .A2(n_173), .B(n_105), .Y(n_728) );
AO31x2_ASAP7_75t_L g729 ( .A1(n_639), .A2(n_87), .A3(n_106), .B(n_108), .Y(n_729) );
OAI21xp5_ASAP7_75t_SL g730 ( .A1(n_687), .A2(n_112), .B(n_113), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_604), .Y(n_731) );
BUFx10_ASAP7_75t_L g732 ( .A(n_616), .Y(n_732) );
AOI221x1_ASAP7_75t_L g733 ( .A1(n_638), .A2(n_114), .B1(n_115), .B2(n_119), .C(n_120), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_661), .A2(n_122), .B(n_123), .Y(n_734) );
CKINVDCx5p33_ASAP7_75t_R g735 ( .A(n_632), .Y(n_735) );
OAI22xp33_ASAP7_75t_L g736 ( .A1(n_580), .A2(n_125), .B1(n_126), .B2(n_127), .Y(n_736) );
OR2x2_ASAP7_75t_L g737 ( .A(n_609), .B(n_130), .Y(n_737) );
OAI21xp5_ASAP7_75t_L g738 ( .A1(n_614), .A2(n_137), .B(n_138), .Y(n_738) );
O2A1O1Ixp5_ASAP7_75t_SL g739 ( .A1(n_669), .A2(n_139), .B(n_140), .C(n_143), .Y(n_739) );
BUFx10_ASAP7_75t_L g740 ( .A(n_616), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g741 ( .A1(n_624), .A2(n_144), .B(n_146), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_580), .A2(n_148), .B1(n_149), .B2(n_151), .Y(n_742) );
INVx3_ASAP7_75t_L g743 ( .A(n_629), .Y(n_743) );
A2O1A1Ixp33_ASAP7_75t_L g744 ( .A1(n_610), .A2(n_152), .B(n_153), .C(n_154), .Y(n_744) );
O2A1O1Ixp33_ASAP7_75t_L g745 ( .A1(n_692), .A2(n_156), .B(n_159), .C(n_160), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_651), .A2(n_166), .B(n_169), .Y(n_746) );
CKINVDCx5p33_ASAP7_75t_R g747 ( .A(n_581), .Y(n_747) );
OAI21xp5_ASAP7_75t_L g748 ( .A1(n_659), .A2(n_186), .B(n_187), .Y(n_748) );
O2A1O1Ixp33_ASAP7_75t_SL g749 ( .A1(n_681), .A2(n_189), .B(n_191), .C(n_194), .Y(n_749) );
CKINVDCx6p67_ASAP7_75t_R g750 ( .A(n_686), .Y(n_750) );
AO31x2_ASAP7_75t_L g751 ( .A1(n_640), .A2(n_199), .A3(n_202), .B(n_203), .Y(n_751) );
NOR2xp33_ASAP7_75t_SL g752 ( .A(n_638), .B(n_204), .Y(n_752) );
AND2x4_ASAP7_75t_L g753 ( .A(n_629), .B(n_258), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_690), .Y(n_754) );
INVx4_ASAP7_75t_L g755 ( .A(n_629), .Y(n_755) );
AO31x2_ASAP7_75t_L g756 ( .A1(n_658), .A2(n_205), .A3(n_208), .B(n_209), .Y(n_756) );
INVx2_ASAP7_75t_SL g757 ( .A(n_591), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_671), .A2(n_673), .B(n_613), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_660), .A2(n_212), .B1(n_213), .B2(n_216), .Y(n_759) );
A2O1A1Ixp33_ASAP7_75t_L g760 ( .A1(n_668), .A2(n_217), .B(n_220), .C(n_221), .Y(n_760) );
NAND2xp33_ASAP7_75t_L g761 ( .A(n_589), .B(n_225), .Y(n_761) );
AO31x2_ASAP7_75t_L g762 ( .A1(n_664), .A2(n_226), .A3(n_230), .B(n_232), .Y(n_762) );
INVx3_ASAP7_75t_L g763 ( .A(n_670), .Y(n_763) );
OAI21x1_ASAP7_75t_L g764 ( .A1(n_645), .A2(n_239), .B(n_240), .Y(n_764) );
A2O1A1Ixp33_ASAP7_75t_L g765 ( .A1(n_608), .A2(n_612), .B(n_611), .C(n_617), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_587), .A2(n_675), .B1(n_684), .B2(n_622), .Y(n_766) );
A2O1A1Ixp33_ASAP7_75t_L g767 ( .A1(n_631), .A2(n_648), .B(n_633), .C(n_667), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_622), .B(n_601), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_582), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_689), .B(n_625), .Y(n_770) );
CKINVDCx8_ASAP7_75t_R g771 ( .A(n_670), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g772 ( .A(n_644), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_590), .Y(n_773) );
INVx2_ASAP7_75t_L g774 ( .A(n_599), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_621), .A2(n_598), .B1(n_600), .B2(n_628), .Y(n_775) );
OAI22xp33_ASAP7_75t_L g776 ( .A1(n_676), .A2(n_691), .B1(n_596), .B2(n_595), .Y(n_776) );
O2A1O1Ixp33_ASAP7_75t_L g777 ( .A1(n_619), .A2(n_623), .B(n_657), .C(n_625), .Y(n_777) );
CKINVDCx16_ASAP7_75t_R g778 ( .A(n_666), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_685), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g780 ( .A1(n_665), .A2(n_643), .B(n_652), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_586), .B(n_620), .Y(n_781) );
OAI21x1_ASAP7_75t_L g782 ( .A1(n_677), .A2(n_680), .B(n_685), .Y(n_782) );
BUFx6f_ASAP7_75t_L g783 ( .A(n_607), .Y(n_783) );
AO31x2_ASAP7_75t_L g784 ( .A1(n_655), .A2(n_682), .A3(n_672), .B(n_678), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_670), .B(n_679), .Y(n_785) );
INVxp67_ASAP7_75t_L g786 ( .A(n_642), .Y(n_786) );
INVxp67_ASAP7_75t_L g787 ( .A(n_679), .Y(n_787) );
CKINVDCx16_ASAP7_75t_R g788 ( .A(n_679), .Y(n_788) );
NAND2x1p5_ASAP7_75t_L g789 ( .A(n_607), .B(n_618), .Y(n_789) );
OR2x6_ASAP7_75t_L g790 ( .A(n_607), .B(n_618), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_618), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g792 ( .A1(n_627), .A2(n_474), .B(n_484), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_627), .B(n_540), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_627), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_588), .A2(n_461), .B1(n_466), .B2(n_539), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_626), .A2(n_521), .B1(n_461), .B2(n_455), .Y(n_796) );
A2O1A1Ixp33_ASAP7_75t_L g797 ( .A1(n_615), .A2(n_662), .B(n_656), .C(n_654), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_688), .Y(n_798) );
AO32x2_ASAP7_75t_L g799 ( .A1(n_683), .A2(n_669), .A3(n_652), .B1(n_596), .B2(n_595), .Y(n_799) );
OAI21x1_ASAP7_75t_L g800 ( .A1(n_634), .A2(n_636), .B(n_635), .Y(n_800) );
BUFx3_ASAP7_75t_L g801 ( .A(n_583), .Y(n_801) );
AND2x4_ASAP7_75t_L g802 ( .A(n_583), .B(n_603), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_688), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_674), .Y(n_804) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_583), .Y(n_805) );
A2O1A1Ixp33_ASAP7_75t_L g806 ( .A1(n_615), .A2(n_662), .B(n_656), .C(n_654), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_588), .A2(n_461), .B1(n_466), .B2(n_539), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_588), .A2(n_461), .B1(n_466), .B2(n_539), .Y(n_808) );
CKINVDCx5p33_ASAP7_75t_R g809 ( .A(n_584), .Y(n_809) );
OAI22xp33_ASAP7_75t_L g810 ( .A1(n_580), .A2(n_497), .B1(n_499), .B2(n_461), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_592), .B(n_540), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_592), .B(n_540), .Y(n_812) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_589), .Y(n_813) );
AO21x2_ASAP7_75t_L g814 ( .A1(n_653), .A2(n_640), .B(n_639), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_688), .Y(n_815) );
BUFx12f_ASAP7_75t_L g816 ( .A(n_632), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_592), .B(n_540), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g818 ( .A(n_816), .Y(n_818) );
BUFx2_ASAP7_75t_L g819 ( .A(n_698), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_770), .A2(n_807), .B1(n_808), .B2(n_795), .Y(n_820) );
OR2x2_ASAP7_75t_L g821 ( .A(n_805), .B(n_801), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_778), .A2(n_737), .B1(n_750), .B2(n_709), .Y(n_822) );
INVxp67_ASAP7_75t_L g823 ( .A(n_707), .Y(n_823) );
AOI21xp5_ASAP7_75t_L g824 ( .A1(n_797), .A2(n_806), .B(n_767), .Y(n_824) );
OA21x2_ASAP7_75t_L g825 ( .A1(n_733), .A2(n_695), .B(n_725), .Y(n_825) );
OAI21xp5_ASAP7_75t_L g826 ( .A1(n_758), .A2(n_765), .B(n_734), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_694), .B(n_754), .Y(n_827) );
NOR3xp33_ASAP7_75t_L g828 ( .A(n_720), .B(n_777), .C(n_723), .Y(n_828) );
BUFx3_ASAP7_75t_L g829 ( .A(n_771), .Y(n_829) );
OA21x2_ASAP7_75t_L g830 ( .A1(n_706), .A2(n_728), .B(n_780), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_711), .Y(n_831) );
NOR2x1_ASAP7_75t_R g832 ( .A(n_721), .B(n_809), .Y(n_832) );
AOI21xp33_ASAP7_75t_L g833 ( .A1(n_745), .A2(n_776), .B(n_775), .Y(n_833) );
OR2x2_ASAP7_75t_L g834 ( .A(n_757), .B(n_699), .Y(n_834) );
INVx1_ASAP7_75t_SL g835 ( .A(n_732), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_731), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_798), .B(n_803), .Y(n_837) );
INVx4_ASAP7_75t_L g838 ( .A(n_788), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_815), .B(n_768), .Y(n_839) );
BUFx4f_ASAP7_75t_SL g840 ( .A(n_732), .Y(n_840) );
AOI21xp5_ASAP7_75t_L g841 ( .A1(n_717), .A2(n_792), .B(n_752), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_810), .B(n_766), .Y(n_842) );
OA21x2_ASAP7_75t_L g843 ( .A1(n_748), .A2(n_741), .B(n_738), .Y(n_843) );
INVx3_ASAP7_75t_L g844 ( .A(n_755), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_804), .Y(n_845) );
BUFx4f_ASAP7_75t_L g846 ( .A(n_802), .Y(n_846) );
OAI21xp5_ASAP7_75t_L g847 ( .A1(n_739), .A2(n_786), .B(n_715), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_802), .B(n_747), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_703), .B(n_704), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_701), .Y(n_850) );
AOI21xp33_ASAP7_75t_L g851 ( .A1(n_693), .A2(n_730), .B(n_814), .Y(n_851) );
OAI21xp5_ASAP7_75t_L g852 ( .A1(n_744), .A2(n_705), .B(n_724), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_796), .B(n_774), .Y(n_853) );
OA21x2_ASAP7_75t_L g854 ( .A1(n_764), .A2(n_760), .B(n_746), .Y(n_854) );
CKINVDCx5p33_ASAP7_75t_R g855 ( .A(n_700), .Y(n_855) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_735), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_769), .B(n_773), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_719), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_781), .B(n_779), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_791), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_719), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_712), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_718), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_702), .A2(n_772), .B1(n_811), .B2(n_812), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_817), .A2(n_710), .B1(n_697), .B2(n_793), .Y(n_865) );
OAI21xp5_ASAP7_75t_L g866 ( .A1(n_726), .A2(n_716), .B(n_722), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_740), .B(n_696), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_740), .B(n_784), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_714), .A2(n_727), .B1(n_713), .B2(n_755), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_784), .B(n_785), .Y(n_870) );
OAI21x1_ASAP7_75t_SL g871 ( .A1(n_742), .A2(n_759), .B(n_794), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_743), .B(n_787), .Y(n_872) );
OR2x6_ASAP7_75t_L g873 ( .A(n_753), .B(n_790), .Y(n_873) );
AO221x2_ASAP7_75t_L g874 ( .A1(n_736), .A2(n_799), .B1(n_729), .B2(n_784), .C(n_756), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_743), .Y(n_875) );
AO21x2_ASAP7_75t_L g876 ( .A1(n_814), .A2(n_761), .B(n_749), .Y(n_876) );
BUFx3_ASAP7_75t_L g877 ( .A(n_763), .Y(n_877) );
AOI21xp5_ASAP7_75t_L g878 ( .A1(n_789), .A2(n_708), .B(n_783), .Y(n_878) );
AOI21xp5_ASAP7_75t_L g879 ( .A1(n_813), .A2(n_799), .B(n_756), .Y(n_879) );
AOI21xp5_ASAP7_75t_L g880 ( .A1(n_756), .A2(n_762), .B(n_751), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_751), .B(n_762), .Y(n_881) );
AND2x2_ASAP7_75t_L g882 ( .A(n_770), .B(n_494), .Y(n_882) );
CKINVDCx5p33_ASAP7_75t_R g883 ( .A(n_816), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_709), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_770), .B(n_494), .Y(n_885) );
OAI21xp5_ASAP7_75t_L g886 ( .A1(n_767), .A2(n_758), .B(n_797), .Y(n_886) );
AOI21xp5_ASAP7_75t_L g887 ( .A1(n_797), .A2(n_806), .B(n_767), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_770), .B(n_494), .Y(n_888) );
INVx3_ASAP7_75t_L g889 ( .A(n_771), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_770), .B(n_494), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_711), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_709), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_709), .Y(n_893) );
AOI21xp5_ASAP7_75t_L g894 ( .A1(n_797), .A2(n_806), .B(n_767), .Y(n_894) );
OA21x2_ASAP7_75t_L g895 ( .A1(n_800), .A2(n_782), .B(n_733), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_711), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_709), .Y(n_897) );
AOI21xp5_ASAP7_75t_L g898 ( .A1(n_797), .A2(n_806), .B(n_767), .Y(n_898) );
AOI21xp5_ASAP7_75t_L g899 ( .A1(n_797), .A2(n_806), .B(n_767), .Y(n_899) );
CKINVDCx20_ASAP7_75t_R g900 ( .A(n_809), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_770), .B(n_494), .Y(n_901) );
INVx5_ASAP7_75t_SL g902 ( .A(n_790), .Y(n_902) );
AOI21xp5_ASAP7_75t_L g903 ( .A1(n_797), .A2(n_806), .B(n_767), .Y(n_903) );
INVx3_ASAP7_75t_L g904 ( .A(n_771), .Y(n_904) );
AOI21xp5_ASAP7_75t_L g905 ( .A1(n_797), .A2(n_806), .B(n_767), .Y(n_905) );
INVxp67_ASAP7_75t_L g906 ( .A(n_805), .Y(n_906) );
AOI21xp5_ASAP7_75t_L g907 ( .A1(n_797), .A2(n_806), .B(n_767), .Y(n_907) );
AND2x4_ASAP7_75t_L g908 ( .A(n_802), .B(n_583), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_694), .B(n_754), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_694), .B(n_754), .Y(n_910) );
AOI22xp5_ASAP7_75t_L g911 ( .A1(n_770), .A2(n_626), .B1(n_597), .B2(n_494), .Y(n_911) );
AOI21xp5_ASAP7_75t_L g912 ( .A1(n_797), .A2(n_806), .B(n_767), .Y(n_912) );
AOI21xp33_ASAP7_75t_SL g913 ( .A1(n_700), .A2(n_772), .B(n_721), .Y(n_913) );
INVxp67_ASAP7_75t_L g914 ( .A(n_805), .Y(n_914) );
A2O1A1Ixp33_ASAP7_75t_L g915 ( .A1(n_797), .A2(n_806), .B(n_777), .C(n_730), .Y(n_915) );
OR2x2_ASAP7_75t_L g916 ( .A(n_805), .B(n_494), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_709), .Y(n_917) );
HB1xp67_ASAP7_75t_L g918 ( .A(n_788), .Y(n_918) );
OR2x2_ASAP7_75t_L g919 ( .A(n_805), .B(n_494), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_709), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_694), .B(n_754), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_795), .A2(n_461), .B1(n_808), .B2(n_807), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_709), .Y(n_923) );
AO21x2_ASAP7_75t_L g924 ( .A1(n_780), .A2(n_734), .B(n_725), .Y(n_924) );
INVx4_ASAP7_75t_SL g925 ( .A(n_753), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_858), .Y(n_926) );
OAI21xp5_ASAP7_75t_L g927 ( .A1(n_828), .A2(n_833), .B(n_915), .Y(n_927) );
AO21x2_ASAP7_75t_L g928 ( .A1(n_880), .A2(n_881), .B(n_879), .Y(n_928) );
OR2x2_ASAP7_75t_L g929 ( .A(n_890), .B(n_882), .Y(n_929) );
INVx2_ASAP7_75t_SL g930 ( .A(n_846), .Y(n_930) );
OAI22xp5_ASAP7_75t_SL g931 ( .A1(n_855), .A2(n_822), .B1(n_840), .B2(n_911), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_885), .B(n_888), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_849), .A2(n_922), .B1(n_842), .B2(n_901), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_831), .B(n_836), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_891), .B(n_896), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_861), .Y(n_936) );
AO21x2_ASAP7_75t_L g937 ( .A1(n_824), .A2(n_899), .B(n_907), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_857), .Y(n_938) );
HB1xp67_ASAP7_75t_L g939 ( .A(n_918), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_857), .Y(n_940) );
OA21x2_ASAP7_75t_L g941 ( .A1(n_887), .A2(n_903), .B(n_905), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_839), .B(n_827), .Y(n_942) );
AND2x4_ASAP7_75t_L g943 ( .A(n_925), .B(n_873), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_839), .B(n_827), .Y(n_944) );
OAI31xp33_ASAP7_75t_L g945 ( .A1(n_822), .A2(n_922), .A3(n_862), .B(n_863), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_870), .Y(n_946) );
OAI322xp33_ASAP7_75t_L g947 ( .A1(n_850), .A2(n_823), .A3(n_894), .B1(n_898), .B2(n_912), .C1(n_910), .C2(n_837), .Y(n_947) );
OR2x2_ASAP7_75t_L g948 ( .A(n_820), .B(n_837), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_870), .Y(n_949) );
BUFx3_ASAP7_75t_L g950 ( .A(n_829), .Y(n_950) );
AND2x4_ASAP7_75t_L g951 ( .A(n_925), .B(n_873), .Y(n_951) );
BUFx3_ASAP7_75t_L g952 ( .A(n_819), .Y(n_952) );
NOR2x1_ASAP7_75t_SL g953 ( .A(n_873), .B(n_925), .Y(n_953) );
AO21x2_ASAP7_75t_L g954 ( .A1(n_886), .A2(n_826), .B(n_851), .Y(n_954) );
NOR2xp33_ASAP7_75t_L g955 ( .A(n_856), .B(n_867), .Y(n_955) );
INVx2_ASAP7_75t_L g956 ( .A(n_860), .Y(n_956) );
INVx2_ASAP7_75t_SL g957 ( .A(n_846), .Y(n_957) );
INVx2_ASAP7_75t_L g958 ( .A(n_895), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_909), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_909), .B(n_910), .Y(n_960) );
AND2x4_ASAP7_75t_SL g961 ( .A(n_838), .B(n_908), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_921), .B(n_845), .Y(n_962) );
INVx4_ASAP7_75t_L g963 ( .A(n_889), .Y(n_963) );
HB1xp67_ASAP7_75t_L g964 ( .A(n_821), .Y(n_964) );
AO21x2_ASAP7_75t_L g965 ( .A1(n_833), .A2(n_847), .B(n_868), .Y(n_965) );
NOR2xp33_ASAP7_75t_L g966 ( .A(n_848), .B(n_838), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_859), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_859), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_874), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_865), .B(n_919), .Y(n_970) );
AO21x2_ASAP7_75t_L g971 ( .A1(n_841), .A2(n_852), .B(n_924), .Y(n_971) );
AOI21xp5_ASAP7_75t_SL g972 ( .A1(n_874), .A2(n_843), .B(n_830), .Y(n_972) );
AOI22xp5_ASAP7_75t_L g973 ( .A1(n_853), .A2(n_897), .B1(n_923), .B2(n_893), .Y(n_973) );
AOI22xp33_ASAP7_75t_SL g974 ( .A1(n_902), .A2(n_889), .B1(n_904), .B2(n_852), .Y(n_974) );
INVxp33_ASAP7_75t_L g975 ( .A(n_832), .Y(n_975) );
AOI221xp5_ASAP7_75t_L g976 ( .A1(n_913), .A2(n_864), .B1(n_906), .B2(n_914), .C(n_884), .Y(n_976) );
INVx3_ASAP7_75t_L g977 ( .A(n_844), .Y(n_977) );
NOR2xp33_ASAP7_75t_SL g978 ( .A(n_818), .B(n_883), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_892), .B(n_917), .Y(n_979) );
AO21x2_ASAP7_75t_L g980 ( .A1(n_924), .A2(n_876), .B(n_871), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_916), .B(n_920), .Y(n_981) );
INVx4_ASAP7_75t_L g982 ( .A(n_904), .Y(n_982) );
AOI21xp5_ASAP7_75t_SL g983 ( .A1(n_843), .A2(n_830), .B(n_825), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_853), .Y(n_984) );
INVx3_ASAP7_75t_L g985 ( .A(n_844), .Y(n_985) );
OR2x6_ASAP7_75t_L g986 ( .A(n_878), .B(n_875), .Y(n_986) );
AO21x2_ASAP7_75t_L g987 ( .A1(n_876), .A2(n_866), .B(n_825), .Y(n_987) );
HB1xp67_ASAP7_75t_L g988 ( .A(n_834), .Y(n_988) );
BUFx2_ASAP7_75t_L g989 ( .A(n_872), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_877), .B(n_902), .Y(n_990) );
BUFx2_ASAP7_75t_L g991 ( .A(n_835), .Y(n_991) );
OA21x2_ASAP7_75t_L g992 ( .A1(n_854), .A2(n_869), .B(n_835), .Y(n_992) );
OAI21xp5_ASAP7_75t_L g993 ( .A1(n_854), .A2(n_900), .B(n_902), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_858), .Y(n_994) );
HB1xp67_ASAP7_75t_L g995 ( .A(n_918), .Y(n_995) );
AO21x2_ASAP7_75t_L g996 ( .A1(n_880), .A2(n_881), .B(n_879), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_858), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_858), .Y(n_998) );
OAI31xp33_ASAP7_75t_L g999 ( .A1(n_822), .A2(n_720), .A3(n_810), .B(n_527), .Y(n_999) );
OR2x6_ASAP7_75t_L g1000 ( .A(n_873), .B(n_922), .Y(n_1000) );
OR2x2_ASAP7_75t_L g1001 ( .A(n_969), .B(n_948), .Y(n_1001) );
HB1xp67_ASAP7_75t_L g1002 ( .A(n_964), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_926), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_999), .A2(n_1000), .B1(n_933), .B2(n_945), .Y(n_1004) );
OR2x2_ASAP7_75t_L g1005 ( .A(n_969), .B(n_948), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_960), .B(n_962), .Y(n_1006) );
OR2x6_ASAP7_75t_L g1007 ( .A(n_1000), .B(n_943), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_946), .B(n_949), .Y(n_1008) );
AND2x4_ASAP7_75t_L g1009 ( .A(n_1000), .B(n_946), .Y(n_1009) );
AOI31xp33_ASAP7_75t_L g1010 ( .A1(n_974), .A2(n_943), .A3(n_951), .B(n_993), .Y(n_1010) );
OR2x2_ASAP7_75t_L g1011 ( .A(n_949), .B(n_929), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_936), .B(n_994), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_936), .B(n_994), .Y(n_1013) );
BUFx3_ASAP7_75t_L g1014 ( .A(n_952), .Y(n_1014) );
OR2x2_ASAP7_75t_L g1015 ( .A(n_929), .B(n_984), .Y(n_1015) );
HB1xp67_ASAP7_75t_L g1016 ( .A(n_952), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_997), .B(n_998), .Y(n_1017) );
NOR2x1_ASAP7_75t_L g1018 ( .A(n_943), .B(n_951), .Y(n_1018) );
NOR2xp33_ASAP7_75t_L g1019 ( .A(n_931), .B(n_932), .Y(n_1019) );
AND2x4_ASAP7_75t_L g1020 ( .A(n_1000), .B(n_986), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_984), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_1000), .B(n_934), .Y(n_1022) );
NOR2xp33_ASAP7_75t_L g1023 ( .A(n_966), .B(n_955), .Y(n_1023) );
OR2x2_ASAP7_75t_L g1024 ( .A(n_989), .B(n_959), .Y(n_1024) );
BUFx3_ASAP7_75t_L g1025 ( .A(n_951), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_934), .B(n_935), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_938), .B(n_940), .Y(n_1027) );
AOI21xp5_ASAP7_75t_L g1028 ( .A1(n_927), .A2(n_947), .B(n_983), .Y(n_1028) );
AOI222xp33_ASAP7_75t_L g1029 ( .A1(n_970), .A2(n_944), .B1(n_942), .B2(n_967), .C1(n_968), .C2(n_976), .Y(n_1029) );
HB1xp67_ASAP7_75t_L g1030 ( .A(n_989), .Y(n_1030) );
INVx2_ASAP7_75t_L g1031 ( .A(n_958), .Y(n_1031) );
INVxp33_ASAP7_75t_L g1032 ( .A(n_978), .Y(n_1032) );
INVx2_ASAP7_75t_SL g1033 ( .A(n_991), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_967), .A2(n_968), .B1(n_995), .B2(n_939), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_956), .B(n_937), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_937), .B(n_979), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_937), .B(n_979), .Y(n_1037) );
AND2x4_ASAP7_75t_L g1038 ( .A(n_986), .B(n_953), .Y(n_1038) );
NOR2x1_ASAP7_75t_L g1039 ( .A(n_977), .B(n_985), .Y(n_1039) );
INVxp67_ASAP7_75t_SL g1040 ( .A(n_953), .Y(n_1040) );
NOR2x1_ASAP7_75t_SL g1041 ( .A(n_986), .B(n_963), .Y(n_1041) );
HB1xp67_ASAP7_75t_L g1042 ( .A(n_988), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_954), .B(n_941), .Y(n_1043) );
OR2x2_ASAP7_75t_L g1044 ( .A(n_991), .B(n_954), .Y(n_1044) );
NOR2xp33_ASAP7_75t_R g1045 ( .A(n_930), .B(n_957), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1003), .Y(n_1046) );
HB1xp67_ASAP7_75t_L g1047 ( .A(n_1030), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1003), .Y(n_1048) );
AND2x2_ASAP7_75t_SL g1049 ( .A(n_1020), .B(n_992), .Y(n_1049) );
BUFx3_ASAP7_75t_L g1050 ( .A(n_1014), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_1008), .B(n_973), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_1036), .B(n_996), .Y(n_1052) );
INVxp67_ASAP7_75t_L g1053 ( .A(n_1016), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1036), .B(n_996), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_1037), .B(n_996), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_1037), .B(n_928), .Y(n_1056) );
INVx1_ASAP7_75t_SL g1057 ( .A(n_1014), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_1035), .B(n_928), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_1006), .B(n_928), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_1006), .B(n_965), .Y(n_1060) );
AND2x4_ASAP7_75t_L g1061 ( .A(n_1020), .B(n_980), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_1008), .B(n_973), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_1012), .B(n_965), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1012), .B(n_965), .Y(n_1064) );
OR2x2_ASAP7_75t_L g1065 ( .A(n_1001), .B(n_992), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_1013), .B(n_971), .Y(n_1066) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_1004), .A2(n_977), .B1(n_985), .B2(n_930), .Y(n_1067) );
BUFx3_ASAP7_75t_L g1068 ( .A(n_1014), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_1035), .B(n_971), .Y(n_1069) );
INVx2_ASAP7_75t_L g1070 ( .A(n_1031), .Y(n_1070) );
BUFx2_ASAP7_75t_L g1071 ( .A(n_1038), .Y(n_1071) );
OR2x2_ASAP7_75t_L g1072 ( .A(n_1005), .B(n_941), .Y(n_1072) );
NAND2x1_ASAP7_75t_SL g1073 ( .A(n_1038), .B(n_985), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1074 ( .A(n_1027), .B(n_941), .Y(n_1074) );
INVx2_ASAP7_75t_SL g1075 ( .A(n_1038), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1017), .B(n_980), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1017), .B(n_980), .Y(n_1077) );
OR2x2_ASAP7_75t_L g1078 ( .A(n_1011), .B(n_987), .Y(n_1078) );
NOR2xp33_ASAP7_75t_L g1079 ( .A(n_1019), .B(n_963), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_1021), .B(n_972), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1059), .B(n_1009), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1059), .B(n_1009), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1046), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1046), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g1085 ( .A(n_1047), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1048), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1048), .Y(n_1087) );
INVx3_ASAP7_75t_L g1088 ( .A(n_1071), .Y(n_1088) );
INVx2_ASAP7_75t_L g1089 ( .A(n_1070), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1060), .B(n_1029), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_1053), .B(n_1029), .Y(n_1091) );
OR2x6_ASAP7_75t_L g1092 ( .A(n_1071), .B(n_1007), .Y(n_1092) );
NOR2x1_ASAP7_75t_L g1093 ( .A(n_1050), .B(n_1010), .Y(n_1093) );
AND2x4_ASAP7_75t_SL g1094 ( .A(n_1075), .B(n_1038), .Y(n_1094) );
HB1xp67_ASAP7_75t_L g1095 ( .A(n_1047), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_1052), .B(n_1009), .Y(n_1096) );
OR2x2_ASAP7_75t_L g1097 ( .A(n_1078), .B(n_1044), .Y(n_1097) );
AND2x4_ASAP7_75t_L g1098 ( .A(n_1075), .B(n_1061), .Y(n_1098) );
NAND2xp5_ASAP7_75t_SL g1099 ( .A(n_1057), .B(n_1010), .Y(n_1099) );
INVx1_ASAP7_75t_SL g1100 ( .A(n_1057), .Y(n_1100) );
AND2x2_ASAP7_75t_SL g1101 ( .A(n_1049), .B(n_1020), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1052), .B(n_1009), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1103 ( .A(n_1053), .B(n_1002), .Y(n_1103) );
OAI211xp5_ASAP7_75t_L g1104 ( .A1(n_1079), .A2(n_1045), .B(n_1034), .C(n_1023), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1054), .B(n_1022), .Y(n_1105) );
AND2x4_ASAP7_75t_SL g1106 ( .A(n_1075), .B(n_1007), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1054), .B(n_1043), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1055), .B(n_1043), .Y(n_1108) );
OAI22xp33_ASAP7_75t_L g1109 ( .A1(n_1067), .A2(n_1007), .B1(n_1040), .B2(n_1032), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1110 ( .A(n_1051), .B(n_1042), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1051), .B(n_1026), .Y(n_1111) );
NOR2xp33_ASAP7_75t_L g1112 ( .A(n_1079), .B(n_975), .Y(n_1112) );
AND2x4_ASAP7_75t_L g1113 ( .A(n_1061), .B(n_1007), .Y(n_1113) );
OR2x2_ASAP7_75t_L g1114 ( .A(n_1097), .B(n_1072), .Y(n_1114) );
INVxp67_ASAP7_75t_L g1115 ( .A(n_1085), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1107), .B(n_1055), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1117 ( .A(n_1097), .B(n_1072), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_1090), .B(n_1063), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1091), .B(n_1063), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1107), .B(n_1056), .Y(n_1120) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1089), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1083), .Y(n_1122) );
OAI211xp5_ASAP7_75t_L g1123 ( .A1(n_1093), .A2(n_1104), .B(n_1099), .C(n_1112), .Y(n_1123) );
NAND2x1p5_ASAP7_75t_L g1124 ( .A(n_1101), .B(n_1050), .Y(n_1124) );
NAND2x1p5_ASAP7_75t_L g1125 ( .A(n_1101), .B(n_1050), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_1108), .B(n_1064), .Y(n_1126) );
INVxp67_ASAP7_75t_L g1127 ( .A(n_1095), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1083), .Y(n_1128) );
HB1xp67_ASAP7_75t_L g1129 ( .A(n_1100), .Y(n_1129) );
OAI32xp33_ASAP7_75t_L g1130 ( .A1(n_1088), .A2(n_1067), .A3(n_1068), .B1(n_1024), .B2(n_1062), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_1108), .B(n_1064), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1084), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1133 ( .A(n_1110), .B(n_1056), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1111), .B(n_1076), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1105), .B(n_1069), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1105), .B(n_1069), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1081), .B(n_1069), .Y(n_1137) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_1103), .B(n_1076), .Y(n_1138) );
OR2x2_ASAP7_75t_L g1139 ( .A(n_1088), .B(n_1065), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1081), .B(n_1058), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1086), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1086), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_1087), .B(n_1077), .Y(n_1143) );
AO22x1_ASAP7_75t_L g1144 ( .A1(n_1129), .A2(n_1088), .B1(n_1018), .B2(n_1098), .Y(n_1144) );
AOI221xp5_ASAP7_75t_L g1145 ( .A1(n_1130), .A2(n_1109), .B1(n_1028), .B2(n_1082), .C(n_1096), .Y(n_1145) );
OAI21xp5_ASAP7_75t_L g1146 ( .A1(n_1123), .A2(n_1033), .B(n_1018), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1114), .Y(n_1147) );
OAI21xp5_ASAP7_75t_L g1148 ( .A1(n_1115), .A2(n_1033), .B(n_1073), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1116), .B(n_1082), .Y(n_1149) );
INVx2_ASAP7_75t_L g1150 ( .A(n_1121), .Y(n_1150) );
BUFx2_ASAP7_75t_L g1151 ( .A(n_1124), .Y(n_1151) );
OA21x2_ASAP7_75t_L g1152 ( .A1(n_1119), .A2(n_1074), .B(n_1080), .Y(n_1152) );
NAND2xp5_ASAP7_75t_SL g1153 ( .A(n_1124), .B(n_1094), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1114), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1116), .B(n_1096), .Y(n_1155) );
NOR2x1_ASAP7_75t_SL g1156 ( .A(n_1139), .B(n_1092), .Y(n_1156) );
OAI221xp5_ASAP7_75t_SL g1157 ( .A1(n_1118), .A2(n_1092), .B1(n_1007), .B2(n_1102), .C(n_1062), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_1120), .B(n_1077), .Y(n_1158) );
OAI22xp33_ASAP7_75t_L g1159 ( .A1(n_1124), .A2(n_1092), .B1(n_1068), .B2(n_1025), .Y(n_1159) );
NAND2xp5_ASAP7_75t_SL g1160 ( .A(n_1125), .B(n_1094), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1120), .B(n_1066), .Y(n_1161) );
OAI21xp5_ASAP7_75t_L g1162 ( .A1(n_1127), .A2(n_1073), .B(n_1039), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1117), .Y(n_1163) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1117), .Y(n_1164) );
AOI221xp5_ASAP7_75t_L g1165 ( .A1(n_1157), .A2(n_1130), .B1(n_1138), .B2(n_1133), .C(n_1134), .Y(n_1165) );
OAI211xp5_ASAP7_75t_SL g1166 ( .A1(n_1145), .A2(n_1146), .B(n_1160), .C(n_1153), .Y(n_1166) );
NOR2x1_ASAP7_75t_L g1167 ( .A(n_1151), .B(n_1068), .Y(n_1167) );
OAI21xp5_ASAP7_75t_L g1168 ( .A1(n_1146), .A2(n_1125), .B(n_1139), .Y(n_1168) );
A2O1A1Ixp33_ASAP7_75t_L g1169 ( .A1(n_1151), .A2(n_1106), .B(n_1113), .C(n_1098), .Y(n_1169) );
AOI222xp33_ASAP7_75t_L g1170 ( .A1(n_1147), .A2(n_1143), .B1(n_1135), .B2(n_1136), .C1(n_1137), .C2(n_1140), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1147), .Y(n_1171) );
XNOR2x1_ASAP7_75t_L g1172 ( .A(n_1144), .B(n_1125), .Y(n_1172) );
AOI21xp5_ASAP7_75t_L g1173 ( .A1(n_1144), .A2(n_1041), .B(n_1092), .Y(n_1173) );
OAI32xp33_ASAP7_75t_L g1174 ( .A1(n_1164), .A2(n_1126), .A3(n_1131), .B1(n_1136), .B2(n_1135), .Y(n_1174) );
AOI21xp33_ASAP7_75t_L g1175 ( .A1(n_1159), .A2(n_950), .B(n_1044), .Y(n_1175) );
AOI21xp5_ASAP7_75t_SL g1176 ( .A1(n_1156), .A2(n_1041), .B(n_1098), .Y(n_1176) );
AOI222xp33_ASAP7_75t_L g1177 ( .A1(n_1154), .A2(n_1137), .B1(n_1140), .B2(n_1142), .C1(n_1132), .C2(n_1128), .Y(n_1177) );
AOI21x1_ASAP7_75t_L g1178 ( .A1(n_1148), .A2(n_1121), .B(n_1039), .Y(n_1178) );
NOR4xp75_ASAP7_75t_L g1179 ( .A(n_1168), .B(n_1162), .C(n_1158), .D(n_1161), .Y(n_1179) );
NOR2xp33_ASAP7_75t_SL g1180 ( .A(n_1173), .B(n_950), .Y(n_1180) );
OAI22xp5_ASAP7_75t_L g1181 ( .A1(n_1169), .A2(n_1164), .B1(n_1163), .B2(n_1154), .Y(n_1181) );
NAND2xp33_ASAP7_75t_R g1182 ( .A(n_1173), .B(n_1152), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1177), .B(n_1152), .Y(n_1183) );
XOR2xp5_ASAP7_75t_L g1184 ( .A(n_1172), .B(n_1156), .Y(n_1184) );
AOI21xp5_ASAP7_75t_L g1185 ( .A1(n_1166), .A2(n_1152), .B(n_1163), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1170), .B(n_1149), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1167), .B(n_1149), .Y(n_1187) );
AOI22xp5_ASAP7_75t_L g1188 ( .A1(n_1165), .A2(n_1152), .B1(n_1113), .B2(n_1155), .Y(n_1188) );
NAND3xp33_ASAP7_75t_SL g1189 ( .A(n_1180), .B(n_1171), .C(n_982), .Y(n_1189) );
NAND2xp5_ASAP7_75t_SL g1190 ( .A(n_1180), .B(n_1178), .Y(n_1190) );
NOR3xp33_ASAP7_75t_L g1191 ( .A(n_1183), .B(n_1174), .C(n_1175), .Y(n_1191) );
NOR2xp67_ASAP7_75t_L g1192 ( .A(n_1185), .B(n_1150), .Y(n_1192) );
AND4x1_ASAP7_75t_L g1193 ( .A(n_1188), .B(n_1176), .C(n_1155), .D(n_990), .Y(n_1193) );
NAND3xp33_ASAP7_75t_SL g1194 ( .A(n_1179), .B(n_982), .C(n_963), .Y(n_1194) );
NOR3xp33_ASAP7_75t_L g1195 ( .A(n_1181), .B(n_982), .C(n_981), .Y(n_1195) );
NAND3xp33_ASAP7_75t_SL g1196 ( .A(n_1191), .B(n_1184), .C(n_1186), .Y(n_1196) );
NOR2x2_ASAP7_75t_L g1197 ( .A(n_1193), .B(n_1182), .Y(n_1197) );
XNOR2xp5_ASAP7_75t_L g1198 ( .A(n_1194), .B(n_1187), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1189), .Y(n_1199) );
AND4x1_ASAP7_75t_L g1200 ( .A(n_1195), .B(n_990), .C(n_961), .D(n_1102), .Y(n_1200) );
XNOR2xp5_ASAP7_75t_L g1201 ( .A(n_1196), .B(n_1190), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1198), .B(n_1192), .Y(n_1202) );
INVx1_ASAP7_75t_SL g1203 ( .A(n_1199), .Y(n_1203) );
XNOR2xp5_ASAP7_75t_L g1204 ( .A(n_1200), .B(n_961), .Y(n_1204) );
XNOR2xp5_ASAP7_75t_L g1205 ( .A(n_1201), .B(n_1197), .Y(n_1205) );
BUFx2_ASAP7_75t_L g1206 ( .A(n_1202), .Y(n_1206) );
XNOR2xp5_ASAP7_75t_L g1207 ( .A(n_1204), .B(n_1197), .Y(n_1207) );
BUFx2_ASAP7_75t_L g1208 ( .A(n_1206), .Y(n_1208) );
OAI22x1_ASAP7_75t_L g1209 ( .A1(n_1205), .A2(n_1203), .B1(n_1113), .B2(n_1150), .Y(n_1209) );
INVxp67_ASAP7_75t_SL g1210 ( .A(n_1208), .Y(n_1210) );
AOI221xp5_ASAP7_75t_L g1211 ( .A1(n_1209), .A2(n_1207), .B1(n_1150), .B2(n_977), .C(n_1141), .Y(n_1211) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1210), .Y(n_1212) );
AOI21xp5_ASAP7_75t_L g1213 ( .A1(n_1212), .A2(n_1211), .B(n_1015), .Y(n_1213) );
AOI21xp5_ASAP7_75t_L g1214 ( .A1(n_1213), .A2(n_1122), .B(n_1080), .Y(n_1214) );
endmodule