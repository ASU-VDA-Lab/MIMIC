module fake_jpeg_28940_n_542 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_542);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_542;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_59),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_61),
.B(n_102),
.Y(n_118)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_64),
.B(n_66),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

BUFx4f_ASAP7_75t_SL g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_70),
.Y(n_160)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_83),
.Y(n_157)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_26),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_99),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_0),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_101),
.Y(n_141)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_98),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_20),
.B(n_1),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_100),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_20),
.B(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_26),
.B(n_2),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_47),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_104),
.B(n_106),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_99),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_150),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_86),
.B1(n_103),
.B2(n_97),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_117),
.A2(n_129),
.B1(n_130),
.B2(n_132),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

AND2x4_ASAP7_75t_L g125 ( 
.A(n_55),
.B(n_40),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_125),
.B(n_40),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_89),
.A2(n_29),
.B1(n_48),
.B2(n_37),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_69),
.A2(n_29),
.B1(n_48),
.B2(n_37),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_78),
.A2(n_29),
.B1(n_48),
.B2(n_37),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_53),
.B(n_51),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_158),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_58),
.A2(n_45),
.B1(n_36),
.B2(n_29),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_138),
.A2(n_140),
.B1(n_90),
.B2(n_88),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_54),
.A2(n_45),
.B1(n_48),
.B2(n_37),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_59),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_93),
.A2(n_45),
.B1(n_47),
.B2(n_24),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_152),
.A2(n_40),
.B1(n_24),
.B2(n_41),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_65),
.B(n_51),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_56),
.B(n_49),
.C(n_44),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_24),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_169),
.A2(n_218),
.B1(n_152),
.B2(n_129),
.Y(n_236)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_171),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g172 ( 
.A1(n_119),
.A2(n_105),
.B1(n_79),
.B2(n_92),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_172),
.A2(n_206),
.B1(n_221),
.B2(n_143),
.Y(n_255)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_173),
.Y(n_239)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_174),
.Y(n_241)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_175),
.Y(n_246)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_177),
.Y(n_251)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_178),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_165),
.A2(n_57),
.B1(n_63),
.B2(n_100),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_179),
.A2(n_190),
.B1(n_203),
.B2(n_213),
.Y(n_243)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_180),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_110),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_181),
.B(n_194),
.Y(n_233)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_185),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_118),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_186),
.B(n_192),
.Y(n_229)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_187),
.Y(n_264)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_188),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_189),
.B(n_215),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_131),
.A2(n_73),
.B1(n_76),
.B2(n_83),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_191),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_30),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_30),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_193),
.B(n_196),
.Y(n_271)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_120),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_197),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_166),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_147),
.B(n_35),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_201),
.Y(n_240)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_199),
.Y(n_247)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_122),
.B(n_35),
.Y(n_201)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_204),
.B(n_207),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_123),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_108),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_208),
.B(n_209),
.Y(n_268)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_122),
.B(n_49),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_210),
.B(n_228),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_110),
.B(n_44),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_211),
.Y(n_253)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_112),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_159),
.B(n_87),
.C(n_80),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_154),
.C(n_149),
.Y(n_256)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_121),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_114),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_217),
.Y(n_244)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_148),
.A2(n_45),
.B1(n_52),
.B2(n_41),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_161),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_223),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_107),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_220),
.A2(n_224),
.B1(n_227),
.B2(n_127),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_151),
.A2(n_52),
.B1(n_41),
.B2(n_38),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_113),
.A2(n_52),
.B1(n_38),
.B2(n_27),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_222),
.A2(n_132),
.B1(n_130),
.B2(n_160),
.Y(n_274)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_126),
.Y(n_223)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_145),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_112),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_226),
.Y(n_248)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_126),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_123),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_236),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_182),
.B(n_125),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_242),
.B(n_257),
.C(n_260),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_250),
.B(n_255),
.Y(n_285)
);

OA22x2_ASAP7_75t_SL g254 ( 
.A1(n_202),
.A2(n_125),
.B1(n_138),
.B2(n_140),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_254),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_256),
.B(n_9),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_127),
.C(n_143),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_181),
.B(n_109),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_262),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_214),
.B(n_176),
.C(n_178),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_169),
.A2(n_27),
.B(n_38),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_261),
.A2(n_219),
.B(n_4),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_180),
.B(n_109),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_212),
.B(n_149),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_266),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_206),
.B(n_27),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_179),
.B(n_3),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_267),
.Y(n_286)
);

AND2x2_ASAP7_75t_SL g269 ( 
.A(n_195),
.B(n_40),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_185),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_200),
.B(n_3),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_272),
.B(n_17),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_274),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_304)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_277),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_222),
.B(n_190),
.C(n_205),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_278),
.A2(n_279),
.B(n_288),
.Y(n_334)
);

AND2x4_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_215),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_280),
.B(n_296),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_217),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_281),
.B(n_291),
.C(n_297),
.Y(n_339)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_232),
.Y(n_282)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_282),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_234),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_283),
.B(n_293),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_266),
.A2(n_172),
.B1(n_216),
.B2(n_203),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_284),
.A2(n_298),
.B1(n_306),
.B2(n_317),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_267),
.A2(n_261),
.B(n_237),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_287),
.A2(n_244),
.B(n_269),
.Y(n_337)
);

AO21x2_ASAP7_75t_L g289 ( 
.A1(n_236),
.A2(n_224),
.B(n_225),
.Y(n_289)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_289),
.A2(n_258),
.B(n_264),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_205),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_290),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_191),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_238),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_274),
.A2(n_170),
.B(n_209),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_294),
.A2(n_308),
.B(n_12),
.Y(n_353)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_237),
.B(n_199),
.C(n_32),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_256),
.B(n_213),
.C(n_154),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_254),
.A2(n_42),
.B1(n_32),
.B2(n_5),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_299),
.A2(n_312),
.B1(n_270),
.B2(n_252),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_249),
.B(n_32),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_300),
.B(n_303),
.Y(n_325)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_232),
.Y(n_301)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_301),
.Y(n_332)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_302),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_238),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_304),
.A2(n_269),
.B1(n_230),
.B2(n_270),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_257),
.B(n_233),
.C(n_229),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_305),
.B(n_310),
.C(n_286),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_254),
.A2(n_32),
.B1(n_6),
.B2(n_7),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_237),
.A2(n_32),
.B1(n_6),
.B2(n_8),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_250),
.B(n_5),
.C(n_8),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_316),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_254),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_275),
.Y(n_313)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_313),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_231),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_314),
.Y(n_358)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_235),
.Y(n_315)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_315),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_272),
.B(n_265),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_255),
.A2(n_243),
.B1(n_271),
.B2(n_248),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_318),
.B(n_11),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_253),
.B(n_11),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_235),
.Y(n_345)
);

AOI32xp33_ASAP7_75t_L g320 ( 
.A1(n_287),
.A2(n_253),
.A3(n_240),
.B1(n_268),
.B2(n_230),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_320),
.B(n_352),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_321),
.A2(n_298),
.B1(n_306),
.B2(n_289),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_322),
.A2(n_331),
.B1(n_335),
.B2(n_357),
.Y(n_364)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_295),
.B(n_244),
.C(n_276),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_328),
.B(n_347),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_291),
.B(n_244),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_329),
.B(n_339),
.C(n_281),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_309),
.A2(n_248),
.B1(n_252),
.B2(n_270),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_309),
.A2(n_247),
.B1(n_245),
.B2(n_264),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_336),
.A2(n_279),
.B1(n_304),
.B2(n_302),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g373 ( 
.A(n_337),
.B(n_280),
.CI(n_318),
.CON(n_373),
.SN(n_373)
);

AOI32xp33_ASAP7_75t_SL g338 ( 
.A1(n_278),
.A2(n_258),
.A3(n_276),
.B1(n_245),
.B2(n_247),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_338),
.A2(n_353),
.B(n_294),
.Y(n_359)
);

XNOR2x1_ASAP7_75t_L g382 ( 
.A(n_341),
.B(n_318),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_319),
.B(n_231),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_342),
.B(n_354),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_345),
.B(n_346),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_307),
.B(n_273),
.Y(n_346)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_279),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_348),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_307),
.B(n_273),
.Y(n_349)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_349),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_292),
.B(n_251),
.Y(n_350)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_350),
.Y(n_390)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_292),
.Y(n_351)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_351),
.Y(n_392)
);

BUFx5_ASAP7_75t_L g352 ( 
.A(n_313),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_251),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_288),
.A2(n_246),
.B(n_241),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_355),
.A2(n_285),
.B(n_308),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_312),
.A2(n_246),
.B1(n_241),
.B2(n_239),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_359),
.A2(n_387),
.B(n_345),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_295),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_360),
.B(n_368),
.C(n_375),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_361),
.A2(n_362),
.B(n_366),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_334),
.A2(n_289),
.B(n_285),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_324),
.A2(n_289),
.B1(n_299),
.B2(n_317),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_363),
.A2(n_383),
.B1(n_385),
.B2(n_322),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_334),
.A2(n_289),
.B(n_285),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_367),
.B(n_388),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_325),
.B(n_305),
.Y(n_372)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_372),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_373),
.B(n_378),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_327),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_376),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_330),
.B(n_297),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_327),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_330),
.B(n_296),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_344),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_380),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_350),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_381),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_337),
.C(n_323),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_328),
.B(n_329),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_332),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_324),
.A2(n_310),
.B1(n_279),
.B2(n_284),
.Y(n_385)
);

OAI31xp33_ASAP7_75t_L g386 ( 
.A1(n_353),
.A2(n_311),
.A3(n_314),
.B(n_315),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g396 ( 
.A(n_386),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_356),
.A2(n_239),
.B1(n_13),
.B2(n_15),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_336),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_351),
.B(n_12),
.Y(n_389)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_389),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_326),
.B(n_323),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_393),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_326),
.B(n_12),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_393),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_394),
.B(n_416),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_384),
.B(n_341),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_398),
.B(n_400),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_360),
.B(n_354),
.C(n_346),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_402),
.B(n_407),
.C(n_409),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_370),
.B(n_349),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_415),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_404),
.A2(n_410),
.B1(n_419),
.B2(n_367),
.Y(n_427)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_392),
.Y(n_406)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_406),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_355),
.C(n_331),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_369),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_408),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_375),
.B(n_335),
.C(n_347),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_338),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_379),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_336),
.Y(n_417)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_417),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_418),
.B(n_373),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_363),
.A2(n_332),
.B1(n_358),
.B2(n_333),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_392),
.Y(n_420)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_420),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_383),
.A2(n_358),
.B1(n_333),
.B2(n_340),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_422),
.Y(n_426)
);

NAND2x1_ASAP7_75t_SL g423 ( 
.A(n_377),
.B(n_352),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_423),
.A2(n_359),
.B(n_366),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_382),
.B(n_340),
.C(n_343),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_424),
.B(n_370),
.C(n_373),
.Y(n_441)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_427),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_396),
.A2(n_410),
.B1(n_385),
.B2(n_388),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_429),
.A2(n_438),
.B1(n_440),
.B2(n_422),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_405),
.B(n_380),
.Y(n_430)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_430),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_423),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_431),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_417),
.B(n_381),
.Y(n_432)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_432),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_397),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_434),
.B(n_439),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_404),
.A2(n_371),
.B1(n_364),
.B2(n_387),
.Y(n_435)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_435),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_436),
.A2(n_411),
.B(n_343),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_413),
.A2(n_362),
.B1(n_361),
.B2(n_377),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_414),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_408),
.A2(n_369),
.B1(n_390),
.B2(n_364),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_441),
.B(n_451),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_406),
.Y(n_443)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_443),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_401),
.B(n_389),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_445),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_446),
.B(n_395),
.Y(n_459)
);

AOI21xp33_ASAP7_75t_L g448 ( 
.A1(n_414),
.A2(n_365),
.B(n_386),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_448),
.A2(n_421),
.B1(n_390),
.B2(n_411),
.Y(n_464)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_420),
.Y(n_449)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_449),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_399),
.B(n_365),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_452),
.A2(n_461),
.B1(n_426),
.B2(n_470),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_451),
.B(n_399),
.C(n_424),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_453),
.B(n_454),
.C(n_455),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_398),
.C(n_407),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_402),
.C(n_409),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g485 ( 
.A(n_459),
.B(n_464),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_441),
.B(n_418),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_460),
.B(n_465),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_444),
.B(n_400),
.C(n_403),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_463),
.B(n_468),
.C(n_472),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_444),
.B(n_415),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_395),
.C(n_412),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_442),
.B(n_412),
.C(n_419),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_438),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_439),
.Y(n_474)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_474),
.Y(n_505)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_467),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_475),
.B(n_476),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_432),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_462),
.Y(n_477)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_477),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_458),
.B(n_434),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_478),
.B(n_480),
.Y(n_502)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_462),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_479),
.A2(n_425),
.B1(n_449),
.B2(n_447),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_455),
.B(n_450),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_433),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_447),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_483),
.A2(n_489),
.B1(n_490),
.B2(n_488),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_453),
.B(n_426),
.C(n_431),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_487),
.B(n_454),
.C(n_456),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_461),
.A2(n_436),
.B(n_433),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_488),
.A2(n_473),
.B(n_437),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_452),
.A2(n_437),
.B1(n_429),
.B2(n_440),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_490),
.B(n_472),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_491),
.B(n_493),
.Y(n_515)
);

INVxp33_ASAP7_75t_L g514 ( 
.A(n_492),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_484),
.B(n_468),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_495),
.B(n_497),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_484),
.A2(n_463),
.B(n_471),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_496),
.A2(n_13),
.B(n_15),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_456),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_485),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_474),
.A2(n_482),
.B(n_476),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_500),
.A2(n_13),
.B(n_16),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_501),
.A2(n_16),
.B1(n_17),
.B2(n_505),
.Y(n_518)
);

BUFx24_ASAP7_75t_SL g503 ( 
.A(n_483),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_503),
.B(n_489),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_481),
.B(n_460),
.C(n_465),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_504),
.B(n_486),
.C(n_485),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_425),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_502),
.B(n_481),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_510),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_508),
.B(n_509),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_511),
.B(n_512),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_459),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_446),
.C(n_15),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_513),
.B(n_499),
.Y(n_522)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_516),
.Y(n_521)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_517),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_518),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_522),
.B(n_523),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_519),
.B(n_494),
.Y(n_523)
);

A2O1A1Ixp33_ASAP7_75t_L g528 ( 
.A1(n_514),
.A2(n_500),
.B(n_497),
.C(n_491),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_528),
.B(n_509),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_527),
.B(n_514),
.Y(n_529)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_529),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_515),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_531),
.B(n_533),
.C(n_515),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_532),
.A2(n_530),
.B(n_513),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_528),
.A2(n_508),
.B(n_526),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_534),
.B(n_531),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_536),
.A2(n_524),
.B(n_521),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_537),
.B(n_538),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_539),
.B(n_535),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_520),
.B1(n_504),
.B2(n_493),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_520),
.Y(n_542)
);


endmodule