module real_aes_16711_n_10 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
output n_10;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_13;
wire n_41;
wire n_34;
wire n_12;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_50;
wire n_29;
wire n_20;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
INVx2_ASAP7_75t_L g19 ( .A(n_0), .Y(n_19) );
INVx1_ASAP7_75t_L g23 ( .A(n_1), .Y(n_23) );
BUFx3_ASAP7_75t_L g35 ( .A(n_2), .Y(n_35) );
AND2x2_ASAP7_75t_L g14 ( .A(n_3), .B(n_9), .Y(n_14) );
BUFx6f_ASAP7_75t_L g30 ( .A(n_4), .Y(n_30) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
AND2x2_ASAP7_75t_L g39 ( .A(n_5), .B(n_23), .Y(n_39) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_6), .B(n_17), .Y(n_16) );
BUFx6f_ASAP7_75t_L g28 ( .A(n_7), .Y(n_28) );
INVx1_ASAP7_75t_L g33 ( .A(n_8), .Y(n_33) );
AOI221xp5_ASAP7_75t_L g10 ( .A1(n_11), .A2(n_34), .B1(n_36), .B2(n_40), .C(n_47), .Y(n_10) );
NAND3xp33_ASAP7_75t_L g11 ( .A(n_12), .B(n_24), .C(n_31), .Y(n_11) );
AOI221xp5_ASAP7_75t_SL g12 ( .A1(n_13), .A2(n_15), .B1(n_16), .B2(n_20), .C(n_21), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_14), .Y(n_13) );
AND2x2_ASAP7_75t_L g38 ( .A(n_14), .B(n_39), .Y(n_38) );
INVx1_ASAP7_75t_L g20 ( .A(n_15), .Y(n_20) );
NOR2xp33_ASAP7_75t_L g49 ( .A(n_15), .B(n_21), .Y(n_49) );
INVxp67_ASAP7_75t_SL g50 ( .A(n_16), .Y(n_50) );
INVx2_ASAP7_75t_SL g17 ( .A(n_18), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
INVx1_ASAP7_75t_L g21 ( .A(n_22), .Y(n_21) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
INVx1_ASAP7_75t_L g24 ( .A(n_25), .Y(n_24) );
INVx3_ASAP7_75t_L g25 ( .A(n_26), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_27), .B(n_29), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_28), .Y(n_27) );
OR2x2_ASAP7_75t_L g44 ( .A(n_28), .B(n_30), .Y(n_44) );
INVx1_ASAP7_75t_L g29 ( .A(n_30), .Y(n_29) );
INVx1_ASAP7_75t_L g31 ( .A(n_32), .Y(n_31) );
NOR2xp33_ASAP7_75t_L g36 ( .A(n_32), .B(n_37), .Y(n_36) );
INVx1_ASAP7_75t_L g32 ( .A(n_33), .Y(n_32) );
BUFx2_ASAP7_75t_L g34 ( .A(n_35), .Y(n_34) );
INVx2_ASAP7_75t_L g46 ( .A(n_35), .Y(n_46) );
INVxp67_ASAP7_75t_L g37 ( .A(n_38), .Y(n_37) );
INVx3_ASAP7_75t_L g40 ( .A(n_41), .Y(n_40) );
OR2x6_ASAP7_75t_L g41 ( .A(n_42), .B(n_45), .Y(n_41) );
INVx2_ASAP7_75t_L g42 ( .A(n_43), .Y(n_42) );
INVx3_ASAP7_75t_L g43 ( .A(n_44), .Y(n_43) );
INVxp67_ASAP7_75t_L g45 ( .A(n_46), .Y(n_45) );
INVx1_ASAP7_75t_L g47 ( .A(n_48), .Y(n_47) );
NAND2xp5_ASAP7_75t_L g48 ( .A(n_49), .B(n_50), .Y(n_48) );
endmodule