module real_jpeg_11372_n_17 (n_301, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_301;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_249;
wire n_286;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_243;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_295;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_4),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_4),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_43),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_4),
.A2(n_43),
.B1(n_63),
.B2(n_64),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_6),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_56),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_56),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_7),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_8),
.A2(n_63),
.B1(n_64),
.B2(n_72),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_8),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_72),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_72),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_9),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_9),
.A2(n_63),
.B1(n_64),
.B2(n_87),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_9),
.A2(n_39),
.B1(n_40),
.B2(n_87),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_87),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_10),
.A2(n_63),
.B1(n_64),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_10),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_153),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_153),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_153),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_12),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_12),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_62),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_62),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_13),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_13),
.B(n_29),
.C(n_67),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_13),
.B(n_85),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_13),
.A2(n_97),
.B(n_157),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_13),
.A2(n_46),
.B(n_84),
.C(n_184),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_141),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_13),
.B(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_13),
.B(n_39),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_14),
.A2(n_39),
.B1(n_40),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_14),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_106),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_14),
.A2(n_63),
.B1(n_64),
.B2(n_106),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_106),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_15),
.A2(n_35),
.B1(n_63),
.B2(n_64),
.Y(n_78)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_128),
.B1(n_298),
.B2(n_299),
.Y(n_18)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_19),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_126),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_109),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_21),
.B(n_109),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_75),
.C(n_91),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_22),
.A2(n_23),
.B1(n_75),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_58),
.B2(n_74),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_36),
.B1(n_37),
.B2(n_57),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_26),
.A2(n_37),
.B(n_74),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_26),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_32),
.B(n_33),
.Y(n_26)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_27),
.A2(n_32),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_27),
.B(n_158),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_27),
.A2(n_32),
.B1(n_96),
.B2(n_246),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_28),
.A2(n_29),
.B1(n_67),
.B2(n_68),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_28),
.B(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_32),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_32),
.B(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_34),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_44),
.B(n_50),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_38),
.A2(n_44),
.B1(n_52),
.B2(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_40),
.B1(n_45),
.B2(n_49),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_40),
.A2(n_52),
.B(n_141),
.C(n_228),
.Y(n_227)
);

AOI32xp33_ASAP7_75t_L g241 ( 
.A1(n_40),
.A2(n_46),
.A3(n_49),
.B1(n_229),
.B2(n_242),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_44),
.B(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_44),
.B(n_55),
.Y(n_108)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_44),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_44),
.A2(n_50),
.B(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_44),
.A2(n_52),
.B1(n_105),
.B2(n_256),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_44)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NAND2xp33_ASAP7_75t_SL g242 ( 
.A(n_45),
.B(n_47),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_47),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_52),
.A2(n_105),
.B(n_107),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_65),
.B1(n_70),
.B2(n_73),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_65),
.B1(n_73),
.B2(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

AO22x1_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_64),
.B1(n_83),
.B2(n_84),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_63),
.B(n_145),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_64),
.A2(n_83),
.B(n_141),
.Y(n_184)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_65),
.A2(n_73),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_65),
.B(n_143),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_65),
.A2(n_73),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_65),
.A2(n_73),
.B1(n_101),
.B2(n_235),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_69),
.A2(n_71),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_69),
.A2(n_152),
.B(n_154),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_69),
.B(n_141),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_69),
.A2(n_154),
.B(n_234),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_73),
.B(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_75),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_79),
.B(n_90),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_79),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_SL g139 ( 
.A1(n_77),
.A2(n_140),
.B(n_142),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_77),
.A2(n_142),
.B(n_217),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_86),
.B1(n_88),
.B2(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_80),
.A2(n_189),
.B(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_80),
.A2(n_88),
.B1(n_204),
.B2(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_80),
.A2(n_190),
.B(n_232),
.Y(n_254)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_85),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_81),
.B(n_191),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_85),
.B(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_88),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_88),
.A2(n_103),
.B(n_205),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_91),
.B(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_102),
.C(n_104),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_92),
.A2(n_93),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_99),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_94),
.A2(n_99),
.B1(n_100),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_94),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_97),
.A2(n_156),
.B(n_157),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_97),
.A2(n_98),
.B1(n_186),
.B2(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_97),
.A2(n_98),
.B1(n_212),
.B2(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_98),
.A2(n_163),
.B(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_98),
.B(n_141),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_98),
.A2(n_171),
.B(n_186),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_102),
.B(n_104),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_108),
.B(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_125),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_117),
.Y(n_124)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_128),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_292),
.B(n_297),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_280),
.B(n_291),
.Y(n_130)
);

OAI321xp33_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_248),
.A3(n_273),
.B1(n_278),
.B2(n_279),
.C(n_301),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_221),
.B(n_247),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_198),
.B(n_220),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_179),
.B(n_197),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_159),
.B(n_178),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_146),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_137),
.B(n_146),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_144),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_138),
.A2(n_139),
.B1(n_144),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_144),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_155),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_151),
.C(n_155),
.Y(n_180)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_156),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_167),
.B(n_177),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_165),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_172),
.B(n_176),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_169),
.B(n_170),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_180),
.B(n_181),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_187),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_192),
.C(n_196),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_185),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_187)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_199),
.B(n_200),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_213),
.B2(n_214),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_216),
.C(n_218),
.Y(n_222)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_207),
.C(n_211),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_222),
.B(n_223),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_237),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_224),
.B(n_238),
.C(n_239),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_230),
.B2(n_236),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_231),
.C(n_233),
.Y(n_262)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_230),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_244),
.Y(n_258)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_263),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_263),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_259),
.C(n_262),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_250),
.A2(n_251),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_258),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_257),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_257),
.C(n_258),
.Y(n_272)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_255),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_259),
.B(n_262),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_261),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_272),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_267),
.C(n_272),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_270),
.C(n_271),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_274),
.B(n_275),
.Y(n_278)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_290),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_290),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_285),
.C(n_286),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_294),
.Y(n_297)
);


endmodule