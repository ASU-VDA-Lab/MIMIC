module fake_jpeg_6599_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_L g45 ( 
.A1(n_17),
.A2(n_8),
.B(n_15),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_18),
.C(n_25),
.Y(n_60)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_19),
.B1(n_21),
.B2(n_30),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_36),
.B1(n_31),
.B2(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_34),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_60),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_27),
.B1(n_19),
.B2(n_21),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_27),
.B1(n_21),
.B2(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_43),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_27),
.B1(n_36),
.B2(n_30),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_27),
.B1(n_36),
.B2(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_46),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_68),
.A2(n_86),
.B1(n_90),
.B2(n_93),
.Y(n_115)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_74),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_47),
.B1(n_41),
.B2(n_42),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_79),
.B1(n_80),
.B2(n_87),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_29),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_75),
.B(n_95),
.Y(n_130)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_47),
.B1(n_41),
.B2(n_42),
.Y(n_80)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_42),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_40),
.B(n_38),
.Y(n_121)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_84),
.Y(n_108)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_36),
.B1(n_37),
.B2(n_44),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_92),
.Y(n_102)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_31),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_37),
.B1(n_44),
.B2(n_43),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_55),
.Y(n_105)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_98),
.Y(n_119)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_31),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_29),
.Y(n_111)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_66),
.Y(n_124)
);

OA22x2_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_43),
.B1(n_38),
.B2(n_40),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_44),
.B(n_37),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_43),
.C(n_39),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_128),
.C(n_33),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_70),
.A2(n_43),
.B(n_24),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_122),
.B(n_127),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_18),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_113),
.A2(n_124),
.B1(n_72),
.B2(n_32),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_40),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_121),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_82),
.A2(n_39),
.B(n_40),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_38),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_39),
.Y(n_160)
);

AOI32xp33_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_38),
.A3(n_39),
.B1(n_50),
.B2(n_37),
.Y(n_126)
);

FAx1_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_128),
.CI(n_119),
.CON(n_159),
.SN(n_159)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_39),
.B(n_24),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_71),
.A2(n_24),
.B(n_34),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_133),
.B(n_134),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_104),
.Y(n_134)
);

BUFx4f_ASAP7_75t_SL g135 ( 
.A(n_124),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_140),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_68),
.B1(n_97),
.B2(n_80),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_137),
.A2(n_144),
.B1(n_147),
.B2(n_131),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_91),
.Y(n_139)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_29),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_149),
.Y(n_167)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_146),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_143),
.B(n_111),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_98),
.B1(n_89),
.B2(n_84),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_90),
.Y(n_145)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_93),
.B1(n_100),
.B2(n_85),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_129),
.B(n_88),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_151),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_109),
.A2(n_23),
.B1(n_33),
.B2(n_32),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_150),
.A2(n_159),
.B1(n_161),
.B2(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_155),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_39),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_113),
.B(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_108),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_39),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_160),
.C(n_131),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

AO22x2_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_17),
.B1(n_35),
.B2(n_66),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_158),
.A2(n_129),
.B1(n_112),
.B2(n_115),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_163),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_164),
.B(n_141),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_135),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_166),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_184),
.C(n_154),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_174),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_191),
.B1(n_193),
.B2(n_141),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_135),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_112),
.B1(n_111),
.B2(n_120),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_186),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_158),
.A2(n_120),
.B1(n_118),
.B2(n_107),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_118),
.B1(n_107),
.B2(n_104),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_157),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_179),
.A2(n_0),
.B(n_1),
.Y(n_222)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_182),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_150),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_136),
.A2(n_108),
.B1(n_33),
.B2(n_23),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_149),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_189),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_138),
.A2(n_32),
.B1(n_23),
.B2(n_25),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_138),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_192),
.Y(n_204)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

OA21x2_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_35),
.B(n_50),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_25),
.B1(n_28),
.B2(n_22),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_195),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_175),
.B(n_132),
.Y(n_200)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_207),
.C(n_210),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_202),
.A2(n_212),
.B1(n_217),
.B2(n_218),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_184),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_160),
.C(n_152),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_194),
.B(n_154),
.Y(n_209)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_164),
.B(n_152),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_183),
.A2(n_28),
.B1(n_22),
.B2(n_35),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_190),
.A2(n_35),
.B1(n_50),
.B2(n_11),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_225),
.B(n_187),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_185),
.A2(n_103),
.B1(n_73),
.B2(n_50),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_173),
.A2(n_103),
.B1(n_73),
.B2(n_2),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_220),
.A2(n_223),
.B(n_165),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_172),
.B1(n_163),
.B2(n_174),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_222),
.A2(n_187),
.B(n_169),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_0),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_7),
.C(n_14),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_226),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_220),
.A2(n_219),
.B1(n_206),
.B2(n_166),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_227),
.A2(n_230),
.B1(n_245),
.B2(n_223),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_162),
.B1(n_179),
.B2(n_176),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_171),
.B1(n_188),
.B2(n_193),
.Y(n_231)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_231),
.Y(n_265)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_224),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_237),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_201),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_238),
.A2(n_239),
.B(n_246),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_204),
.A2(n_193),
.B(n_179),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_203),
.A2(n_169),
.B1(n_165),
.B2(n_167),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_167),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_237),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_224),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_214),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_207),
.B(n_167),
.C(n_1),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_210),
.C(n_205),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_248),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_266),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_257),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_244),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_202),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_213),
.C(n_198),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_264),
.C(n_267),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_259),
.A2(n_268),
.B1(n_229),
.B2(n_247),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_234),
.B(n_225),
.Y(n_261)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_215),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_272),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_199),
.C(n_216),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_235),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_217),
.C(n_218),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_239),
.A2(n_197),
.B(n_221),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_212),
.C(n_222),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_232),
.C(n_240),
.Y(n_285)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_238),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_271),
.A2(n_241),
.B1(n_242),
.B2(n_233),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_16),
.Y(n_272)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_273),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_275),
.A2(n_276),
.B(n_278),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_263),
.A2(n_228),
.B(n_251),
.Y(n_278)
);

NOR2xp67_ASAP7_75t_SL g279 ( 
.A(n_253),
.B(n_251),
.Y(n_279)
);

XOR2x1_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_12),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_240),
.Y(n_281)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_287),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_290),
.C(n_9),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_16),
.Y(n_287)
);

XOR2x2_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_0),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_288),
.B(n_1),
.Y(n_298)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_258),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_9),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_280),
.A2(n_265),
.B1(n_260),
.B2(n_267),
.Y(n_291)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_291),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_284),
.Y(n_293)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_293),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_286),
.B(n_272),
.Y(n_294)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_294),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_295),
.A2(n_298),
.B(n_3),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_278),
.A2(n_264),
.B1(n_255),
.B2(n_254),
.Y(n_296)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_296),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_274),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_277),
.B(n_282),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_301),
.A2(n_304),
.B(n_13),
.Y(n_309)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_282),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_306),
.A2(n_307),
.B(n_310),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_277),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_309),
.A2(n_317),
.B1(n_298),
.B2(n_4),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_274),
.B(n_13),
.Y(n_310)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_313),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_14),
.B(n_16),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_3),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_291),
.C(n_305),
.Y(n_318)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_318),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_314),
.Y(n_319)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_319),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_301),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_325),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_322),
.B(n_324),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_302),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_302),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_326),
.B(n_3),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_328),
.A2(n_331),
.B(n_321),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_323),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_333),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_318),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_325),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_334),
.B(n_335),
.Y(n_337)
);

OAI321xp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_332),
.A3(n_330),
.B1(n_327),
.B2(n_6),
.C(n_5),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_4),
.C(n_5),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_6),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_6),
.C(n_339),
.Y(n_341)
);


endmodule