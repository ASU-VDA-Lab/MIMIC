module fake_jpeg_4933_n_177 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_15),
.Y(n_49)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_26),
.B1(n_28),
.B2(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_47),
.B1(n_51),
.B2(n_17),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_26),
.B1(n_14),
.B2(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_49),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_26),
.B1(n_14),
.B2(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_17),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_63),
.Y(n_78)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_67),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_16),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_41),
.B1(n_40),
.B2(n_42),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_23),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_23),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_25),
.B(n_10),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_71),
.B1(n_79),
.B2(n_64),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_69),
.A2(n_58),
.B1(n_61),
.B2(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_42),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_41),
.B1(n_43),
.B2(n_48),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_67),
.B1(n_16),
.B2(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_63),
.B(n_41),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_83),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_53),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_54),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_68),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_91),
.B1(n_96),
.B2(n_16),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_64),
.B1(n_62),
.B2(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_85),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_70),
.B1(n_81),
.B2(n_75),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_77),
.C(n_74),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_98),
.C(n_100),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_80),
.C(n_78),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_25),
.B(n_53),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_16),
.B(n_20),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_31),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_54),
.C(n_31),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_82),
.C(n_73),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_107),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

AOI322xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_72),
.A3(n_98),
.B1(n_90),
.B2(n_94),
.C1(n_87),
.C2(n_100),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_72),
.B(n_79),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_25),
.B(n_19),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_16),
.Y(n_110)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_111),
.A2(n_65),
.B1(n_19),
.B2(n_20),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_19),
.B(n_20),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_97),
.B(n_101),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_115),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_67),
.Y(n_116)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_130),
.B(n_0),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_65),
.B1(n_19),
.B2(n_30),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_125),
.A2(n_116),
.B1(n_112),
.B2(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_104),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_128),
.A2(n_131),
.B1(n_46),
.B2(n_20),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_65),
.B1(n_20),
.B2(n_46),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_132),
.B(n_134),
.Y(n_150)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_102),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_136),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_141),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_111),
.B1(n_106),
.B2(n_108),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_122),
.B1(n_124),
.B2(n_127),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_103),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_140),
.C(n_129),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_113),
.C(n_46),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_143),
.B(n_119),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_136),
.C(n_12),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_152),
.B1(n_150),
.B2(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_151),
.Y(n_160)
);

AOI31xp67_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_122),
.A3(n_118),
.B(n_3),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_SL g157 ( 
.A(n_148),
.B(n_11),
.C(n_3),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_140),
.Y(n_151)
);

OAI22x1_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_118),
.B1(n_2),
.B2(n_3),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_153),
.Y(n_154)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_158),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_156),
.B(n_4),
.Y(n_164)
);

AOI31xp33_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_4),
.A3(n_5),
.B(n_6),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_152),
.A2(n_151),
.B1(n_146),
.B2(n_11),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_146),
.B(n_1),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_161),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_1),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_156),
.B(n_157),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_163),
.A2(n_7),
.B(n_8),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_5),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_7),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_170),
.B(n_171),
.C(n_163),
.Y(n_173)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_166),
.Y(n_175)
);

NOR2xp67_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_162),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_9),
.B(n_172),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.Y(n_177)
);


endmodule