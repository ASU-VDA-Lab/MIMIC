module fake_jpeg_6799_n_252 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_45;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_36),
.Y(n_43)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_13),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_25),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_28),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx6p67_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_25),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_23),
.B1(n_27),
.B2(n_19),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_23),
.B1(n_35),
.B2(n_21),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_66),
.B1(n_67),
.B2(n_44),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_28),
.C(n_29),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_43),
.C(n_51),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_57),
.Y(n_73)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_47),
.Y(n_88)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_21),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_69),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_42),
.B(n_29),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_20),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_36),
.Y(n_87)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_83),
.B1(n_87),
.B2(n_78),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_74),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_42),
.B1(n_40),
.B2(n_48),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_63),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_40),
.B1(n_38),
.B2(n_41),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_42),
.B1(n_32),
.B2(n_30),
.Y(n_77)
);

NOR2x1p5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_46),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_70),
.B(n_68),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_50),
.B(n_43),
.C(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_86),
.Y(n_99)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_54),
.C(n_64),
.Y(n_101)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_65),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_95),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_69),
.B1(n_33),
.B2(n_30),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_96),
.B1(n_104),
.B2(n_108),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_60),
.B(n_59),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_54),
.B1(n_64),
.B2(n_40),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_73),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_106),
.C(n_87),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_81),
.B1(n_80),
.B2(n_77),
.Y(n_112)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_109),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_61),
.C(n_41),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_62),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_71),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_88),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_117),
.B1(n_121),
.B2(n_125),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_104),
.A2(n_72),
.B1(n_80),
.B2(n_79),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_113),
.A2(n_127),
.B1(n_38),
.B2(n_105),
.Y(n_148)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_119),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_77),
.B1(n_79),
.B2(n_63),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_130),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_93),
.B(n_109),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_100),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_91),
.B1(n_86),
.B2(n_85),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_110),
.B1(n_101),
.B2(n_103),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_74),
.Y(n_126)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_33),
.B1(n_32),
.B2(n_30),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_131),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_28),
.Y(n_129)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_96),
.Y(n_130)
);

BUFx24_ASAP7_75t_SL g131 ( 
.A(n_106),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_130),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_137),
.Y(n_155)
);

OAI21x1_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_94),
.B(n_106),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_133),
.A2(n_116),
.B1(n_126),
.B2(n_122),
.Y(n_157)
);

XNOR2x1_ASAP7_75t_SL g134 ( 
.A(n_124),
.B(n_108),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_134),
.A2(n_144),
.B(n_153),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_115),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_135),
.B(n_150),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_151),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_108),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_114),
.B(n_97),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_141),
.B(n_111),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_94),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_147),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_26),
.Y(n_166)
);

AO22x2_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_99),
.B1(n_100),
.B2(n_97),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_31),
.B1(n_15),
.B2(n_18),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_99),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_127),
.B1(n_123),
.B2(n_116),
.Y(n_160)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_28),
.B(n_17),
.C(n_62),
.D(n_16),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_113),
.A2(n_38),
.B1(n_33),
.B2(n_32),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_90),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_140),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_158),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_134),
.C(n_149),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_132),
.C(n_142),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_157),
.B(n_14),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

NOR2x1_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_14),
.B(n_1),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_139),
.B(n_18),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_164),
.B(n_174),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_168),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_14),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_144),
.A2(n_45),
.B(n_65),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_171),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_172),
.B(n_173),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_176),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_137),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_167),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_183),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_147),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_166),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_185),
.A2(n_189),
.B(n_160),
.Y(n_198)
);

AO21x2_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_158),
.B(n_157),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_188),
.A2(n_18),
.B1(n_15),
.B2(n_26),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_156),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_SL g218 ( 
.A(n_192),
.B(n_194),
.C(n_196),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_165),
.C(n_170),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_174),
.B1(n_159),
.B2(n_169),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_197),
.A2(n_206),
.B1(n_188),
.B2(n_185),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_145),
.C(n_163),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_203),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_47),
.B1(n_16),
.B2(n_13),
.Y(n_216)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_0),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_90),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_10),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_8),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_188),
.A2(n_18),
.B1(n_15),
.B2(n_31),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_208),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_193),
.A2(n_187),
.B1(n_178),
.B2(n_190),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_178),
.B1(n_184),
.B2(n_45),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_216),
.B1(n_16),
.B2(n_12),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_206),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_0),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_8),
.Y(n_219)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_45),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_214),
.A2(n_205),
.B(n_195),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_217),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_219),
.B(n_220),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_210),
.A2(n_205),
.B1(n_47),
.B2(n_2),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_222),
.B(n_225),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_195),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_228),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_215),
.B(n_12),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_227),
.A2(n_209),
.B(n_212),
.Y(n_231)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_232),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_216),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_218),
.C(n_207),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_236),
.C(n_226),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_12),
.B(n_11),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_235),
.A2(n_9),
.B(n_2),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_11),
.C(n_9),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_239),
.B(n_240),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_47),
.C(n_11),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_1),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_242),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_229),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_SL g245 ( 
.A1(n_240),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_3),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_5),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_244),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g249 ( 
.A(n_248),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_250),
.B1(n_243),
.B2(n_6),
.Y(n_251)
);

OAI221xp5_ASAP7_75t_SL g252 ( 
.A1(n_251),
.A2(n_6),
.B1(n_7),
.B2(n_219),
.C(n_213),
.Y(n_252)
);


endmodule