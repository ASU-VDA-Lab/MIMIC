module fake_jpeg_22736_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_0),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_47),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_51),
.Y(n_79)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_19),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_76),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_33),
.B1(n_31),
.B2(n_17),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_22),
.B1(n_29),
.B2(n_30),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_33),
.B1(n_31),
.B2(n_17),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_33),
.B1(n_31),
.B2(n_17),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_31),
.B1(n_18),
.B2(n_24),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_26),
.B1(n_29),
.B2(n_22),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_29),
.B1(n_18),
.B2(n_24),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_26),
.B1(n_32),
.B2(n_21),
.Y(n_95)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_25),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_41),
.B(n_35),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_83),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_80),
.B(n_89),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_82),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_26),
.B1(n_24),
.B2(n_18),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_86),
.A2(n_95),
.B1(n_107),
.B2(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_28),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_91),
.B(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_32),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_67),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_97),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_63),
.A2(n_16),
.B1(n_21),
.B2(n_32),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_101),
.B1(n_114),
.B2(n_56),
.Y(n_119)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_25),
.B1(n_20),
.B2(n_27),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_55),
.A2(n_28),
.B1(n_27),
.B2(n_21),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_105),
.B1(n_110),
.B2(n_113),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_0),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_106),
.B(n_111),
.Y(n_123)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_58),
.A2(n_28),
.B1(n_25),
.B2(n_20),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_20),
.B(n_1),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_51),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_49),
.A2(n_23),
.B1(n_46),
.B2(n_48),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_0),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_63),
.A2(n_23),
.B1(n_48),
.B2(n_10),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_59),
.A2(n_54),
.B(n_2),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g115 ( 
.A(n_81),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_117),
.B(n_141),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_111),
.Y(n_166)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_108),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_109),
.B1(n_79),
.B2(n_89),
.Y(n_148)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

AOI32xp33_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_53),
.A3(n_54),
.B1(n_40),
.B2(n_44),
.Y(n_129)
);

AOI31xp33_ASAP7_75t_L g165 ( 
.A1(n_129),
.A2(n_83),
.A3(n_111),
.B(n_54),
.Y(n_165)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_90),
.A2(n_53),
.B1(n_75),
.B2(n_44),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_140),
.B1(n_100),
.B2(n_94),
.Y(n_151)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_135),
.A2(n_118),
.B1(n_144),
.B2(n_131),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_90),
.A2(n_37),
.B1(n_40),
.B2(n_23),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_82),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_82),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_142),
.B(n_143),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_146),
.B(n_149),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_148),
.B(n_150),
.Y(n_199)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_151),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_123),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_163),
.Y(n_191)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_158),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_125),
.B1(n_133),
.B2(n_137),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_159),
.B1(n_164),
.B2(n_135),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_139),
.A2(n_92),
.B1(n_85),
.B2(n_98),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_162),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_106),
.B(n_77),
.C(n_103),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_161),
.A2(n_165),
.B(n_166),
.Y(n_185)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_83),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_80),
.B1(n_79),
.B2(n_87),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_93),
.B(n_91),
.Y(n_167)
);

HAxp5_ASAP7_75t_SL g213 ( 
.A(n_167),
.B(n_170),
.CON(n_213),
.SN(n_213)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_127),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_171),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_103),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_175),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_129),
.A2(n_86),
.B(n_87),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_116),
.A2(n_112),
.B(n_78),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_23),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_120),
.B(n_99),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_19),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_119),
.B(n_99),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_128),
.A2(n_101),
.B1(n_84),
.B2(n_54),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_128),
.A2(n_84),
.B1(n_112),
.B2(n_78),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_130),
.A2(n_78),
.B1(n_66),
.B2(n_74),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_130),
.A2(n_13),
.B(n_14),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_88),
.B1(n_10),
.B2(n_3),
.Y(n_204)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_180),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_117),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_184),
.C(n_159),
.Y(n_219)
);

AND2x6_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_143),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_182),
.A2(n_186),
.B(n_6),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_127),
.C(n_142),
.Y(n_184)
);

OA21x2_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_141),
.B(n_124),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_192),
.Y(n_218)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

INVxp67_ASAP7_75t_SL g189 ( 
.A(n_160),
.Y(n_189)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_202),
.B1(n_145),
.B2(n_177),
.Y(n_214)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_193),
.B(n_195),
.Y(n_241)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_196),
.A2(n_200),
.B(n_208),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_162),
.A2(n_138),
.B1(n_144),
.B2(n_118),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_145),
.B1(n_176),
.B2(n_173),
.Y(n_216)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_120),
.B1(n_138),
.B2(n_124),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_204),
.A2(n_210),
.B1(n_169),
.B2(n_172),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_146),
.B(n_59),
.Y(n_207)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_209),
.A2(n_211),
.B(n_161),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_149),
.B(n_37),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_168),
.B(n_1),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_212),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_214),
.A2(n_216),
.B1(n_223),
.B2(n_228),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_201),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_225),
.C(n_232),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_220),
.A2(n_226),
.B(n_238),
.Y(n_264)
);

AOI22x1_ASAP7_75t_SL g222 ( 
.A1(n_186),
.A2(n_166),
.B1(n_163),
.B2(n_172),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_222),
.A2(n_192),
.B1(n_200),
.B2(n_206),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_213),
.A2(n_166),
.B1(n_163),
.B2(n_155),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_74),
.C(n_73),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_185),
.A2(n_19),
.B(n_73),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_19),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_230),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_213),
.A2(n_74),
.B1(n_73),
.B2(n_66),
.Y(n_228)
);

OAI32xp33_ASAP7_75t_L g230 ( 
.A1(n_191),
.A2(n_19),
.A3(n_66),
.B1(n_4),
.B2(n_5),
.Y(n_230)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_182),
.B(n_19),
.C(n_3),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_2),
.C(n_3),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_234),
.C(n_235),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_197),
.B(n_3),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_4),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_191),
.B(n_4),
.C(n_5),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_240),
.C(n_6),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_6),
.C(n_7),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_238),
.A2(n_186),
.B(n_195),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_242),
.A2(n_226),
.B(n_220),
.Y(n_269)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_239),
.Y(n_243)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_245),
.Y(n_279)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_252),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_247),
.A2(n_251),
.B(n_258),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_229),
.B(n_187),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_248),
.B(n_250),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_215),
.B(n_193),
.Y(n_250)
);

OA22x2_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_205),
.B1(n_190),
.B2(n_209),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_207),
.C(n_211),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_218),
.A2(n_196),
.B1(n_202),
.B2(n_199),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_259),
.B1(n_261),
.B2(n_228),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_221),
.B(n_198),
.Y(n_254)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_241),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_255),
.Y(n_272)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_263),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_217),
.A2(n_194),
.B1(n_183),
.B2(n_204),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_232),
.A2(n_194),
.B1(n_188),
.B2(n_180),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_216),
.A2(n_203),
.B1(n_7),
.B2(n_8),
.Y(n_262)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g265 ( 
.A(n_236),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_236),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_264),
.B(n_223),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_268),
.B(n_271),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_269),
.A2(n_247),
.B(n_251),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_219),
.C(n_225),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_274),
.C(n_276),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_235),
.C(n_231),
.Y(n_274)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_234),
.C(n_222),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_237),
.C(n_233),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_282),
.C(n_249),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_227),
.C(n_240),
.Y(n_282)
);

XNOR2x1_ASAP7_75t_L g284 ( 
.A(n_242),
.B(n_7),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_284),
.A2(n_265),
.B1(n_251),
.B2(n_263),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_249),
.B(n_256),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_256),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_253),
.Y(n_287)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_287),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_272),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_292),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_SL g312 ( 
.A(n_289),
.B(n_294),
.C(n_295),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_268),
.Y(n_308)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_296),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_271),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_265),
.C(n_259),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_286),
.C(n_291),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_281),
.B(n_243),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_300),
.B(n_301),
.Y(n_306)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_267),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_304),
.C(n_311),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_274),
.C(n_280),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_314),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_SL g309 ( 
.A(n_294),
.B(n_284),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_309),
.B(n_310),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_295),
.A2(n_283),
.B1(n_262),
.B2(n_278),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_289),
.C(n_297),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_277),
.B(n_278),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_269),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_7),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_251),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_316),
.B(n_324),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_305),
.A2(n_276),
.B1(n_282),
.B2(n_279),
.Y(n_317)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_317),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_315),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_8),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_322),
.B(n_323),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_8),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_8),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_303),
.C(n_311),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_327),
.A2(n_331),
.B(n_321),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_318),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_316),
.B(n_304),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_330),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_308),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_331),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_333),
.B(n_334),
.Y(n_337)
);

NAND4xp25_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_325),
.C(n_320),
.D(n_328),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_338),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_336),
.B1(n_326),
.B2(n_337),
.Y(n_340)
);

O2A1O1Ixp33_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_325),
.B(n_332),
.C(n_9),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_9),
.Y(n_342)
);


endmodule