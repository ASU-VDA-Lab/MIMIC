module fake_netlist_5_2044_n_1639 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_167, n_234, n_343, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1639);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_167;
input n_234;
input n_343;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1639;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_569;
wire n_920;
wire n_1289;
wire n_1517;
wire n_370;
wire n_976;
wire n_1449;
wire n_1566;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_1598;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_696;
wire n_550;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_944;
wire n_1623;
wire n_1565;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1617;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1591;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_1575;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1536;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_325),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_19),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_308),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_61),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_337),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_166),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_200),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_288),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_138),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_40),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_350),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_4),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_120),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_261),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_105),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_272),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_81),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_97),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_236),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_87),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_40),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_109),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_39),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_177),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_118),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_221),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_119),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_224),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_22),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_146),
.Y(n_390)
);

BUFx10_ASAP7_75t_L g391 ( 
.A(n_302),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_233),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_201),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_125),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_163),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_55),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_343),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_240),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_85),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_113),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_297),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_275),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_15),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_9),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_33),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_127),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_46),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_148),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_9),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_278),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_289),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_310),
.Y(n_412)
);

BUFx5_ASAP7_75t_L g413 ( 
.A(n_157),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_347),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_25),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_250),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_154),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_255),
.Y(n_418)
);

BUFx10_ASAP7_75t_L g419 ( 
.A(n_182),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_135),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_53),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_139),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_104),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_22),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_248),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_326),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_341),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_96),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_228),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_295),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_327),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_223),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_173),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_168),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_196),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_239),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_4),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_144),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_50),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_194),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_181),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_359),
.Y(n_442)
);

BUFx10_ASAP7_75t_L g443 ( 
.A(n_206),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_214),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_18),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_286),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_90),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_89),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_185),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_79),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_222),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_211),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_309),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_150),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_191),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_176),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_164),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_218),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_265),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_108),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_210),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_76),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_95),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_111),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_103),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_270),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_123),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_39),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_198),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_266),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_226),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_13),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_209),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_56),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_6),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_305),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_153),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_23),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_212),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_192),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_131),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_0),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_116),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_351),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_23),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_3),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_58),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_189),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_342),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_101),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_60),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_11),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_235),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_152),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_78),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_73),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_20),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_287),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_55),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_26),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_59),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_294),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_75),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_203),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_64),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_358),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_251),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_129),
.Y(n_508)
);

BUFx2_ASAP7_75t_SL g509 ( 
.A(n_324),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_303),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_128),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_300),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_259),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_279),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_322),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_243),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_335),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_312),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_102),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_304),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_171),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_258),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_159),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_328),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_225),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_213),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_290),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_88),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_16),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_338),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_298),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_175),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_117),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_13),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_121),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_149),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_332),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_37),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_59),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_186),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_281),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_215),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_30),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_27),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_241),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_184),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_32),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_315),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_316),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_307),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_254),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_202),
.Y(n_552)
);

INVx1_ASAP7_75t_SL g553 ( 
.A(n_114),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_242),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_15),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_46),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_38),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_249),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_331),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_282),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_37),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_54),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_126),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_165),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_130),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_66),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_348),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_306),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_84),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_293),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_2),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_299),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_7),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_188),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_267),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_141),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_346),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_27),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_208),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_61),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_230),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_205),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_353),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_6),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_363),
.Y(n_585)
);

INVxp33_ASAP7_75t_SL g586 ( 
.A(n_364),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_580),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_580),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_439),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_439),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_375),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_361),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_365),
.Y(n_593)
);

NOR2xp67_ASAP7_75t_L g594 ( 
.A(n_486),
.B(n_0),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_435),
.B(n_1),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_372),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_403),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_381),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_366),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_405),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_415),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_367),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_421),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_437),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_374),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_378),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_474),
.Y(n_607)
);

NOR2xp67_ASAP7_75t_L g608 ( 
.A(n_486),
.B(n_1),
.Y(n_608)
);

BUFx6f_ASAP7_75t_SL g609 ( 
.A(n_391),
.Y(n_609)
);

INVxp67_ASAP7_75t_SL g610 ( 
.A(n_461),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_382),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_482),
.Y(n_612)
);

CKINVDCx16_ASAP7_75t_R g613 ( 
.A(n_377),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_487),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_499),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_384),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_500),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_505),
.Y(n_618)
);

NOR2xp67_ASAP7_75t_L g619 ( 
.A(n_534),
.B(n_2),
.Y(n_619)
);

INVxp67_ASAP7_75t_SL g620 ( 
.A(n_560),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_539),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_386),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_544),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_557),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_369),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_380),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_562),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_571),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_410),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_387),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_390),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_393),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_573),
.Y(n_633)
);

INVxp33_ASAP7_75t_SL g634 ( 
.A(n_362),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_584),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_478),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_375),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_447),
.B(n_477),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_385),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_370),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_385),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_395),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_397),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_398),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_446),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_400),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_446),
.Y(n_647)
);

INVxp33_ASAP7_75t_SL g648 ( 
.A(n_383),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_516),
.B(n_3),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_490),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_411),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_490),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_498),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_389),
.Y(n_654)
);

INVxp33_ASAP7_75t_SL g655 ( 
.A(n_396),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_498),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_561),
.Y(n_657)
);

CKINVDCx16_ASAP7_75t_R g658 ( 
.A(n_401),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_394),
.B(n_5),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_462),
.Y(n_660)
);

NOR2xp67_ASAP7_75t_L g661 ( 
.A(n_426),
.B(n_5),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_462),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_519),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_484),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_519),
.Y(n_665)
);

NOR2xp67_ASAP7_75t_L g666 ( 
.A(n_426),
.B(n_7),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_558),
.B(n_436),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_404),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_414),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_416),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_407),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_563),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_409),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_484),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_514),
.Y(n_675)
);

INVxp33_ASAP7_75t_SL g676 ( 
.A(n_424),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_412),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_R g678 ( 
.A(n_514),
.B(n_527),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_417),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_423),
.Y(n_680)
);

NAND2xp33_ASAP7_75t_R g681 ( 
.A(n_583),
.B(n_427),
.Y(n_681)
);

NOR2xp67_ASAP7_75t_L g682 ( 
.A(n_436),
.B(n_8),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_563),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_579),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_527),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_579),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_458),
.B(n_552),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_428),
.Y(n_688)
);

NOR2xp67_ASAP7_75t_L g689 ( 
.A(n_458),
.B(n_8),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_413),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_429),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_445),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_431),
.Y(n_693)
);

CKINVDCx16_ASAP7_75t_R g694 ( 
.A(n_473),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_552),
.B(n_10),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_368),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_371),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_468),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_R g699 ( 
.A(n_582),
.B(n_432),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_493),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_373),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_376),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_472),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_379),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_433),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_388),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_475),
.Y(n_707)
);

NOR2xp67_ASAP7_75t_L g708 ( 
.A(n_567),
.B(n_11),
.Y(n_708)
);

INVxp33_ASAP7_75t_SL g709 ( 
.A(n_485),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_392),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_567),
.B(n_12),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_434),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_531),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_399),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_554),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_491),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_402),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_438),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_440),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_492),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_406),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_441),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_420),
.Y(n_723)
);

NOR2xp67_ASAP7_75t_L g724 ( 
.A(n_497),
.B(n_12),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_501),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_422),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_444),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_448),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_425),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_413),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_529),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_469),
.B(n_14),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_538),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_413),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_543),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_449),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_430),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_442),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_454),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_589),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_654),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_591),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_696),
.B(n_581),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_590),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_657),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_591),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_697),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_701),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_596),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_702),
.B(n_450),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_668),
.B(n_418),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_586),
.A2(n_638),
.B1(n_595),
.B2(n_613),
.Y(n_752)
);

NAND2xp33_ASAP7_75t_SL g753 ( 
.A(n_678),
.B(n_547),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_704),
.Y(n_754)
);

AND2x2_ASAP7_75t_SL g755 ( 
.A(n_658),
.B(n_408),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_725),
.B(n_391),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_640),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_706),
.B(n_710),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_714),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_694),
.B(n_391),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_717),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_721),
.B(n_451),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_598),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_610),
.B(n_456),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_592),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_732),
.B(n_419),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_723),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_600),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_649),
.B(n_548),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_671),
.B(n_419),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_601),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_726),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_673),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_603),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_604),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_729),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_698),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_620),
.B(n_465),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_661),
.B(n_419),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_607),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_612),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_737),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_614),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_615),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_720),
.B(n_443),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_738),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_617),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_667),
.B(n_553),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_618),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_621),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_623),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_739),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_624),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_627),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_628),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_659),
.B(n_593),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_633),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_637),
.B(n_453),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_635),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_587),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_692),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_707),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_588),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_690),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_639),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_641),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_687),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_690),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_730),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_730),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_645),
.Y(n_811)
);

CKINVDCx8_ASAP7_75t_R g812 ( 
.A(n_599),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_734),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_734),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_647),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_650),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_652),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_653),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_656),
.B(n_555),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_663),
.Y(n_820)
);

INVx4_ASAP7_75t_L g821 ( 
.A(n_602),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_665),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_672),
.B(n_455),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_678),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_683),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_605),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_684),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_686),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_692),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_634),
.B(n_648),
.Y(n_830)
);

CKINVDCx16_ASAP7_75t_R g831 ( 
.A(n_585),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_695),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_666),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_682),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_689),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_708),
.B(n_724),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_711),
.B(n_457),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_619),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_594),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_608),
.B(n_466),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_655),
.B(n_443),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_606),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_736),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_611),
.Y(n_844)
);

INVx4_ASAP7_75t_L g845 ( 
.A(n_843),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_808),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_769),
.A2(n_681),
.B1(n_699),
.B2(n_676),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_755),
.B(n_769),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_804),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_745),
.B(n_616),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_800),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_766),
.B(n_709),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_807),
.B(n_622),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_807),
.B(n_630),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_808),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_808),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_810),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_765),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_810),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_745),
.B(n_631),
.Y(n_860)
);

INVx4_ASAP7_75t_L g861 ( 
.A(n_843),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_741),
.B(n_819),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_741),
.B(n_632),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_788),
.B(n_642),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_807),
.B(n_643),
.Y(n_865)
);

INVxp67_ASAP7_75t_SL g866 ( 
.A(n_746),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_804),
.Y(n_867)
);

OR2x6_ASAP7_75t_L g868 ( 
.A(n_844),
.B(n_509),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_SL g869 ( 
.A(n_812),
.B(n_625),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_742),
.B(n_467),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_803),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_794),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_788),
.B(n_644),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_832),
.B(n_646),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_797),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_814),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_814),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_814),
.Y(n_878)
);

INVx4_ASAP7_75t_SL g879 ( 
.A(n_770),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_832),
.B(n_651),
.Y(n_880)
);

AND2x6_ASAP7_75t_L g881 ( 
.A(n_751),
.B(n_408),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_747),
.Y(n_882)
);

AND2x2_ASAP7_75t_SL g883 ( 
.A(n_824),
.B(n_831),
.Y(n_883)
);

BUFx4f_ASAP7_75t_L g884 ( 
.A(n_832),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_748),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_798),
.B(n_669),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_837),
.B(n_670),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_751),
.B(n_679),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_740),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_764),
.A2(n_778),
.B1(n_837),
.B2(n_840),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_798),
.B(n_680),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_824),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_823),
.B(n_688),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_805),
.B(n_471),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_821),
.B(n_691),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_802),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_744),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_817),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_754),
.Y(n_899)
);

INVxp67_ASAP7_75t_SL g900 ( 
.A(n_817),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_802),
.Y(n_901)
);

INVx1_ASAP7_75t_SL g902 ( 
.A(n_801),
.Y(n_902)
);

OR2x6_ASAP7_75t_L g903 ( 
.A(n_829),
.B(n_479),
.Y(n_903)
);

OR2x6_ASAP7_75t_L g904 ( 
.A(n_760),
.B(n_483),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_809),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_820),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_820),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_826),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_759),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_777),
.B(n_693),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_761),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_767),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_830),
.B(n_705),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_813),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_830),
.B(n_712),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_772),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_820),
.Y(n_917)
);

OR2x6_ASAP7_75t_L g918 ( 
.A(n_842),
.B(n_488),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_768),
.Y(n_919)
);

INVx4_ASAP7_75t_L g920 ( 
.A(n_815),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_785),
.B(n_718),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_776),
.Y(n_922)
);

AND2x6_ASAP7_75t_L g923 ( 
.A(n_756),
.B(n_408),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_782),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_786),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_777),
.B(n_719),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_792),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_828),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_763),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_823),
.B(n_722),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_743),
.B(n_727),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_764),
.A2(n_452),
.B1(n_503),
.B2(n_408),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_806),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_743),
.B(n_728),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_774),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_750),
.B(n_703),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_811),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_768),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_919),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_858),
.Y(n_940)
);

AO22x2_ASAP7_75t_L g941 ( 
.A1(n_848),
.A2(n_841),
.B1(n_779),
.B2(n_778),
.Y(n_941)
);

AO22x2_ASAP7_75t_L g942 ( 
.A1(n_862),
.A2(n_779),
.B1(n_838),
.B2(n_836),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_884),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_884),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_919),
.Y(n_945)
);

AO22x2_ASAP7_75t_L g946 ( 
.A1(n_913),
.A2(n_836),
.B1(n_839),
.B2(n_840),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_852),
.A2(n_796),
.B1(n_753),
.B2(n_752),
.Y(n_947)
);

NOR2xp67_ASAP7_75t_L g948 ( 
.A(n_845),
.B(n_842),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_849),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_916),
.Y(n_950)
);

AO22x2_ASAP7_75t_L g951 ( 
.A1(n_915),
.A2(n_834),
.B1(n_835),
.B2(n_833),
.Y(n_951)
);

AO22x2_ASAP7_75t_L g952 ( 
.A1(n_873),
.A2(n_495),
.B1(n_496),
.B2(n_489),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_919),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_938),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_925),
.Y(n_955)
);

BUFx8_ASAP7_75t_L g956 ( 
.A(n_896),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_860),
.Y(n_957)
);

OAI221xp5_ASAP7_75t_L g958 ( 
.A1(n_890),
.A2(n_762),
.B1(n_750),
.B2(n_758),
.C(n_827),
.Y(n_958)
);

AO22x2_ASAP7_75t_L g959 ( 
.A1(n_850),
.A2(n_520),
.B1(n_522),
.B2(n_510),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_887),
.B(n_716),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_937),
.Y(n_961)
);

NAND2x1p5_ASAP7_75t_L g962 ( 
.A(n_845),
.B(n_816),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_872),
.Y(n_963)
);

NAND2x1p5_ASAP7_75t_L g964 ( 
.A(n_861),
.B(n_825),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_936),
.A2(n_731),
.B1(n_733),
.B2(n_716),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_847),
.A2(n_735),
.B1(n_629),
.B2(n_677),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_861),
.B(n_822),
.Y(n_967)
);

AO22x2_ASAP7_75t_L g968 ( 
.A1(n_864),
.A2(n_526),
.B1(n_530),
.B2(n_525),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_875),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_863),
.B(n_757),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_849),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_867),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_882),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_879),
.B(n_815),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_885),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_920),
.B(n_818),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_917),
.B(n_749),
.Y(n_977)
);

AO22x2_ASAP7_75t_L g978 ( 
.A1(n_902),
.A2(n_568),
.B1(n_569),
.B2(n_546),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_899),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_931),
.A2(n_934),
.B1(n_888),
.B2(n_930),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_909),
.Y(n_981)
);

AO22x2_ASAP7_75t_L g982 ( 
.A1(n_921),
.A2(n_574),
.B1(n_572),
.B2(n_660),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_901),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_866),
.B(n_818),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_867),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_893),
.B(n_757),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_911),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_881),
.A2(n_926),
.B1(n_910),
.B2(n_880),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_881),
.B(n_773),
.Y(n_989)
);

BUFx8_ASAP7_75t_L g990 ( 
.A(n_892),
.Y(n_990)
);

BUFx6f_ASAP7_75t_SL g991 ( 
.A(n_883),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_912),
.Y(n_992)
);

OAI221xp5_ASAP7_75t_L g993 ( 
.A1(n_932),
.A2(n_758),
.B1(n_784),
.B2(n_787),
.C(n_780),
.Y(n_993)
);

OAI221xp5_ASAP7_75t_L g994 ( 
.A1(n_922),
.A2(n_924),
.B1(n_927),
.B2(n_891),
.C(n_886),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_851),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_929),
.B(n_626),
.Y(n_996)
);

AO22x2_ASAP7_75t_L g997 ( 
.A1(n_870),
.A2(n_662),
.B1(n_664),
.B2(n_660),
.Y(n_997)
);

OAI221xp5_ASAP7_75t_L g998 ( 
.A1(n_853),
.A2(n_854),
.B1(n_865),
.B2(n_874),
.C(n_871),
.Y(n_998)
);

CKINVDCx14_ASAP7_75t_R g999 ( 
.A(n_908),
.Y(n_999)
);

NAND2x1p5_ASAP7_75t_L g1000 ( 
.A(n_917),
.B(n_749),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_933),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_935),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_905),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_895),
.B(n_773),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_928),
.B(n_700),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_889),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_897),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_914),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_881),
.B(n_771),
.Y(n_1009)
);

OAI221xp5_ASAP7_75t_L g1010 ( 
.A1(n_904),
.A2(n_790),
.B1(n_789),
.B2(n_799),
.C(n_783),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_846),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_869),
.Y(n_1012)
);

AO22x2_ASAP7_75t_L g1013 ( 
.A1(n_870),
.A2(n_664),
.B1(n_674),
.B2(n_662),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_894),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_894),
.B(n_713),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_881),
.B(n_783),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_900),
.B(n_799),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_923),
.A2(n_715),
.B1(n_459),
.B2(n_463),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_868),
.A2(n_675),
.B1(n_685),
.B2(n_674),
.Y(n_1019)
);

BUFx8_ASAP7_75t_L g1020 ( 
.A(n_938),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_906),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_923),
.A2(n_460),
.B1(n_470),
.B2(n_464),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_846),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_906),
.Y(n_1024)
);

AO22x2_ASAP7_75t_L g1025 ( 
.A1(n_904),
.A2(n_685),
.B1(n_675),
.B2(n_636),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_907),
.Y(n_1026)
);

AO22x2_ASAP7_75t_L g1027 ( 
.A1(n_918),
.A2(n_636),
.B1(n_597),
.B2(n_17),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_907),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_868),
.B(n_775),
.Y(n_1029)
);

AO22x2_ASAP7_75t_L g1030 ( 
.A1(n_918),
.A2(n_597),
.B1(n_609),
.B2(n_17),
.Y(n_1030)
);

AO22x2_ASAP7_75t_L g1031 ( 
.A1(n_903),
.A2(n_609),
.B1(n_18),
.B2(n_14),
.Y(n_1031)
);

AO22x2_ASAP7_75t_L g1032 ( 
.A1(n_903),
.A2(n_20),
.B1(n_16),
.B2(n_19),
.Y(n_1032)
);

AO22x2_ASAP7_75t_L g1033 ( 
.A1(n_857),
.A2(n_25),
.B1(n_21),
.B2(n_24),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_988),
.B(n_938),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_948),
.B(n_898),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_980),
.B(n_923),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_986),
.B(n_957),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_970),
.B(n_947),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_1004),
.B(n_898),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_943),
.B(n_898),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_944),
.B(n_846),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_1012),
.B(n_855),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_989),
.B(n_855),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_974),
.B(n_855),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_967),
.B(n_856),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_960),
.B(n_1029),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_950),
.B(n_878),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_955),
.B(n_856),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_961),
.B(n_859),
.Y(n_1049)
);

NAND2xp33_ASAP7_75t_SL g1050 ( 
.A(n_991),
.B(n_476),
.Y(n_1050)
);

NAND2xp33_ASAP7_75t_SL g1051 ( 
.A(n_940),
.B(n_480),
.Y(n_1051)
);

NAND2xp33_ASAP7_75t_SL g1052 ( 
.A(n_939),
.B(n_481),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_984),
.B(n_877),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_963),
.B(n_876),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_969),
.B(n_876),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_973),
.B(n_975),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_979),
.B(n_775),
.Y(n_1057)
);

NAND2xp33_ASAP7_75t_SL g1058 ( 
.A(n_939),
.B(n_494),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_981),
.B(n_775),
.Y(n_1059)
);

NAND2xp33_ASAP7_75t_SL g1060 ( 
.A(n_945),
.B(n_502),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_987),
.B(n_781),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_992),
.B(n_781),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_1014),
.B(n_795),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_995),
.B(n_781),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_1001),
.B(n_791),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_983),
.B(n_791),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_945),
.B(n_791),
.Y(n_1067)
);

NAND2xp33_ASAP7_75t_SL g1068 ( 
.A(n_1015),
.B(n_504),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_966),
.B(n_793),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_965),
.B(n_793),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_1006),
.B(n_793),
.Y(n_1071)
);

NAND2xp33_ASAP7_75t_SL g1072 ( 
.A(n_1009),
.B(n_506),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_996),
.B(n_795),
.Y(n_1073)
);

NAND2xp33_ASAP7_75t_SL g1074 ( 
.A(n_1016),
.B(n_507),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_1007),
.B(n_795),
.Y(n_1075)
);

NAND2xp33_ASAP7_75t_SL g1076 ( 
.A(n_976),
.B(n_508),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_1018),
.B(n_511),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_1017),
.B(n_512),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_962),
.B(n_513),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_964),
.B(n_515),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_1002),
.B(n_517),
.Y(n_1081)
);

NAND2xp33_ASAP7_75t_SL g1082 ( 
.A(n_1005),
.B(n_518),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_999),
.B(n_578),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_1003),
.B(n_521),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_958),
.B(n_523),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_978),
.B(n_556),
.Y(n_1086)
);

NAND2xp33_ASAP7_75t_SL g1087 ( 
.A(n_1019),
.B(n_524),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_949),
.B(n_528),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_1008),
.B(n_532),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_971),
.B(n_533),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_978),
.B(n_566),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_977),
.B(n_535),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_982),
.B(n_443),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_1000),
.B(n_537),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_972),
.B(n_540),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_985),
.B(n_541),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_1021),
.B(n_542),
.Y(n_1097)
);

NAND2xp33_ASAP7_75t_SL g1098 ( 
.A(n_1024),
.B(n_545),
.Y(n_1098)
);

NAND2xp33_ASAP7_75t_SL g1099 ( 
.A(n_1026),
.B(n_1028),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_1022),
.B(n_549),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_982),
.B(n_942),
.Y(n_1101)
);

NAND2xp33_ASAP7_75t_SL g1102 ( 
.A(n_953),
.B(n_550),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_998),
.B(n_551),
.Y(n_1103)
);

NAND2xp33_ASAP7_75t_SL g1104 ( 
.A(n_954),
.B(n_559),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_1011),
.B(n_452),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_1023),
.B(n_452),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_1020),
.B(n_564),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_990),
.B(n_565),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_942),
.B(n_570),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_951),
.B(n_71),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_956),
.B(n_575),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_946),
.B(n_576),
.Y(n_1112)
);

NAND2xp33_ASAP7_75t_SL g1113 ( 
.A(n_941),
.B(n_577),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1047),
.Y(n_1114)
);

CKINVDCx16_ASAP7_75t_R g1115 ( 
.A(n_1083),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1053),
.A2(n_946),
.B(n_951),
.Y(n_1116)
);

NAND2x1p5_ASAP7_75t_L g1117 ( 
.A(n_1073),
.B(n_452),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1038),
.A2(n_994),
.B1(n_941),
.B2(n_968),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1036),
.A2(n_993),
.B(n_1010),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1037),
.B(n_959),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1056),
.Y(n_1121)
);

NOR2x1_ASAP7_75t_SL g1122 ( 
.A(n_1034),
.B(n_503),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1085),
.A2(n_959),
.B(n_952),
.C(n_503),
.Y(n_1123)
);

OR2x6_ASAP7_75t_L g1124 ( 
.A(n_1110),
.B(n_1013),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_1110),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1046),
.B(n_952),
.Y(n_1126)
);

AO21x2_ASAP7_75t_L g1127 ( 
.A1(n_1109),
.A2(n_1033),
.B(n_413),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_1075),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_1051),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_1075),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_1063),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1063),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_1070),
.Y(n_1133)
);

O2A1O1Ixp5_ASAP7_75t_SL g1134 ( 
.A1(n_1039),
.A2(n_1031),
.B(n_1032),
.C(n_1030),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1101),
.B(n_1027),
.Y(n_1135)
);

NOR2x1p5_ASAP7_75t_L g1136 ( 
.A(n_1093),
.B(n_1013),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1103),
.A2(n_413),
.B(n_536),
.Y(n_1137)
);

AO31x2_ASAP7_75t_L g1138 ( 
.A1(n_1112),
.A2(n_536),
.A3(n_1025),
.B(n_1027),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_1086),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_1044),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_1091),
.Y(n_1141)
);

AO31x2_ASAP7_75t_L g1142 ( 
.A1(n_1059),
.A2(n_1025),
.A3(n_997),
.B(n_26),
.Y(n_1142)
);

AOI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1043),
.A2(n_74),
.B(n_72),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1048),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1113),
.A2(n_21),
.B(n_24),
.C(n_28),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1042),
.B(n_28),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1069),
.A2(n_178),
.B1(n_357),
.B2(n_356),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1088),
.B(n_29),
.Y(n_1148)
);

O2A1O1Ixp5_ASAP7_75t_L g1149 ( 
.A1(n_1078),
.A2(n_174),
.B(n_355),
.C(n_354),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1105),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1105),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1090),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_1099),
.A2(n_29),
.A3(n_30),
.B(n_31),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_1045),
.B(n_77),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1052),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_1072),
.Y(n_1156)
);

INVxp67_ASAP7_75t_SL g1157 ( 
.A(n_1066),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1035),
.A2(n_82),
.B(n_80),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1106),
.Y(n_1159)
);

INVx3_ASAP7_75t_SL g1160 ( 
.A(n_1108),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1087),
.B(n_31),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1077),
.A2(n_1100),
.B(n_1096),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_SL g1163 ( 
.A1(n_1074),
.A2(n_86),
.B(n_83),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1040),
.B(n_33),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1106),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1095),
.A2(n_92),
.B(n_91),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_1076),
.A2(n_34),
.A3(n_35),
.B(n_36),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1049),
.A2(n_94),
.B(n_93),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1092),
.A2(n_99),
.B(n_98),
.Y(n_1169)
);

NAND2xp33_ASAP7_75t_L g1170 ( 
.A(n_1094),
.B(n_100),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1054),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1055),
.A2(n_107),
.B(n_106),
.Y(n_1172)
);

AO21x2_ASAP7_75t_L g1173 ( 
.A1(n_1097),
.A2(n_112),
.B(n_110),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1071),
.A2(n_122),
.B(n_115),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_SL g1175 ( 
.A1(n_1107),
.A2(n_34),
.B(n_36),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1041),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1081),
.A2(n_219),
.B(n_352),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1067),
.B(n_124),
.Y(n_1178)
);

NOR2xp67_ASAP7_75t_L g1179 ( 
.A(n_1079),
.B(n_1080),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1057),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_1061),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1114),
.B(n_1062),
.Y(n_1182)
);

CKINVDCx6p67_ASAP7_75t_R g1183 ( 
.A(n_1160),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1131),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_1137),
.A2(n_1065),
.B(n_1064),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1125),
.A2(n_1084),
.B1(n_1089),
.B2(n_1111),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1133),
.B(n_1050),
.Y(n_1187)
);

AND2x2_ASAP7_75t_SL g1188 ( 
.A(n_1161),
.B(n_1068),
.Y(n_1188)
);

INVx1_ASAP7_75t_SL g1189 ( 
.A(n_1139),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1152),
.B(n_1082),
.Y(n_1190)
);

OA21x2_ASAP7_75t_L g1191 ( 
.A1(n_1116),
.A2(n_1098),
.B(n_1102),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1121),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1131),
.Y(n_1193)
);

INVx6_ASAP7_75t_SL g1194 ( 
.A(n_1124),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1118),
.A2(n_1104),
.B1(n_1060),
.B2(n_1058),
.Y(n_1195)
);

INVx4_ASAP7_75t_SL g1196 ( 
.A(n_1153),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1141),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1145),
.A2(n_38),
.B(n_41),
.C(n_42),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1152),
.B(n_41),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1171),
.Y(n_1200)
);

OR2x6_ASAP7_75t_L g1201 ( 
.A(n_1131),
.B(n_132),
.Y(n_1201)
);

OR2x2_ASAP7_75t_L g1202 ( 
.A(n_1135),
.B(n_42),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1132),
.B(n_43),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1168),
.A2(n_227),
.B(n_349),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1132),
.B(n_43),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_SL g1206 ( 
.A1(n_1124),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1115),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1162),
.A2(n_229),
.B(n_345),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1128),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1128),
.B(n_44),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1126),
.B(n_45),
.Y(n_1211)
);

OA21x2_ASAP7_75t_L g1212 ( 
.A1(n_1119),
.A2(n_231),
.B(n_344),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1171),
.Y(n_1213)
);

OAI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1120),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1157),
.B(n_48),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1138),
.B(n_49),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1150),
.Y(n_1217)
);

AO21x2_ASAP7_75t_L g1218 ( 
.A1(n_1122),
.A2(n_232),
.B(n_340),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1150),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1151),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1148),
.A2(n_220),
.B(n_339),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1172),
.A2(n_217),
.B(n_336),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1151),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1140),
.Y(n_1224)
);

NOR2x1_ASAP7_75t_L g1225 ( 
.A(n_1179),
.B(n_133),
.Y(n_1225)
);

NAND4xp25_ASAP7_75t_L g1226 ( 
.A(n_1146),
.B(n_50),
.C(n_51),
.D(n_52),
.Y(n_1226)
);

AOI221xp5_ASAP7_75t_L g1227 ( 
.A1(n_1175),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.C(n_54),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1143),
.A2(n_238),
.B(n_334),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1130),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1130),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1140),
.Y(n_1231)
);

AO22x1_ASAP7_75t_L g1232 ( 
.A1(n_1154),
.A2(n_1129),
.B1(n_1155),
.B2(n_1178),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1170),
.A2(n_244),
.B(n_333),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1123),
.A2(n_57),
.B(n_60),
.C(n_62),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1138),
.B(n_62),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1176),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1144),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_SL g1238 ( 
.A1(n_1177),
.A2(n_246),
.B(n_330),
.C(n_329),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1176),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_1164),
.Y(n_1240)
);

NOR2xp67_ASAP7_75t_L g1241 ( 
.A(n_1156),
.B(n_134),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1166),
.A2(n_245),
.B(n_323),
.Y(n_1242)
);

NAND2x1p5_ASAP7_75t_L g1243 ( 
.A(n_1140),
.B(n_136),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1138),
.B(n_63),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1154),
.B(n_360),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1181),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1159),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1181),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1181),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1159),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1180),
.B(n_137),
.Y(n_1251)
);

OR2x6_ASAP7_75t_L g1252 ( 
.A(n_1178),
.B(n_140),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1165),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1165),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1234),
.A2(n_1169),
.A3(n_1158),
.B(n_1153),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1217),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1217),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1200),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1219),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_1183),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1240),
.B(n_1156),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1232),
.B(n_1134),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1213),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1224),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1192),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1246),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1219),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1216),
.B(n_1127),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1220),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1197),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1220),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1237),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1207),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1223),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1223),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1247),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1188),
.A2(n_1136),
.B1(n_1117),
.B2(n_1147),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1186),
.A2(n_1127),
.B1(n_1173),
.B2(n_1174),
.Y(n_1278)
);

INVx4_ASAP7_75t_SL g1279 ( 
.A(n_1201),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1245),
.B(n_1173),
.Y(n_1280)
);

AND2x4_ASAP7_75t_SL g1281 ( 
.A(n_1251),
.B(n_1163),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1235),
.B(n_1153),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1244),
.B(n_1167),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1193),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1247),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1250),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1250),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1254),
.B(n_1142),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1254),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1242),
.A2(n_1149),
.B(n_256),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1239),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1203),
.Y(n_1292)
);

AO21x2_ASAP7_75t_L g1293 ( 
.A1(n_1221),
.A2(n_1167),
.B(n_1142),
.Y(n_1293)
);

AO21x1_ASAP7_75t_L g1294 ( 
.A1(n_1198),
.A2(n_1167),
.B(n_1142),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1246),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1204),
.A2(n_252),
.B(n_320),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1211),
.B(n_1245),
.Y(n_1297)
);

INVxp67_ASAP7_75t_SL g1298 ( 
.A(n_1231),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1187),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_1299)
);

OAI21xp33_ASAP7_75t_L g1300 ( 
.A1(n_1227),
.A2(n_68),
.B(n_69),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1205),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1246),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1212),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1196),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1189),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1212),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1190),
.B(n_142),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1252),
.B(n_321),
.Y(n_1308)
);

BUFx12f_ASAP7_75t_L g1309 ( 
.A(n_1202),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1228),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1222),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1252),
.B(n_257),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1251),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1199),
.B(n_70),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1210),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1208),
.A2(n_253),
.B(n_143),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1182),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1209),
.Y(n_1318)
);

O2A1O1Ixp33_ASAP7_75t_SL g1319 ( 
.A1(n_1214),
.A2(n_70),
.B(n_145),
.C(n_147),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1229),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1195),
.A2(n_151),
.B(n_155),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1248),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1191),
.A2(n_156),
.B(n_158),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1248),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1201),
.B(n_1196),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1249),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1231),
.Y(n_1327)
);

INVxp67_ASAP7_75t_L g1328 ( 
.A(n_1273),
.Y(n_1328)
);

NAND2xp33_ASAP7_75t_R g1329 ( 
.A(n_1305),
.B(n_1249),
.Y(n_1329)
);

XOR2xp5_ASAP7_75t_L g1330 ( 
.A(n_1260),
.B(n_1243),
.Y(n_1330)
);

XNOR2xp5_ASAP7_75t_L g1331 ( 
.A(n_1260),
.B(n_1226),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1297),
.B(n_1268),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1317),
.B(n_1215),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_R g1334 ( 
.A(n_1305),
.B(n_1184),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1297),
.B(n_1206),
.Y(n_1335)
);

XOR2xp5_ASAP7_75t_L g1336 ( 
.A(n_1313),
.B(n_1225),
.Y(n_1336)
);

OR2x6_ASAP7_75t_L g1337 ( 
.A(n_1325),
.B(n_1241),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1291),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_R g1339 ( 
.A(n_1313),
.B(n_1184),
.Y(n_1339)
);

NAND2xp33_ASAP7_75t_R g1340 ( 
.A(n_1308),
.B(n_1191),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1279),
.B(n_1218),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1274),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1268),
.B(n_1236),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1279),
.B(n_1233),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1292),
.B(n_1253),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1276),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1301),
.B(n_1230),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1285),
.Y(n_1348)
);

NAND2xp33_ASAP7_75t_R g1349 ( 
.A(n_1308),
.B(n_1185),
.Y(n_1349)
);

OR2x6_ASAP7_75t_L g1350 ( 
.A(n_1325),
.B(n_1194),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1315),
.B(n_1238),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1270),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1261),
.B(n_1185),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1291),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1256),
.Y(n_1355)
);

NAND2xp33_ASAP7_75t_R g1356 ( 
.A(n_1312),
.B(n_1194),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1314),
.B(n_1272),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1286),
.Y(n_1358)
);

NAND2xp33_ASAP7_75t_R g1359 ( 
.A(n_1312),
.B(n_160),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1279),
.B(n_161),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1256),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_R g1362 ( 
.A(n_1313),
.B(n_162),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_R g1363 ( 
.A(n_1313),
.B(n_319),
.Y(n_1363)
);

XNOR2xp5_ASAP7_75t_L g1364 ( 
.A(n_1270),
.B(n_167),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_1264),
.Y(n_1365)
);

XOR2xp5_ASAP7_75t_L g1366 ( 
.A(n_1277),
.B(n_169),
.Y(n_1366)
);

INVxp33_ASAP7_75t_L g1367 ( 
.A(n_1284),
.Y(n_1367)
);

NAND2xp33_ASAP7_75t_R g1368 ( 
.A(n_1304),
.B(n_170),
.Y(n_1368)
);

NAND2xp33_ASAP7_75t_R g1369 ( 
.A(n_1304),
.B(n_172),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_R g1370 ( 
.A(n_1309),
.B(n_179),
.Y(n_1370)
);

BUFx10_ASAP7_75t_L g1371 ( 
.A(n_1295),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_R g1372 ( 
.A(n_1309),
.B(n_318),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1314),
.B(n_180),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1257),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_R g1375 ( 
.A(n_1266),
.B(n_317),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1279),
.B(n_183),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_SL g1377 ( 
.A(n_1307),
.B(n_187),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1265),
.B(n_190),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1257),
.Y(n_1379)
);

INVxp67_ASAP7_75t_L g1380 ( 
.A(n_1302),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_R g1381 ( 
.A(n_1266),
.B(n_314),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1298),
.B(n_193),
.Y(n_1382)
);

INVxp67_ASAP7_75t_L g1383 ( 
.A(n_1295),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_R g1384 ( 
.A(n_1295),
.B(n_1327),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1259),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1283),
.B(n_195),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_R g1387 ( 
.A(n_1295),
.B(n_197),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_R g1388 ( 
.A(n_1327),
.B(n_313),
.Y(n_1388)
);

XOR2xp5_ASAP7_75t_L g1389 ( 
.A(n_1280),
.B(n_199),
.Y(n_1389)
);

NAND2xp33_ASAP7_75t_R g1390 ( 
.A(n_1280),
.B(n_204),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_R g1391 ( 
.A(n_1262),
.B(n_207),
.Y(n_1391)
);

NAND2xp33_ASAP7_75t_R g1392 ( 
.A(n_1280),
.B(n_1283),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_R g1393 ( 
.A(n_1322),
.B(n_311),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1324),
.B(n_216),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1258),
.B(n_1263),
.Y(n_1395)
);

NAND2xp33_ASAP7_75t_R g1396 ( 
.A(n_1282),
.B(n_234),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1318),
.B(n_237),
.Y(n_1397)
);

NAND2xp33_ASAP7_75t_R g1398 ( 
.A(n_1282),
.B(n_247),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1326),
.B(n_260),
.Y(n_1399)
);

BUFx10_ASAP7_75t_L g1400 ( 
.A(n_1281),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1353),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1332),
.B(n_1293),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1366),
.A2(n_1300),
.B1(n_1321),
.B2(n_1299),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1342),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1361),
.B(n_1259),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_SL g1406 ( 
.A(n_1391),
.B(n_1281),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1346),
.B(n_1293),
.Y(n_1407)
);

OAI222xp33_ASAP7_75t_L g1408 ( 
.A1(n_1389),
.A2(n_1278),
.B1(n_1288),
.B2(n_1320),
.C1(n_1318),
.C2(n_1290),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1348),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1358),
.B(n_1293),
.Y(n_1410)
);

INVxp67_ASAP7_75t_SL g1411 ( 
.A(n_1355),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1374),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1379),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1343),
.B(n_1288),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1385),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1395),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1386),
.B(n_1338),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1341),
.B(n_1289),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1354),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1341),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1357),
.B(n_1289),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1335),
.B(n_1275),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1380),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1351),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1333),
.B(n_1294),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1331),
.A2(n_1294),
.B1(n_1316),
.B2(n_1320),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1378),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1400),
.Y(n_1428)
);

INVxp67_ASAP7_75t_SL g1429 ( 
.A(n_1349),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1347),
.B(n_1287),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1345),
.B(n_1287),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1367),
.B(n_1275),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1400),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1344),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1344),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1373),
.B(n_1271),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1397),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1371),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1371),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1383),
.Y(n_1440)
);

INVxp67_ASAP7_75t_SL g1441 ( 
.A(n_1392),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1337),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1364),
.B(n_1271),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1337),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1365),
.B(n_1267),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1399),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1399),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1360),
.B(n_1267),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1360),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1382),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1377),
.A2(n_1316),
.B1(n_1310),
.B2(n_1311),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1376),
.B(n_1269),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1336),
.B(n_1269),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1382),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1394),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1442),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1426),
.A2(n_1323),
.B(n_1303),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1404),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1401),
.Y(n_1459)
);

NAND2x1p5_ASAP7_75t_SL g1460 ( 
.A(n_1406),
.B(n_1398),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1402),
.B(n_1306),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1432),
.B(n_1328),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1404),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1402),
.B(n_1306),
.Y(n_1464)
);

AOI221xp5_ASAP7_75t_L g1465 ( 
.A1(n_1455),
.A2(n_1319),
.B1(n_1372),
.B2(n_1370),
.C(n_1393),
.Y(n_1465)
);

AOI33xp33_ASAP7_75t_L g1466 ( 
.A1(n_1403),
.A2(n_1455),
.A3(n_1319),
.B1(n_1427),
.B2(n_1416),
.B3(n_1432),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1412),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1418),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1414),
.B(n_1303),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1425),
.B(n_1255),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1442),
.A2(n_1376),
.B1(n_1363),
.B2(n_1362),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1414),
.B(n_1255),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1425),
.B(n_1407),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1421),
.B(n_1352),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1407),
.B(n_1255),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1418),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1409),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1412),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1444),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1412),
.Y(n_1480)
);

AOI221xp5_ASAP7_75t_L g1481 ( 
.A1(n_1408),
.A2(n_1388),
.B1(n_1381),
.B2(n_1375),
.C(n_1330),
.Y(n_1481)
);

OAI33xp33_ASAP7_75t_L g1482 ( 
.A1(n_1427),
.A2(n_1396),
.A3(n_1359),
.B1(n_1329),
.B2(n_1368),
.B3(n_1369),
.Y(n_1482)
);

OAI221xp5_ASAP7_75t_L g1483 ( 
.A1(n_1444),
.A2(n_1390),
.B1(n_1356),
.B2(n_1340),
.C(n_1350),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1409),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1421),
.B(n_1334),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1424),
.Y(n_1486)
);

AOI211xp5_ASAP7_75t_L g1487 ( 
.A1(n_1429),
.A2(n_1387),
.B(n_1339),
.C(n_1384),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1441),
.A2(n_1350),
.B1(n_1310),
.B2(n_1311),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1458),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1463),
.Y(n_1490)
);

NAND2x1p5_ASAP7_75t_L g1491 ( 
.A(n_1457),
.B(n_1449),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1477),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1459),
.B(n_1420),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1484),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1467),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1468),
.B(n_1420),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1467),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1482),
.B(n_1453),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1468),
.B(n_1434),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1486),
.B(n_1453),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1468),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1478),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1456),
.B(n_1435),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1478),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1480),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1480),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1485),
.B(n_1423),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1473),
.Y(n_1508)
);

NAND4xp25_ASAP7_75t_L g1509 ( 
.A(n_1466),
.B(n_1443),
.C(n_1436),
.D(n_1431),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1479),
.B(n_1434),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1473),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1476),
.B(n_1435),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1462),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1500),
.B(n_1474),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1500),
.B(n_1445),
.Y(n_1515)
);

NAND2xp33_ASAP7_75t_SL g1516 ( 
.A(n_1493),
.B(n_1466),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1513),
.B(n_1445),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1489),
.Y(n_1518)
);

OAI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1509),
.A2(n_1481),
.B1(n_1465),
.B2(n_1483),
.C(n_1471),
.Y(n_1519)
);

CKINVDCx20_ASAP7_75t_R g1520 ( 
.A(n_1507),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1490),
.Y(n_1521)
);

INVxp33_ASAP7_75t_SL g1522 ( 
.A(n_1507),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1511),
.B(n_1508),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1498),
.B(n_1461),
.Y(n_1524)
);

NAND2xp33_ASAP7_75t_SL g1525 ( 
.A(n_1503),
.B(n_1460),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1498),
.B(n_1416),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1508),
.B(n_1476),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1499),
.B(n_1487),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1491),
.A2(n_1460),
.B1(n_1446),
.B2(n_1450),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1492),
.B(n_1494),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1510),
.B(n_1464),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1512),
.B(n_1461),
.Y(n_1532)
);

NAND2x1_ASAP7_75t_L g1533 ( 
.A(n_1496),
.B(n_1476),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1499),
.B(n_1472),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1527),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1518),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1533),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1521),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1523),
.B(n_1501),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1530),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1517),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1528),
.B(n_1499),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1524),
.Y(n_1543)
);

INVxp67_ASAP7_75t_SL g1544 ( 
.A(n_1522),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1526),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1525),
.A2(n_1449),
.B1(n_1454),
.B2(n_1447),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1531),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1534),
.B(n_1470),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1526),
.B(n_1496),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1520),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1532),
.B(n_1496),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1515),
.B(n_1470),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_1516),
.Y(n_1553)
);

OAI32xp33_ASAP7_75t_L g1554 ( 
.A1(n_1553),
.A2(n_1519),
.A3(n_1491),
.B1(n_1514),
.B2(n_1475),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_SL g1555 ( 
.A1(n_1544),
.A2(n_1449),
.B1(n_1450),
.B2(n_1454),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1545),
.B(n_1529),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1543),
.A2(n_1529),
.B1(n_1449),
.B2(n_1457),
.Y(n_1557)
);

OAI21xp33_ASAP7_75t_SL g1558 ( 
.A1(n_1537),
.A2(n_1506),
.B(n_1497),
.Y(n_1558)
);

AOI221xp5_ASAP7_75t_L g1559 ( 
.A1(n_1540),
.A2(n_1488),
.B1(n_1504),
.B2(n_1502),
.C(n_1495),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1550),
.B(n_1428),
.Y(n_1560)
);

NAND4xp25_ASAP7_75t_L g1561 ( 
.A(n_1546),
.B(n_1436),
.C(n_1446),
.D(n_1431),
.Y(n_1561)
);

OAI211xp5_ASAP7_75t_SL g1562 ( 
.A1(n_1540),
.A2(n_1451),
.B(n_1440),
.C(n_1430),
.Y(n_1562)
);

OAI221xp5_ASAP7_75t_SL g1563 ( 
.A1(n_1549),
.A2(n_1475),
.B1(n_1454),
.B2(n_1447),
.C(n_1464),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1560),
.B(n_1547),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1556),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1559),
.B(n_1547),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1561),
.B(n_1536),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1555),
.B(n_1541),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1557),
.A2(n_1542),
.B1(n_1537),
.B2(n_1535),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1563),
.B(n_1552),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1562),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1558),
.A2(n_1542),
.B1(n_1535),
.B2(n_1551),
.Y(n_1572)
);

BUFx2_ASAP7_75t_L g1573 ( 
.A(n_1564),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1567),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1572),
.B(n_1542),
.Y(n_1575)
);

INVxp33_ASAP7_75t_SL g1576 ( 
.A(n_1565),
.Y(n_1576)
);

INVx8_ASAP7_75t_L g1577 ( 
.A(n_1566),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1571),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_1568),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1569),
.Y(n_1580)
);

NAND4xp25_ASAP7_75t_L g1581 ( 
.A(n_1580),
.B(n_1554),
.C(n_1570),
.D(n_1538),
.Y(n_1581)
);

NOR4xp75_ASAP7_75t_L g1582 ( 
.A(n_1575),
.B(n_1576),
.C(n_1577),
.D(n_1579),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1573),
.Y(n_1583)
);

NAND4xp25_ASAP7_75t_L g1584 ( 
.A(n_1574),
.B(n_1578),
.C(n_1577),
.D(n_1538),
.Y(n_1584)
);

AOI31xp33_ASAP7_75t_L g1585 ( 
.A1(n_1577),
.A2(n_1551),
.A3(n_1539),
.B(n_1552),
.Y(n_1585)
);

NOR3xp33_ASAP7_75t_L g1586 ( 
.A(n_1579),
.B(n_1428),
.C(n_1433),
.Y(n_1586)
);

NOR3xp33_ASAP7_75t_L g1587 ( 
.A(n_1579),
.B(n_1428),
.C(n_1433),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1577),
.B(n_1539),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1581),
.A2(n_1548),
.B1(n_1433),
.B2(n_1440),
.Y(n_1589)
);

AOI222xp33_ASAP7_75t_L g1590 ( 
.A1(n_1583),
.A2(n_1437),
.B1(n_1472),
.B2(n_1422),
.C1(n_1410),
.C2(n_1447),
.Y(n_1590)
);

AOI211xp5_ASAP7_75t_SL g1591 ( 
.A1(n_1585),
.A2(n_1548),
.B(n_1438),
.C(n_1439),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1588),
.A2(n_1505),
.B1(n_1430),
.B2(n_1422),
.Y(n_1592)
);

NAND4xp25_ASAP7_75t_L g1593 ( 
.A(n_1584),
.B(n_1437),
.C(n_1417),
.D(n_1439),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1593),
.Y(n_1594)
);

NAND3xp33_ASAP7_75t_L g1595 ( 
.A(n_1591),
.B(n_1587),
.C(n_1586),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1589),
.Y(n_1596)
);

NOR2x1_ASAP7_75t_L g1597 ( 
.A(n_1592),
.B(n_1582),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1590),
.A2(n_1457),
.B1(n_1437),
.B2(n_1452),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1589),
.B(n_1438),
.Y(n_1599)
);

XNOR2xp5_ASAP7_75t_L g1600 ( 
.A(n_1597),
.B(n_1452),
.Y(n_1600)
);

NAND3xp33_ASAP7_75t_L g1601 ( 
.A(n_1595),
.B(n_1439),
.C(n_1438),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_R g1602 ( 
.A(n_1596),
.B(n_262),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1594),
.B(n_1505),
.Y(n_1603)
);

NAND2xp33_ASAP7_75t_SL g1604 ( 
.A(n_1599),
.B(n_1448),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1598),
.B(n_1469),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_R g1606 ( 
.A(n_1596),
.B(n_263),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_R g1607 ( 
.A(n_1596),
.B(n_264),
.Y(n_1607)
);

OAI22x1_ASAP7_75t_L g1608 ( 
.A1(n_1600),
.A2(n_1448),
.B1(n_1418),
.B2(n_1417),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1601),
.A2(n_1415),
.B1(n_1413),
.B2(n_1411),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1602),
.B(n_1415),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1603),
.Y(n_1611)
);

BUFx2_ASAP7_75t_SL g1612 ( 
.A(n_1606),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1607),
.B(n_1469),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1604),
.A2(n_1296),
.B(n_1323),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1605),
.A2(n_1418),
.B1(n_1413),
.B2(n_1410),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1605),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1611),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1612),
.B(n_1405),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1610),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1616),
.B(n_1405),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1613),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1615),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1608),
.A2(n_1419),
.B1(n_1405),
.B2(n_1311),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1617),
.A2(n_1609),
.B1(n_1614),
.B2(n_1419),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1620),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1625),
.A2(n_1622),
.B1(n_1621),
.B2(n_1619),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1624),
.A2(n_1618),
.B1(n_1623),
.B2(n_1419),
.Y(n_1627)
);

AOI31xp33_ASAP7_75t_L g1628 ( 
.A1(n_1625),
.A2(n_268),
.A3(n_269),
.B(n_271),
.Y(n_1628)
);

NOR3xp33_ASAP7_75t_L g1629 ( 
.A(n_1628),
.B(n_1296),
.C(n_274),
.Y(n_1629)
);

OR5x1_ASAP7_75t_L g1630 ( 
.A(n_1626),
.B(n_273),
.C(n_276),
.D(n_277),
.E(n_280),
.Y(n_1630)
);

XNOR2xp5_ASAP7_75t_L g1631 ( 
.A(n_1627),
.B(n_283),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1630),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1631),
.B(n_284),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1629),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1633),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1632),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1634),
.Y(n_1637)
);

OAI221xp5_ASAP7_75t_R g1638 ( 
.A1(n_1636),
.A2(n_285),
.B1(n_291),
.B2(n_292),
.C(n_296),
.Y(n_1638)
);

AOI211xp5_ASAP7_75t_L g1639 ( 
.A1(n_1638),
.A2(n_1637),
.B(n_1635),
.C(n_301),
.Y(n_1639)
);


endmodule