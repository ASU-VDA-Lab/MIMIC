module fake_jpeg_23197_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_42),
.Y(n_60)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_29),
.B1(n_25),
.B2(n_19),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_29),
.B1(n_25),
.B2(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_62),
.Y(n_66)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_63),
.B(n_88),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_64),
.A2(n_72),
.B1(n_78),
.B2(n_86),
.Y(n_124)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_67),
.Y(n_96)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

OR2x4_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_30),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_79),
.B(n_35),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_71),
.B(n_35),
.Y(n_118)
);

AO22x1_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_16),
.B1(n_30),
.B2(n_40),
.Y(n_72)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_73),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_42),
.Y(n_94)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_80),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_61),
.A2(n_29),
.B1(n_19),
.B2(n_18),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_42),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_89),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_10),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_16),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_44),
.Y(n_84)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_18),
.B1(n_30),
.B2(n_24),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_18),
.B1(n_44),
.B2(n_39),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_59),
.B(n_49),
.C(n_55),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_58),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_36),
.Y(n_91)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_36),
.Y(n_93)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_94),
.B(n_119),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_36),
.C(n_39),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_66),
.C(n_80),
.Y(n_132)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_109),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_88),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_101),
.Y(n_135)
);

AND2x4_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_30),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_107),
.B(n_92),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_103),
.B(n_111),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_79),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_105),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_72),
.B(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_73),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_121),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_40),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_118),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_59),
.B1(n_49),
.B2(n_16),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_71),
.B1(n_107),
.B2(n_102),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_39),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_122),
.A2(n_76),
.B1(n_67),
.B2(n_57),
.Y(n_134)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_65),
.Y(n_131)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_137),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_126),
.A2(n_140),
.B1(n_110),
.B2(n_104),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_113),
.C(n_114),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_120),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_133),
.A2(n_123),
.B1(n_69),
.B2(n_108),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_69),
.B1(n_75),
.B2(n_116),
.Y(n_153)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_138),
.A2(n_142),
.B(n_147),
.Y(n_178)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_144),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_119),
.A2(n_109),
.B1(n_112),
.B2(n_95),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_90),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_141),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_105),
.A2(n_28),
.B(n_26),
.C(n_32),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_80),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_149),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_124),
.A2(n_21),
.B(n_31),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_99),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_151),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_153),
.A2(n_166),
.B1(n_173),
.B2(n_183),
.Y(n_205)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_164),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_163),
.A2(n_184),
.B(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_169),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_118),
.Y(n_167)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_114),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_168),
.B(n_32),
.Y(n_207)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_174),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_111),
.B(n_118),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_136),
.B(n_133),
.Y(n_198)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_108),
.C(n_106),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_177),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_106),
.B1(n_75),
.B2(n_100),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_146),
.B1(n_89),
.B2(n_135),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_40),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_129),
.Y(n_179)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_135),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_180),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_97),
.C(n_43),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_41),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_126),
.A2(n_97),
.B1(n_121),
.B2(n_82),
.Y(n_183)
);

AND2x4_ASAP7_75t_L g184 ( 
.A(n_125),
.B(n_43),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_161),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_186),
.B(n_217),
.Y(n_233)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_140),
.A3(n_148),
.B1(n_130),
.B2(n_125),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_187),
.B(n_194),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_162),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_189),
.Y(n_224)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_196),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_197),
.C(n_175),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_184),
.A2(n_130),
.B(n_139),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_192),
.A2(n_208),
.B(n_28),
.Y(n_237)
);

OAI32xp33_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_139),
.A3(n_136),
.B1(n_142),
.B2(n_137),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_28),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_209),
.B1(n_210),
.B2(n_181),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_166),
.A2(n_149),
.B1(n_146),
.B2(n_70),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_200),
.A2(n_212),
.B1(n_215),
.B2(n_169),
.Y(n_218)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_202),
.Y(n_221)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_154),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_207),
.B(n_160),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_172),
.A2(n_20),
.B(n_22),
.Y(n_208)
);

OAI22x1_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_129),
.B1(n_70),
.B2(n_31),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_165),
.A2(n_26),
.B1(n_22),
.B2(n_27),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_0),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_156),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_183),
.A2(n_34),
.B1(n_31),
.B2(n_21),
.Y(n_212)
);

CKINVDCx12_ASAP7_75t_R g213 ( 
.A(n_154),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_216),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_178),
.A2(n_34),
.B1(n_41),
.B2(n_43),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_155),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_218),
.A2(n_216),
.B1(n_214),
.B2(n_203),
.Y(n_257)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_177),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_238),
.Y(n_246)
);

HAxp5_ASAP7_75t_SL g250 ( 
.A(n_222),
.B(n_211),
.CON(n_250),
.SN(n_250)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_205),
.A2(n_158),
.B1(n_178),
.B2(n_163),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_223),
.A2(n_192),
.B1(n_204),
.B2(n_209),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_226),
.C(n_227),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_155),
.C(n_164),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_174),
.C(n_171),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_191),
.B(n_158),
.C(n_43),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_198),
.C(n_215),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_214),
.Y(n_258)
);

AOI21xp33_ASAP7_75t_L g234 ( 
.A1(n_188),
.A2(n_10),
.B(n_14),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_234),
.B(n_210),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_185),
.B(n_9),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_243),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_208),
.B(n_211),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_187),
.B(n_41),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_41),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_9),
.Y(n_241)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_206),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_232),
.A2(n_217),
.B1(n_204),
.B2(n_200),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_244),
.A2(n_250),
.B1(n_258),
.B2(n_261),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_247),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_225),
.C(n_239),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_195),
.Y(n_253)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_254),
.Y(n_282)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_237),
.B(n_222),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_194),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_256),
.Y(n_267)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_221),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_230),
.A2(n_201),
.B1(n_31),
.B2(n_21),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_218),
.A2(n_17),
.B1(n_1),
.B2(n_3),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_220),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_247),
.B(n_223),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_270),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_274),
.C(n_276),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_233),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_275),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_244),
.A2(n_242),
.B1(n_227),
.B2(n_240),
.Y(n_269)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

XOR2x2_ASAP7_75t_SL g272 ( 
.A(n_256),
.B(n_250),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_272),
.Y(n_283)
);

XOR2x2_ASAP7_75t_SL g273 ( 
.A(n_256),
.B(n_242),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_273),
.B(n_277),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_226),
.C(n_238),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_222),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_28),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_28),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_8),
.Y(n_281)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_285),
.A2(n_272),
.B1(n_265),
.B2(n_282),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_278),
.B(n_249),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_286),
.Y(n_308)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_270),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_276),
.B(n_264),
.Y(n_290)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_258),
.C(n_263),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_295),
.C(n_8),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_262),
.C(n_255),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_248),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_0),
.Y(n_303)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_298),
.Y(n_311)
);

AOI21x1_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_280),
.B(n_266),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_285),
.B1(n_297),
.B2(n_294),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_254),
.C(n_259),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_304),
.Y(n_310)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_28),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_306),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_8),
.C(n_14),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_7),
.C(n_14),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_309),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_7),
.C(n_12),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_312),
.B(n_313),
.Y(n_321)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g314 ( 
.A1(n_298),
.A2(n_283),
.B(n_292),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_314),
.A2(n_284),
.B(n_288),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_319),
.A2(n_320),
.B(n_323),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_308),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_304),
.C(n_300),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_322),
.B(n_324),
.Y(n_329)
);

OAI31xp33_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_292),
.A3(n_293),
.B(n_4),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_6),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_17),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_325),
.A2(n_17),
.B1(n_5),
.B2(n_6),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_321),
.A2(n_317),
.B1(n_318),
.B2(n_4),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_326),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_328),
.B(n_5),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_326),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_329),
.B(n_327),
.Y(n_333)
);

AOI322xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_331),
.A3(n_321),
.B1(n_6),
.B2(n_9),
.C1(n_11),
.C2(n_3),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_11),
.C(n_1),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_11),
.C(n_3),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_3),
.Y(n_337)
);


endmodule