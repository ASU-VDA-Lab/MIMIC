module fake_jpeg_28592_n_90 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_90);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_90;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_1),
.Y(n_51)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_27),
.Y(n_50)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_33),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_51),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_57),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_25),
.B(n_6),
.C(n_7),
.Y(n_56)
);

AO21x2_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_8),
.B(n_9),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_5),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_12),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_59),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_65),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_69),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_68),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_42),
.B1(n_14),
.B2(n_15),
.Y(n_70)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_71),
.B(n_72),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_13),
.B(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_74),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_24),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_78),
.A2(n_67),
.B(n_21),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_80),
.Y(n_83)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_75),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_85),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_82),
.B1(n_81),
.B2(n_77),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g89 ( 
.A1(n_88),
.A2(n_79),
.B(n_74),
.C(n_73),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_62),
.Y(n_90)
);


endmodule