module real_jpeg_30836_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_0),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_0),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_1),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_1),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_1),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_1),
.B(n_348),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_1),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_1),
.B(n_391),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_2),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_2),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_2),
.B(n_135),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_2),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_2),
.B(n_185),
.Y(n_184)
);

NAND2xp33_ASAP7_75t_SL g205 ( 
.A(n_2),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_2),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_2),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_3),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_3),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_3),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_3),
.B(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_3),
.Y(n_167)
);

NAND2x1_ASAP7_75t_L g304 ( 
.A(n_3),
.B(n_81),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_3),
.B(n_350),
.Y(n_349)
);

NAND2x1_ASAP7_75t_L g406 ( 
.A(n_3),
.B(n_407),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_4),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_4),
.Y(n_280)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_6),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_6),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_6),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_6),
.B(n_300),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_6),
.B(n_300),
.Y(n_305)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_6),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_6),
.B(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_7),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_7),
.Y(n_165)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_7),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_8),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_8),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_8),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_8),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_8),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_8),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_8),
.B(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_9),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_9),
.Y(n_189)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_9),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_10),
.Y(n_389)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_11),
.Y(n_105)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_11),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_12),
.B(n_88),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_12),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_12),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_12),
.B(n_415),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_13),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_13),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_14),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_14),
.B(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_14),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_14),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_14),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_14),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_14),
.B(n_332),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_15),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_15),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_15),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_15),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_15),
.B(n_336),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_15),
.B(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_364),
.Y(n_16)
);

NOR2xp67_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_360),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_252),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_154),
.B(n_251),
.Y(n_19)
);

NOR2xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_108),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_21),
.B(n_108),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_69),
.C(n_90),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_22),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_23),
.B(n_52),
.C(n_67),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_24)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_25),
.B(n_34),
.C(n_35),
.Y(n_115)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_28),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_39),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_52),
.B1(n_67),
.B2(n_68),
.Y(n_40)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_42),
.B(n_47),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_42),
.A2(n_43),
.B1(n_92),
.B2(n_93),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

MAJx2_ASAP7_75t_L g380 ( 
.A(n_43),
.B(n_93),
.C(n_322),
.Y(n_380)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_51),
.Y(n_135)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_51),
.Y(n_266)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_51),
.Y(n_351)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.C(n_62),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_53),
.B(n_62),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_57),
.Y(n_338)
);

XNOR2x2_ASAP7_75t_SL g239 ( 
.A(n_58),
.B(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_65),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_66),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_66),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_69),
.A2(n_70),
.B1(n_90),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_79),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_71),
.B(n_84),
.C(n_89),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

AO22x1_ASAP7_75t_SL g106 ( 
.A1(n_72),
.A2(n_76),
.B1(n_77),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_72),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_72),
.A2(n_107),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_72),
.B(n_278),
.C(n_282),
.Y(n_354)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_74),
.Y(n_169)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22x1_ASAP7_75t_L g419 ( 
.A1(n_76),
.A2(n_77),
.B1(n_420),
.B2(n_422),
.Y(n_419)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_84),
.B1(n_85),
.B2(n_89),
.Y(n_79)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_90),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_99),
.C(n_106),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_91),
.B(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_92),
.A2(n_93),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_93),
.B(n_95),
.Y(n_181)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_98),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_99),
.A2(n_100),
.B1(n_106),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_104),
.Y(n_218)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_104),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_105),
.Y(n_199)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_105),
.Y(n_272)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_106),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_130),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_110),
.B(n_130),
.C(n_255),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_111),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_117),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2x1_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_114),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_115),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_116),
.B(n_259),
.C(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_127),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_SL g289 ( 
.A(n_119),
.B(n_123),
.C(n_127),
.Y(n_289)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_126),
.Y(n_348)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_131),
.B(n_138),
.C(n_152),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_138),
.B1(n_152),
.B2(n_153),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_136),
.B(n_137),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_136),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_137),
.B(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_137),
.B(n_267),
.C(n_273),
.Y(n_344)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

XNOR2x1_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_145),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_140),
.B(n_148),
.C(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx6_ASAP7_75t_L g333 ( 
.A(n_144),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_146),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_146),
.B(n_404),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_150),
.B(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21x1_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_245),
.B(n_250),
.Y(n_154)
);

OAI21x1_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_233),
.B(n_244),
.Y(n_155)
);

AOI21x1_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_202),
.B(n_232),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_176),
.Y(n_157)
);

NOR2x1_ASAP7_75t_L g232 ( 
.A(n_158),
.B(n_176),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_170),
.C(n_173),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_159),
.A2(n_160),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_166),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_166),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_170),
.A2(n_173),
.B1(n_174),
.B2(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_170),
.Y(n_212)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_182),
.B1(n_200),
.B2(n_201),
.Y(n_176)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_178),
.B(n_181),
.C(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_184),
.B(n_191),
.C(n_195),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.Y(n_190)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

OAI21x1_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_213),
.B(n_231),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_209),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_207),
.Y(n_215)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_219),
.B(n_230),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_216),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_224),
.Y(n_297)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_236),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_239),
.C(n_241),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

NOR2xp67_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_249),
.Y(n_250)
);

NOR2x1_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_308),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g362 ( 
.A(n_254),
.B(n_256),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_285),
.Y(n_256)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_257),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_261),
.Y(n_257)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_258),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_274),
.Y(n_261)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_262),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_267),
.B1(n_268),
.B2(n_273),
.Y(n_263)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_264),
.Y(n_273)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_274),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_281),
.B2(n_284),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_280),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_306),
.B2(n_307),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_287),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_292),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_289),
.B(n_290),
.C(n_293),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_298),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_294),
.B(n_304),
.C(n_340),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_303),
.B1(n_304),
.B2(n_305),
.Y(n_298)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx5_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_302),
.Y(n_418)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_310),
.C(n_311),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_308),
.A2(n_362),
.B(n_363),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_312),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_309),
.B(n_312),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_317),
.Y(n_312)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_313),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.C(n_316),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_341),
.B1(n_342),
.B2(n_356),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_339),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_326),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_320),
.B(n_357),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_320),
.B(n_326),
.C(n_359),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_325),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_326),
.A2(n_339),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_326),
.Y(n_358)
);

XOR2x2_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_335),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_330),
.B1(n_331),
.B2(n_334),
.Y(n_327)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_328),
.Y(n_334)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_331),
.Y(n_412)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_334),
.B(n_335),
.C(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_337),
.Y(n_421)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_339),
.Y(n_359)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_342),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_355),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

HB1xp67_ASAP7_75t_SL g399 ( 
.A(n_344),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_345),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_354),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_349),
.B1(n_352),
.B2(n_353),
.Y(n_346)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_347),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_349),
.Y(n_353)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_353),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_354),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_355),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_356),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_423),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_371),
.Y(n_366)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_367),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.C(n_370),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_371),
.Y(n_426)
);

XNOR2x1_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_396),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_393),
.B1(n_394),
.B2(n_395),
.Y(n_373)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_374),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_379),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.C(n_378),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_386),
.B1(n_390),
.B2(n_392),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_384),
.Y(n_391)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_386),
.Y(n_392)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

XNOR2x1_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_401),
.Y(n_396)
);

MAJx2_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.C(n_400),
.Y(n_397)
);

XOR2x2_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_410),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_413),
.Y(n_410)
);

XNOR2x1_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_419),
.Y(n_413)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_420),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);


endmodule