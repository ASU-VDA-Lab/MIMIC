module fake_jpeg_756_n_374 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_374);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_374;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_51),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_52),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_53),
.B(n_64),
.Y(n_126)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_54),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_16),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_56),
.A2(n_69),
.B(n_90),
.C(n_91),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_72),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g119 ( 
.A(n_60),
.Y(n_119)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_0),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_65),
.Y(n_147)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_26),
.B(n_0),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_25),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_77),
.Y(n_104)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g150 ( 
.A(n_76),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_25),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_26),
.B(n_2),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_80),
.B(n_4),
.Y(n_143)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_36),
.Y(n_84)
);

BUFx8_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_32),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_34),
.B(n_2),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_34),
.B(n_2),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_42),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_42),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_30),
.Y(n_137)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_41),
.B(n_43),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_101),
.A2(n_6),
.B(n_10),
.C(n_11),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_61),
.B1(n_76),
.B2(n_62),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_110),
.A2(n_159),
.B1(n_73),
.B2(n_55),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_60),
.A2(n_43),
.B1(n_41),
.B2(n_44),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_124),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_68),
.A2(n_45),
.B1(n_44),
.B2(n_46),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_52),
.A2(n_45),
.B1(n_46),
.B2(n_27),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_52),
.A2(n_24),
.B1(n_30),
.B2(n_27),
.Y(n_124)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_129),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_137),
.B(n_143),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_56),
.B(n_36),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_144),
.Y(n_162)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_51),
.A2(n_36),
.B1(n_33),
.B2(n_28),
.Y(n_146)
);

AO22x1_ASAP7_75t_SL g163 ( 
.A1(n_146),
.A2(n_96),
.B1(n_89),
.B2(n_82),
.Y(n_163)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_79),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_78),
.B(n_5),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_149),
.B(n_6),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_55),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_132),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_168),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_174),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_164),
.Y(n_233)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_165),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_166),
.B(n_167),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_73),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_132),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_106),
.B(n_59),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_169),
.B(n_116),
.C(n_131),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_119),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_176),
.Y(n_216)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_103),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_126),
.B(n_10),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_177),
.B(n_184),
.Y(n_234)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_103),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_198),
.Y(n_223)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_181),
.Y(n_235)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_118),
.B(n_11),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_183),
.B(n_195),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_104),
.B(n_128),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_153),
.A2(n_104),
.B(n_127),
.C(n_134),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_113),
.B(n_159),
.C(n_116),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_109),
.B(n_111),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_187),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_130),
.B(n_158),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_188),
.A2(n_190),
.B1(n_121),
.B2(n_107),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_125),
.A2(n_147),
.B1(n_105),
.B2(n_155),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_114),
.B(n_152),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_191),
.B(n_202),
.Y(n_214)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_193),
.Y(n_213)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_141),
.B(n_123),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_120),
.B(n_147),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_196),
.B(n_162),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_156),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_200),
.Y(n_228)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_136),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_170),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_115),
.B(n_108),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_124),
.B(n_146),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_203),
.B(n_202),
.Y(n_227)
);

OR2x2_ASAP7_75t_SL g240 ( 
.A(n_205),
.B(n_180),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_184),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_217),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_203),
.A2(n_133),
.B1(n_151),
.B2(n_131),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_218),
.A2(n_231),
.B1(n_182),
.B2(n_193),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_189),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_219),
.B(n_224),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_174),
.A2(n_138),
.B(n_154),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_220),
.A2(n_227),
.B(n_169),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_121),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_191),
.A2(n_163),
.B1(n_185),
.B2(n_187),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_228),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_236),
.B(n_243),
.Y(n_282)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_237),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_227),
.A2(n_163),
.B1(n_180),
.B2(n_197),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_252),
.B1(n_256),
.B2(n_218),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_240),
.A2(n_246),
.B1(n_211),
.B2(n_209),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_212),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_241),
.B(n_247),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_224),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_228),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_216),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_248),
.Y(n_262)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_213),
.Y(n_249)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_249),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_192),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_250),
.B(n_253),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_214),
.A2(n_180),
.B(n_175),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_205),
.B(n_211),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_180),
.B1(n_199),
.B2(n_178),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_165),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_213),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_254),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_214),
.A2(n_173),
.B1(n_188),
.B2(n_172),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_204),
.B(n_169),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_258),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_219),
.B(n_200),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_210),
.B(n_201),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_259),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_206),
.Y(n_260)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_204),
.B(n_201),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_217),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_263),
.A2(n_238),
.B(n_254),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_264),
.A2(n_245),
.B1(n_260),
.B2(n_206),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_232),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_270),
.Y(n_289)
);

OAI32xp33_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_209),
.A3(n_208),
.B1(n_233),
.B2(n_223),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_283),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_251),
.A2(n_220),
.B(n_235),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_274),
.A2(n_284),
.B(n_230),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_233),
.C(n_222),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_258),
.C(n_255),
.Y(n_295)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_242),
.B(n_209),
.CI(n_234),
.CON(n_278),
.SN(n_278)
);

A2O1A1O1Ixp25_ASAP7_75t_L g296 ( 
.A1(n_278),
.A2(n_243),
.B(n_236),
.C(n_234),
.D(n_255),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_261),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_248),
.Y(n_285)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_281),
.Y(n_287)
);

AO22x1_ASAP7_75t_SL g283 ( 
.A1(n_246),
.A2(n_239),
.B1(n_240),
.B2(n_256),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_252),
.A2(n_235),
.B(n_222),
.Y(n_284)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

OA21x2_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_237),
.B(n_253),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_286),
.A2(n_291),
.B(n_296),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_262),
.B(n_247),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_288),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_244),
.Y(n_290)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_290),
.Y(n_318)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_293),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_238),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_297),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_304),
.C(n_294),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_213),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_298),
.B(n_272),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_299),
.A2(n_287),
.B1(n_293),
.B2(n_245),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_282),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_300),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_229),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_301),
.A2(n_303),
.B1(n_277),
.B2(n_276),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_302),
.A2(n_263),
.B1(n_271),
.B2(n_284),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_282),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_232),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_306),
.A2(n_286),
.B(n_291),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_289),
.A2(n_283),
.B1(n_269),
.B2(n_264),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_317),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_320),
.C(n_321),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_295),
.Y(n_323)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_315),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_289),
.A2(n_281),
.B1(n_269),
.B2(n_245),
.Y(n_316)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_316),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_283),
.B1(n_275),
.B2(n_270),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_319),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_278),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_278),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_292),
.A2(n_280),
.B1(n_260),
.B2(n_230),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_322),
.B(n_310),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_323),
.B(n_312),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_324),
.A2(n_319),
.B(n_313),
.Y(n_346)
);

BUFx12_ASAP7_75t_L g326 ( 
.A(n_312),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_329),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_327),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_309),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_292),
.Y(n_330)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_330),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_314),
.A2(n_296),
.B(n_299),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_333),
.Y(n_340)
);

NOR2xp67_ASAP7_75t_SL g333 ( 
.A(n_314),
.B(n_297),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_286),
.C(n_287),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_323),
.C(n_311),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_337),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_336),
.C(n_335),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_334),
.A2(n_317),
.B1(n_307),
.B2(n_306),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_343),
.B(n_344),
.Y(n_347)
);

FAx1_ASAP7_75t_SL g344 ( 
.A(n_324),
.B(n_320),
.CI(n_321),
.CON(n_344),
.SN(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_318),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_345),
.B(n_346),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_342),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_349),
.B(n_350),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_339),
.B(n_310),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_352),
.B(n_353),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_338),
.B(n_335),
.C(n_325),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_340),
.B(n_325),
.C(n_328),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_354),
.B(n_328),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_347),
.B(n_346),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_356),
.B(n_360),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_357),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_348),
.A2(n_341),
.B1(n_343),
.B2(n_344),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_359),
.B(n_360),
.C(n_358),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_347),
.B(n_337),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_351),
.B(n_280),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_361),
.B(n_226),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_363),
.B(n_365),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_356),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_366),
.B(n_365),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_364),
.B(n_355),
.C(n_344),
.Y(n_368)
);

O2A1O1Ixp33_ASAP7_75t_SL g370 ( 
.A1(n_368),
.A2(n_367),
.B(n_362),
.C(n_326),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_369),
.A2(n_326),
.B1(n_230),
.B2(n_226),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_370),
.B(n_371),
.C(n_181),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_372),
.A2(n_207),
.B(n_314),
.Y(n_373)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_373),
.Y(n_374)
);


endmodule