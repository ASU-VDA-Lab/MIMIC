module real_jpeg_4592_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g97 ( 
.A(n_0),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_1),
.A2(n_42),
.B1(n_104),
.B2(n_107),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_1),
.A2(n_42),
.B1(n_175),
.B2(n_178),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_1),
.A2(n_42),
.B1(n_203),
.B2(n_207),
.Y(n_202)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_2),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_2),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_2),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_3),
.A2(n_156),
.B1(n_157),
.B2(n_160),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_3),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_3),
.A2(n_156),
.B1(n_236),
.B2(n_238),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_3),
.A2(n_156),
.B1(n_280),
.B2(n_283),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_3),
.A2(n_156),
.B1(n_417),
.B2(n_418),
.Y(n_416)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_4),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_5),
.Y(n_166)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_5),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_5),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_5),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_6),
.Y(n_147)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_9),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_10),
.A2(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_11),
.Y(n_120)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_11),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_11),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_12),
.A2(n_26),
.B1(n_95),
.B2(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_12),
.B(n_31),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_12),
.A2(n_26),
.B1(n_130),
.B2(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_12),
.A2(n_26),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_12),
.A2(n_303),
.B(n_305),
.C(n_313),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_12),
.B(n_329),
.C(n_331),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_12),
.B(n_111),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_12),
.B(n_166),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_12),
.B(n_127),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_13),
.A2(n_41),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_13),
.A2(n_68),
.B1(n_104),
.B2(n_107),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_13),
.A2(n_68),
.B1(n_139),
.B2(n_309),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_13),
.A2(n_68),
.B1(n_339),
.B2(n_343),
.Y(n_338)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_442),
.Y(n_20)
);

OAI221xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_53),
.B1(n_57),
.B2(n_437),
.C(n_440),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_22),
.B(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_22),
.B(n_53),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_23),
.B(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_24),
.B(n_213),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_44),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_28),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_26),
.B(n_29),
.Y(n_28)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_26),
.A2(n_306),
.B(n_309),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_28),
.Y(n_151)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2x1_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_31),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_31),
.B(n_40),
.Y(n_212)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_34),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_35),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_37),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_39),
.B(n_66),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_39),
.A2(n_55),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_44),
.B(n_67),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g152 ( 
.A(n_49),
.B(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_53),
.A2(n_262),
.B1(n_265),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_53),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_53),
.A2(n_265),
.B(n_271),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B(n_56),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_54),
.A2(n_212),
.B(n_416),
.Y(n_433)
);

A2O1A1O1Ixp25_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_395),
.B(n_427),
.C(n_430),
.D(n_436),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_387),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_250),
.C(n_292),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_222),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_194),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_62),
.B(n_194),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_141),
.C(n_179),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_63),
.B(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_73),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_64),
.B(n_74),
.C(n_113),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_65),
.B(n_212),
.Y(n_402)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_71),
.Y(n_417)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_112),
.B1(n_113),
.B2(n_140),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_109),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_76),
.A2(n_111),
.B(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_76),
.B(n_216),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_102),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_77),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_89),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_84),
.B2(n_86),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_80),
.Y(n_304)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_86),
.Y(n_283)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_89),
.B(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_93),
.B1(n_98),
.B2(n_100),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_92),
.Y(n_308)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_96),
.Y(n_206)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_96),
.Y(n_241)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_97),
.Y(n_312)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_99),
.Y(n_237)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_103),
.B(n_111),
.Y(n_181)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_106),
.Y(n_221)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_106),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_108),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_109),
.B(n_260),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_110),
.B(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_111),
.A2(n_183),
.B(n_218),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_112),
.A2(n_113),
.B1(n_422),
.B2(n_423),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_112),
.B(n_402),
.C(n_405),
.Y(n_425)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_113),
.B(n_405),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_113),
.B(n_423),
.C(n_424),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_135),
.B(n_136),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_114),
.A2(n_201),
.B(n_235),
.Y(n_264)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_115),
.B(n_137),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_115),
.B(n_202),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_115),
.B(n_319),
.Y(n_318)
);

NOR2x1_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_127),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_119),
.B1(n_121),
.B2(n_124),
.Y(n_116)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AO22x1_ASAP7_75t_SL g127 ( 
.A1(n_120),
.A2(n_128),
.B1(n_130),
.B2(n_133),
.Y(n_127)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_123),
.Y(n_330)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_126),
.Y(n_207)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_127),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_127),
.B(n_319),
.Y(n_333)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_128),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g331 ( 
.A(n_132),
.Y(n_331)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_135),
.A2(n_235),
.B(n_242),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_135),
.B(n_136),
.Y(n_285)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_141),
.A2(n_142),
.B1(n_179),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_154),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_143),
.B(n_154),
.Y(n_209)
);

AOI32xp33_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.A3(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_150),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_164),
.B(n_167),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_155),
.A2(n_191),
.B(n_198),
.Y(n_197)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_166),
.Y(n_356)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_168),
.A2(n_188),
.B(n_230),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_168),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_169),
.Y(n_361)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_170),
.Y(n_342)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_179),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.C(n_186),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_180),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_181),
.B(n_260),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_181),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_183),
.B(n_218),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_183),
.A2(n_279),
.B(n_406),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_186),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_187),
.B(n_355),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_191),
.B(n_337),
.Y(n_365)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_194),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_194),
.B(n_223),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_196),
.CI(n_208),
.CON(n_194),
.SN(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_199),
.Y(n_244)
);

AND2x2_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_200),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_201),
.B(n_318),
.Y(n_345)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_206),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_211),
.C(n_214),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_222),
.A2(n_390),
.B(n_391),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_224),
.B(n_226),
.C(n_243),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_243),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_234),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_234),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_233),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_228),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_233),
.B(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_242),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_242),
.B(n_333),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_247),
.C(n_248),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_246),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_246),
.B(n_433),
.C(n_434),
.Y(n_439)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_248),
.B(n_433),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_289),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_251),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_267),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_252),
.B(n_267),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_261),
.C(n_266),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_253),
.B(n_261),
.CI(n_266),
.CON(n_290),
.SN(n_290)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_258),
.C(n_259),
.Y(n_288)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_262),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_264),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_262),
.B(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_262),
.A2(n_265),
.B1(n_302),
.B2(n_378),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_288),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_276),
.B2(n_277),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_270),
.B(n_276),
.C(n_288),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_284),
.B(n_287),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_278),
.B(n_284),
.Y(n_287)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_285),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_287),
.A2(n_399),
.B1(n_400),
.B2(n_407),
.Y(n_398)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_287),
.Y(n_407)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_289),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_290),
.B(n_291),
.Y(n_392)
);

BUFx24_ASAP7_75t_SL g444 ( 
.A(n_290),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_320),
.B(n_386),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_297),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_294),
.B(n_297),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.C(n_315),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_298),
.B(n_382),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_301),
.A2(n_315),
.B1(n_316),
.B2(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_301),
.Y(n_383)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_302),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_380),
.B(n_385),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_370),
.B(n_379),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_349),
.B(n_369),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_334),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_324),
.B(n_334),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_332),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_325),
.A2(n_326),
.B1(n_332),
.B2(n_352),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_332),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_344),
.Y(n_334)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_335),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_338),
.B(n_356),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_345),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.Y(n_344)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_345),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_346),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_346),
.B(n_347),
.C(n_372),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_350),
.A2(n_357),
.B(n_368),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_353),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_353),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_364),
.B(n_367),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_363),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_362),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_365),
.B(n_366),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_373),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_373),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_377),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_376),
.C(n_377),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_384),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_381),
.B(n_384),
.Y(n_385)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g387 ( 
.A1(n_388),
.A2(n_389),
.B(n_392),
.C(n_393),
.D(n_394),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_410),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_409),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_397),
.B(n_409),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_408),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_407),
.C(n_408),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_402),
.B1(n_403),
.B2(n_404),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_401),
.A2(n_402),
.B1(n_413),
.B2(n_414),
.Y(n_412)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_402),
.B(n_413),
.C(n_425),
.Y(n_435)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_410),
.A2(n_428),
.B(n_429),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_426),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_426),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_425),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_420),
.B1(n_421),
.B2(n_424),
.Y(n_414)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_415),
.Y(n_424)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_435),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_431),
.B(n_435),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_434),
.Y(n_431)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_439),
.Y(n_441)
);


endmodule