module fake_jpeg_13390_n_147 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_147);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_SL g36 ( 
.A(n_27),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_5),
.B(n_28),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_1),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_1),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_68),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_2),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_72),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_73),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_83),
.Y(n_86)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_63),
.B(n_47),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_46),
.C(n_39),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_60),
.B(n_53),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_87),
.B(n_89),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_48),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_93),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_59),
.B1(n_40),
.B2(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_37),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_42),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_24),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_53),
.B1(n_36),
.B2(n_52),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_53),
.B1(n_41),
.B2(n_60),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_102),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_112)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_2),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_110),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_38),
.C(n_58),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_10),
.C(n_12),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_88),
.B(n_3),
.Y(n_110)
);

FAx1_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_4),
.CI(n_5),
.CON(n_111),
.SN(n_111)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_114),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_8),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_118),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_96),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_119),
.B(n_120),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_8),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_130),
.C(n_129),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_22),
.C(n_23),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_108),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_117),
.B(n_111),
.C(n_112),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_109),
.B(n_30),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_134),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_127),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_133),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_116),
.C(n_113),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_135),
.A2(n_122),
.B(n_31),
.Y(n_137)
);

A2O1A1O1Ixp25_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_123),
.B(n_129),
.C(n_125),
.D(n_126),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_137),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_138),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_131),
.C(n_139),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_140),
.Y(n_147)
);


endmodule