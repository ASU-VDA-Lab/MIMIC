module fake_ariane_2932_n_44 (n_8, n_3, n_2, n_7, n_5, n_1, n_0, n_6, n_4, n_44);

input n_8;
input n_3;
input n_2;
input n_7;
input n_5;
input n_1;
input n_0;
input n_6;
input n_4;

output n_44;

wire n_24;
wire n_22;
wire n_43;
wire n_13;
wire n_27;
wire n_20;
wire n_29;
wire n_17;
wire n_41;
wire n_38;
wire n_18;
wire n_32;
wire n_28;
wire n_37;
wire n_9;
wire n_11;
wire n_34;
wire n_26;
wire n_14;
wire n_36;
wire n_33;
wire n_19;
wire n_30;
wire n_39;
wire n_40;
wire n_31;
wire n_42;
wire n_16;
wire n_12;
wire n_15;
wire n_21;
wire n_23;
wire n_35;
wire n_10;
wire n_25;

CKINVDCx5p33_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_0),
.B(n_8),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_1),
.Y(n_13)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_1),
.Y(n_16)
);

AND2x2_ASAP7_75t_SL g17 ( 
.A(n_13),
.B(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_R g20 ( 
.A(n_9),
.B(n_15),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

OR2x6_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_2),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_17),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_17),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

AOI21xp33_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_23),
.B(n_10),
.Y(n_28)
);

OAI221xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_23),
.B1(n_18),
.B2(n_16),
.C(n_27),
.Y(n_29)
);

OAI221xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_16),
.B1(n_22),
.B2(n_19),
.C(n_12),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_12),
.B1(n_21),
.B2(n_20),
.Y(n_31)
);

AO21x2_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_20),
.B(n_12),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_4),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_12),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_32),
.B(n_31),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_SL g38 ( 
.A1(n_33),
.A2(n_35),
.B(n_36),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_38),
.B(n_25),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_36),
.B1(n_32),
.B2(n_7),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_4),
.Y(n_42)
);

NOR2xp67_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_5),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_8),
.B1(n_41),
.B2(n_10),
.Y(n_44)
);


endmodule