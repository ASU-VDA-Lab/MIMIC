module fake_jpeg_31022_n_147 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_147);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_45),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_25),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_0),
.B(n_1),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_50),
.C(n_59),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_69),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_74),
.Y(n_80)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_64),
.B1(n_63),
.B2(n_55),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_79),
.B1(n_64),
.B2(n_74),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_66),
.B1(n_65),
.B2(n_53),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_74),
.A2(n_61),
.B1(n_54),
.B2(n_55),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_62),
.B(n_4),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_60),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_88),
.B(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_58),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_104),
.B1(n_18),
.B2(n_21),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_0),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_99),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_97),
.B(n_106),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_2),
.Y(n_99)
);

NAND2x1_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_5),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_87),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_101),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_26),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_7),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_105),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_12),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_13),
.B(n_16),
.C(n_17),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_112),
.B1(n_109),
.B2(n_118),
.Y(n_131)
);

AO22x1_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_115),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_122),
.Y(n_134)
);

AOI22x1_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_102),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_117),
.B(n_42),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_43),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_106),
.A2(n_34),
.B(n_35),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_36),
.B(n_38),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_128),
.B(n_130),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_41),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_129),
.B(n_112),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_123),
.B(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_111),
.B(n_116),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_133),
.B1(n_121),
.B2(n_114),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_121),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_135),
.Y(n_140)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_134),
.B(n_126),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_137),
.Y(n_142)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_143),
.B(n_140),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_138),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_139),
.C(n_141),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_127),
.Y(n_147)
);


endmodule