module fake_netlist_6_4945_n_798 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_798);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_798;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_772;
wire n_656;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_127),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_29),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_8),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_5),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_7),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_89),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_125),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_98),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_52),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_48),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_149),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_116),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_96),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_31),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_22),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_132),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_121),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_110),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_126),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_55),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_97),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_26),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_2),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_64),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_92),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_73),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_79),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_35),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_74),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_20),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_44),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_37),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_3),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_123),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_148),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_101),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_30),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_69),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_62),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_135),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_63),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_1),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_28),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_53),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_151),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_25),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_143),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_17),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_24),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_5),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_157),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_159),
.B(n_0),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_158),
.B(n_0),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_186),
.B(n_1),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_2),
.Y(n_217)
);

BUFx8_ASAP7_75t_SL g218 ( 
.A(n_203),
.Y(n_218)
);

AND2x4_ASAP7_75t_L g219 ( 
.A(n_163),
.B(n_27),
.Y(n_219)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_160),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_3),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_4),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_154),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_4),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_174),
.B(n_32),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_182),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_175),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_182),
.Y(n_233)
);

AND2x6_ASAP7_75t_L g234 ( 
.A(n_184),
.B(n_153),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_161),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_188),
.B(n_6),
.Y(n_237)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_156),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_164),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_165),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_183),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_167),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_187),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_6),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_190),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_192),
.B(n_197),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g247 ( 
.A(n_191),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_194),
.B(n_7),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_204),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_8),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_209),
.B(n_210),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_169),
.B(n_9),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_170),
.B(n_9),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_171),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_155),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_222),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g259 ( 
.A1(n_215),
.A2(n_216),
.B1(n_254),
.B2(n_237),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_172),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_214),
.A2(n_203),
.B1(n_155),
.B2(n_185),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_217),
.A2(n_185),
.B1(n_177),
.B2(n_162),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_217),
.A2(n_177),
.B1(n_166),
.B2(n_202),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_221),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_224),
.A2(n_225),
.B1(n_244),
.B2(n_229),
.Y(n_265)
);

AO22x2_ASAP7_75t_L g266 ( 
.A1(n_224),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_225),
.A2(n_208),
.B1(n_206),
.B2(n_200),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_244),
.A2(n_181),
.B1(n_196),
.B2(n_195),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_221),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_223),
.B1(n_220),
.B2(n_232),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_232),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_173),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_220),
.A2(n_199),
.B1(n_193),
.B2(n_189),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_L g274 ( 
.A1(n_220),
.A2(n_180),
.B1(n_179),
.B2(n_178),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_176),
.Y(n_275)
);

AO22x2_ASAP7_75t_L g276 ( 
.A1(n_219),
.A2(n_230),
.B1(n_249),
.B2(n_251),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_256),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_33),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_221),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_221),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_235),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_249),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_220),
.B(n_13),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_251),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_L g285 ( 
.A1(n_220),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_220),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_219),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_287)
);

OA22x2_ASAP7_75t_L g288 ( 
.A1(n_241),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_235),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_235),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_L g291 ( 
.A1(n_223),
.A2(n_23),
.B1(n_25),
.B2(n_34),
.Y(n_291)
);

AND2x2_ASAP7_75t_SL g292 ( 
.A(n_219),
.B(n_230),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_256),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_235),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_230),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_243),
.Y(n_298)
);

OR2x6_ASAP7_75t_L g299 ( 
.A(n_247),
.B(n_43),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_223),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_223),
.B(n_49),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_243),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_236),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_243),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_243),
.Y(n_305)
);

OR2x6_ASAP7_75t_L g306 ( 
.A(n_247),
.B(n_56),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_223),
.B(n_227),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_259),
.B(n_255),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_262),
.B(n_255),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_298),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_246),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_258),
.B(n_223),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_271),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_271),
.B(n_227),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_305),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_255),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_276),
.A2(n_246),
.B(n_236),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_262),
.B(n_255),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_305),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_265),
.B(n_246),
.Y(n_321)
);

BUFx8_ASAP7_75t_L g322 ( 
.A(n_278),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_263),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_257),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_272),
.B(n_212),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_261),
.B(n_236),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_281),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_263),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_296),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_302),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_264),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_265),
.A2(n_234),
.B(n_245),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_276),
.B(n_242),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_269),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_279),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_268),
.B(n_242),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_288),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_275),
.A2(n_234),
.B(n_245),
.Y(n_339)
);

NAND2x1p5_ASAP7_75t_L g340 ( 
.A(n_297),
.B(n_213),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_268),
.B(n_212),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_267),
.B(n_213),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_280),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_289),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_294),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_260),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_295),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_304),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_266),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_304),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_270),
.B(n_238),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_283),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_301),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_297),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_306),
.B(n_233),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_303),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_303),
.Y(n_358)
);

XOR2x2_ASAP7_75t_L g359 ( 
.A(n_277),
.B(n_218),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_274),
.B(n_238),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_291),
.Y(n_361)
);

XOR2x2_ASAP7_75t_L g362 ( 
.A(n_282),
.B(n_226),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_273),
.B(n_238),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_287),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_287),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_293),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_285),
.B(n_238),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_286),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_266),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_300),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_299),
.B(n_233),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_282),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_299),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_315),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_311),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_321),
.B(n_226),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_326),
.B(n_306),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_335),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_325),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_334),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_335),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_346),
.B(n_238),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_284),
.Y(n_383)
);

AND2x2_ASAP7_75t_SL g384 ( 
.A(n_355),
.B(n_284),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_318),
.B(n_234),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_321),
.B(n_228),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_311),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_311),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_332),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_336),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_346),
.B(n_238),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_337),
.B(n_228),
.Y(n_392)
);

AND2x2_ASAP7_75t_SL g393 ( 
.A(n_355),
.B(n_231),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_354),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_343),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_344),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_313),
.B(n_231),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_345),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_342),
.B(n_239),
.Y(n_399)
);

NAND2x1p5_ASAP7_75t_L g400 ( 
.A(n_354),
.B(n_370),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_248),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_325),
.B(n_308),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_308),
.B(n_239),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_340),
.B(n_239),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_341),
.B(n_248),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_358),
.B(n_317),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_347),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_330),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_340),
.B(n_239),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_333),
.B(n_248),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_310),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_312),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_356),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_368),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_318),
.B(n_239),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_353),
.B(n_234),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_364),
.B(n_248),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_316),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_371),
.B(n_234),
.Y(n_420)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_371),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_320),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_365),
.B(n_248),
.Y(n_423)
);

AND2x6_ASAP7_75t_L g424 ( 
.A(n_369),
.B(n_250),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_361),
.B(n_250),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_314),
.B(n_239),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_372),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_324),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_363),
.B(n_234),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_372),
.B(n_250),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_339),
.B(n_240),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_309),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_360),
.A2(n_234),
.B(n_240),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_327),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_328),
.B(n_240),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_348),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_349),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_319),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_351),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_350),
.B(n_250),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_352),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_322),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_366),
.B(n_240),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_373),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_421),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_373),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_420),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_428),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_414),
.B(n_373),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_430),
.B(n_362),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_428),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_376),
.B(n_367),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_414),
.B(n_373),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_L g454 ( 
.A(n_379),
.B(n_363),
.Y(n_454)
);

NAND2x1p5_ASAP7_75t_L g455 ( 
.A(n_375),
.B(n_367),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_379),
.B(n_323),
.Y(n_456)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_388),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_384),
.B(n_323),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_375),
.B(n_329),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_427),
.Y(n_460)
);

OR2x6_ASAP7_75t_L g461 ( 
.A(n_442),
.B(n_350),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_434),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_378),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_376),
.B(n_362),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_384),
.B(n_329),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_434),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_430),
.B(n_359),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_392),
.B(n_359),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_381),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_406),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_381),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_378),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_389),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_402),
.B(n_322),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_389),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_432),
.B(n_250),
.Y(n_476)
);

NAND2x1_ASAP7_75t_SL g477 ( 
.A(n_374),
.B(n_57),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_375),
.B(n_58),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_420),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_386),
.B(n_240),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_402),
.Y(n_481)
);

AND2x2_ASAP7_75t_SL g482 ( 
.A(n_411),
.B(n_59),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_420),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_407),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_390),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_392),
.B(n_240),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_387),
.B(n_60),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_400),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_386),
.B(n_61),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_415),
.B(n_441),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_388),
.Y(n_493)
);

NOR2x1p5_ASAP7_75t_L g494 ( 
.A(n_442),
.B(n_65),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_411),
.B(n_66),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_395),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_407),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_395),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_441),
.B(n_67),
.Y(n_499)
);

INVx3_ASAP7_75t_SL g500 ( 
.A(n_461),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_463),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_447),
.Y(n_502)
);

BUFx12f_ASAP7_75t_L g503 ( 
.A(n_461),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_447),
.B(n_388),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_468),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_456),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_472),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_447),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_444),
.Y(n_509)
);

NOR2x1_ASAP7_75t_R g510 ( 
.A(n_456),
.B(n_383),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_470),
.B(n_418),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_476),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_452),
.B(n_418),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_444),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_469),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_445),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_445),
.Y(n_517)
);

BUFx10_ASAP7_75t_L g518 ( 
.A(n_474),
.Y(n_518)
);

OR2x6_ASAP7_75t_L g519 ( 
.A(n_445),
.B(n_400),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_452),
.A2(n_394),
.B1(n_405),
.B2(n_401),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_479),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_446),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_446),
.Y(n_523)
);

NAND2x1p5_ASAP7_75t_L g524 ( 
.A(n_489),
.B(n_387),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_474),
.Y(n_525)
);

NAND2x1p5_ASAP7_75t_L g526 ( 
.A(n_489),
.B(n_387),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_471),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_479),
.Y(n_528)
);

BUFx4f_ASAP7_75t_SL g529 ( 
.A(n_460),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_479),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_482),
.A2(n_481),
.B1(n_464),
.B2(n_458),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_484),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_484),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_470),
.B(n_491),
.Y(n_534)
);

BUFx6f_ASAP7_75t_SL g535 ( 
.A(n_459),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_484),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_449),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_454),
.B(n_423),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_461),
.Y(n_539)
);

BUFx6f_ASAP7_75t_SL g540 ( 
.A(n_459),
.Y(n_540)
);

CKINVDCx6p67_ASAP7_75t_R g541 ( 
.A(n_450),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_449),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_493),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_453),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_531),
.A2(n_465),
.B1(n_458),
.B2(n_464),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_515),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_515),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_534),
.A2(n_455),
.B1(n_491),
.B2(n_492),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_501),
.Y(n_549)
);

INVx6_ASAP7_75t_L g550 ( 
.A(n_521),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_501),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_527),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_527),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_506),
.A2(n_465),
.B1(n_482),
.B2(n_467),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_506),
.A2(n_438),
.B1(n_499),
.B2(n_380),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_513),
.A2(n_499),
.B1(n_377),
.B2(n_405),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_507),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_529),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_507),
.Y(n_559)
);

INVx1_ASAP7_75t_SL g560 ( 
.A(n_512),
.Y(n_560)
);

INVx6_ASAP7_75t_L g561 ( 
.A(n_521),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_511),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_513),
.A2(n_377),
.B1(n_453),
.B2(n_393),
.Y(n_563)
);

CKINVDCx11_ASAP7_75t_R g564 ( 
.A(n_500),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_519),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_519),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_505),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_528),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_538),
.A2(n_393),
.B1(n_423),
.B2(n_429),
.Y(n_569)
);

NAND2x1p5_ASAP7_75t_L g570 ( 
.A(n_516),
.B(n_517),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_SL g571 ( 
.A1(n_505),
.A2(n_488),
.B1(n_490),
.B2(n_492),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_539),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_538),
.A2(n_429),
.B1(n_383),
.B2(n_451),
.Y(n_573)
);

OAI22xp33_ASAP7_75t_L g574 ( 
.A1(n_525),
.A2(n_488),
.B1(n_466),
.B2(n_448),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_525),
.A2(n_462),
.B1(n_455),
.B2(n_399),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_541),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_500),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_519),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_519),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_538),
.B(n_440),
.Y(n_580)
);

INVx6_ASAP7_75t_L g581 ( 
.A(n_516),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_520),
.A2(n_490),
.B1(n_486),
.B2(n_496),
.Y(n_582)
);

INVx6_ASAP7_75t_L g583 ( 
.A(n_516),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_528),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_528),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_535),
.A2(n_494),
.B1(n_478),
.B2(n_425),
.Y(n_586)
);

CKINVDCx11_ASAP7_75t_R g587 ( 
.A(n_503),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_566),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_546),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_571),
.A2(n_541),
.B1(n_535),
.B2(n_540),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_545),
.A2(n_540),
.B1(n_535),
.B2(n_539),
.Y(n_591)
);

OAI222xp33_ASAP7_75t_L g592 ( 
.A1(n_554),
.A2(n_401),
.B1(n_483),
.B2(n_475),
.C1(n_498),
.C2(n_473),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_567),
.A2(n_503),
.B1(n_544),
.B2(n_542),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_574),
.A2(n_540),
.B1(n_518),
.B2(n_425),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_562),
.B(n_580),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_581),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_556),
.A2(n_518),
.B1(n_429),
.B2(n_443),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_555),
.A2(n_509),
.B1(n_514),
.B2(n_522),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_580),
.B(n_383),
.Y(n_599)
);

BUFx8_ASAP7_75t_SL g600 ( 
.A(n_567),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_575),
.A2(n_509),
.B1(n_514),
.B2(n_522),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_566),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_573),
.A2(n_518),
.B1(n_497),
.B2(n_485),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_566),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_552),
.Y(n_605)
);

NAND3xp33_ASAP7_75t_L g606 ( 
.A(n_586),
.B(n_382),
.C(n_391),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_552),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_563),
.A2(n_523),
.B1(n_544),
.B2(n_542),
.Y(n_608)
);

OAI22x1_ASAP7_75t_L g609 ( 
.A1(n_572),
.A2(n_524),
.B1(n_526),
.B2(n_543),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_547),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_587),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_581),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_549),
.B(n_440),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_548),
.A2(n_504),
.B1(n_537),
.B2(n_487),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_565),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_581),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_569),
.A2(n_504),
.B1(n_537),
.B2(n_397),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_560),
.A2(n_523),
.B1(n_495),
.B2(n_526),
.Y(n_618)
);

BUFx4f_ASAP7_75t_L g619 ( 
.A(n_581),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_564),
.A2(n_504),
.B1(n_397),
.B2(n_478),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_565),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_SL g622 ( 
.A1(n_577),
.A2(n_433),
.B(n_495),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_553),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_557),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_559),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_564),
.A2(n_493),
.B1(n_426),
.B2(n_419),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_568),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_549),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_551),
.B(n_530),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_582),
.A2(n_510),
.B(n_409),
.Y(n_630)
);

BUFx4f_ASAP7_75t_SL g631 ( 
.A(n_558),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_SL g632 ( 
.A1(n_576),
.A2(n_543),
.B1(n_536),
.B2(n_502),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_587),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_551),
.B(n_530),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_578),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_578),
.A2(n_493),
.B1(n_422),
.B2(n_419),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_583),
.Y(n_637)
);

OAI22xp33_ASAP7_75t_L g638 ( 
.A1(n_595),
.A2(n_576),
.B1(n_579),
.B2(n_558),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_SL g639 ( 
.A1(n_593),
.A2(n_579),
.B1(n_583),
.B2(n_524),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_591),
.A2(n_398),
.B1(n_410),
.B2(n_408),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_590),
.A2(n_398),
.B1(n_410),
.B2(n_408),
.Y(n_641)
);

AOI221xp5_ASAP7_75t_SL g642 ( 
.A1(n_626),
.A2(n_585),
.B1(n_584),
.B2(n_396),
.C(n_422),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_620),
.A2(n_583),
.B1(n_526),
.B2(n_524),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_599),
.B(n_477),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_597),
.A2(n_396),
.B1(n_403),
.B2(n_437),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_594),
.A2(n_617),
.B1(n_614),
.B2(n_619),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_606),
.A2(n_437),
.B1(n_439),
.B2(n_530),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_608),
.A2(n_439),
.B1(n_532),
.B2(n_583),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_605),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_SL g650 ( 
.A1(n_601),
.A2(n_561),
.B1(n_550),
.B2(n_517),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_598),
.A2(n_424),
.B1(n_480),
.B2(n_532),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_619),
.A2(n_457),
.B1(n_570),
.B2(n_532),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_618),
.A2(n_404),
.B1(n_521),
.B2(n_533),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_600),
.A2(n_521),
.B1(n_533),
.B2(n_424),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_600),
.A2(n_521),
.B1(n_533),
.B2(n_424),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_619),
.A2(n_457),
.B1(n_570),
.B2(n_508),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_603),
.A2(n_533),
.B1(n_424),
.B2(n_480),
.Y(n_657)
);

OAI221xp5_ASAP7_75t_SL g658 ( 
.A1(n_630),
.A2(n_508),
.B1(n_502),
.B2(n_436),
.C(n_416),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_636),
.A2(n_457),
.B1(n_517),
.B2(n_550),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_615),
.A2(n_533),
.B1(n_424),
.B2(n_536),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_615),
.A2(n_424),
.B1(n_536),
.B2(n_457),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_621),
.A2(n_561),
.B1(n_550),
.B2(n_412),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_613),
.B(n_561),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_621),
.A2(n_413),
.B1(n_412),
.B2(n_385),
.Y(n_664)
);

OAI222xp33_ASAP7_75t_L g665 ( 
.A1(n_635),
.A2(n_385),
.B1(n_417),
.B2(n_413),
.C1(n_412),
.C2(n_431),
.Y(n_665)
);

OAI211xp5_ASAP7_75t_L g666 ( 
.A1(n_622),
.A2(n_413),
.B(n_435),
.C(n_71),
.Y(n_666)
);

NAND4xp25_ASAP7_75t_L g667 ( 
.A(n_624),
.B(n_385),
.C(n_417),
.D(n_72),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_613),
.B(n_629),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_635),
.B(n_68),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_627),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_632),
.A2(n_417),
.B1(n_75),
.B2(n_76),
.Y(n_671)
);

OAI222xp33_ASAP7_75t_L g672 ( 
.A1(n_611),
.A2(n_70),
.B1(n_77),
.B2(n_78),
.C1(n_80),
.C2(n_81),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_602),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_673)
);

OAI22x1_ASAP7_75t_L g674 ( 
.A1(n_589),
.A2(n_610),
.B1(n_623),
.B2(n_625),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_SL g675 ( 
.A1(n_611),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_638),
.B(n_592),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_642),
.B(n_588),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_670),
.B(n_607),
.Y(n_678)
);

NAND4xp25_ASAP7_75t_L g679 ( 
.A(n_658),
.B(n_634),
.C(n_629),
.D(n_628),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_668),
.B(n_605),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_674),
.B(n_607),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_674),
.B(n_602),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g683 ( 
.A1(n_641),
.A2(n_633),
.B1(n_631),
.B2(n_637),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_663),
.B(n_602),
.Y(n_684)
);

NAND4xp25_ASAP7_75t_L g685 ( 
.A(n_667),
.B(n_634),
.C(n_637),
.D(n_616),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_649),
.B(n_588),
.Y(n_686)
);

OAI221xp5_ASAP7_75t_L g687 ( 
.A1(n_667),
.A2(n_633),
.B1(n_637),
.B2(n_616),
.C(n_612),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_649),
.B(n_604),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_644),
.B(n_639),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_669),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_669),
.B(n_604),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_646),
.B(n_604),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_651),
.Y(n_693)
);

NAND3xp33_ASAP7_75t_L g694 ( 
.A(n_666),
.B(n_604),
.C(n_588),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_651),
.B(n_604),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_640),
.B(n_588),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_653),
.B(n_588),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_643),
.B(n_616),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_648),
.B(n_609),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_650),
.B(n_609),
.Y(n_700)
);

OA21x2_ASAP7_75t_L g701 ( 
.A1(n_665),
.A2(n_612),
.B(n_596),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_647),
.B(n_596),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_662),
.B(n_88),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_645),
.B(n_657),
.Y(n_704)
);

NOR3xp33_ASAP7_75t_L g705 ( 
.A(n_687),
.B(n_672),
.C(n_675),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_681),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_684),
.B(n_654),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_682),
.Y(n_708)
);

NOR2x1_ASAP7_75t_L g709 ( 
.A(n_694),
.B(n_652),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_678),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_691),
.B(n_655),
.Y(n_711)
);

NAND3xp33_ASAP7_75t_L g712 ( 
.A(n_676),
.B(n_673),
.C(n_671),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_676),
.A2(n_656),
.B1(n_659),
.B2(n_664),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_700),
.B(n_660),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_690),
.B(n_661),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_680),
.B(n_90),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_706),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_708),
.B(n_693),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_709),
.B(n_689),
.Y(n_719)
);

OA22x2_ASAP7_75t_L g720 ( 
.A1(n_713),
.A2(n_689),
.B1(n_683),
.B2(n_692),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_710),
.B(n_688),
.Y(n_721)
);

AND2x4_ASAP7_75t_SL g722 ( 
.A(n_707),
.B(n_697),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_711),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_715),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_714),
.Y(n_725)
);

XNOR2xp5_ASAP7_75t_L g726 ( 
.A(n_720),
.B(n_712),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_717),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_724),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_722),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_724),
.B(n_698),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_721),
.Y(n_731)
);

OA22x2_ASAP7_75t_L g732 ( 
.A1(n_726),
.A2(n_722),
.B1(n_723),
.B2(n_725),
.Y(n_732)
);

OA22x2_ASAP7_75t_L g733 ( 
.A1(n_726),
.A2(n_723),
.B1(n_720),
.B2(n_719),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_729),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_727),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_728),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_735),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_735),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_734),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_736),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_739),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_737),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_741),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_742),
.Y(n_744)
);

NAND4xp25_ASAP7_75t_SL g745 ( 
.A(n_742),
.B(n_739),
.C(n_733),
.D(n_705),
.Y(n_745)
);

OAI221xp5_ASAP7_75t_L g746 ( 
.A1(n_743),
.A2(n_719),
.B1(n_744),
.B2(n_732),
.C(n_745),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_745),
.A2(n_732),
.B1(n_740),
.B2(n_738),
.Y(n_747)
);

NOR2x1_ASAP7_75t_L g748 ( 
.A(n_745),
.B(n_730),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_745),
.B(n_731),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_743),
.Y(n_750)
);

AO22x2_ASAP7_75t_L g751 ( 
.A1(n_744),
.A2(n_712),
.B1(n_705),
.B2(n_716),
.Y(n_751)
);

NOR3xp33_ASAP7_75t_L g752 ( 
.A(n_746),
.B(n_716),
.C(n_703),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_750),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_751),
.A2(n_685),
.B1(n_718),
.B2(n_679),
.Y(n_754)
);

AND3x4_ASAP7_75t_L g755 ( 
.A(n_748),
.B(n_698),
.C(n_677),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_747),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_749),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_750),
.Y(n_758)
);

AO22x2_ASAP7_75t_L g759 ( 
.A1(n_756),
.A2(n_677),
.B1(n_702),
.B2(n_699),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_753),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_758),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_L g762 ( 
.A(n_757),
.B(n_704),
.C(n_686),
.Y(n_762)
);

AND4x1_ASAP7_75t_L g763 ( 
.A(n_752),
.B(n_696),
.C(n_697),
.D(n_695),
.Y(n_763)
);

AO22x2_ASAP7_75t_L g764 ( 
.A1(n_755),
.A2(n_701),
.B1(n_93),
.B2(n_94),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_754),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_756),
.A2(n_701),
.B1(n_95),
.B2(n_99),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_760),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_761),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_765),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_762),
.Y(n_770)
);

NOR3xp33_ASAP7_75t_L g771 ( 
.A(n_766),
.B(n_91),
.C(n_100),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_764),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_763),
.Y(n_773)
);

NOR2x1_ASAP7_75t_L g774 ( 
.A(n_759),
.B(n_701),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_769),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_773),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_772),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_770),
.Y(n_778)
);

OAI22x1_ASAP7_75t_L g779 ( 
.A1(n_767),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_768),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_780)
);

OAI22x1_ASAP7_75t_L g781 ( 
.A1(n_774),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_781)
);

AOI31xp33_ASAP7_75t_L g782 ( 
.A1(n_771),
.A2(n_120),
.A3(n_122),
.B(n_124),
.Y(n_782)
);

OAI22xp33_ASAP7_75t_L g783 ( 
.A1(n_771),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_778),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_775),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_781),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_777),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_779),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_776),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_782),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_785),
.A2(n_783),
.B1(n_780),
.B2(n_140),
.Y(n_791)
);

AOI211xp5_ASAP7_75t_L g792 ( 
.A1(n_785),
.A2(n_134),
.B(n_137),
.C(n_141),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_784),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_791),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_794),
.A2(n_786),
.B1(n_790),
.B2(n_788),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_795),
.Y(n_796)
);

OA22x2_ASAP7_75t_L g797 ( 
.A1(n_796),
.A2(n_787),
.B1(n_789),
.B2(n_793),
.Y(n_797)
);

AOI211xp5_ASAP7_75t_L g798 ( 
.A1(n_797),
.A2(n_792),
.B(n_146),
.C(n_147),
.Y(n_798)
);


endmodule