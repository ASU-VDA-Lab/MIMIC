module fake_jpeg_24277_n_45 (n_3, n_2, n_1, n_0, n_4, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx5_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

INVx8_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx11_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_2),
.Y(n_13)
);

OAI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_14),
.A2(n_7),
.B1(n_9),
.B2(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_15),
.B(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_1),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_16),
.A2(n_18),
.B(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp67_ASAP7_75t_SL g24 ( 
.A(n_20),
.B(n_19),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_4),
.C(n_5),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_10),
.C(n_5),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_24),
.B(n_25),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_15),
.B1(n_7),
.B2(n_9),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_20),
.C(n_17),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_16),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_21),
.B1(n_8),
.B2(n_11),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_22),
.B1(n_19),
.B2(n_18),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_33),
.C(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_35),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_11),
.Y(n_40)
);

FAx1_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_11),
.CI(n_33),
.CON(n_37),
.SN(n_37)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_34),
.Y(n_39)
);

A2O1A1O1Ixp25_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_40),
.B(n_37),
.C(n_38),
.D(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_38),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_36),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_43),
.C(n_40),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_37),
.Y(n_45)
);


endmodule