module fake_netlist_1_10342_n_999 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_999);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_999;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_964;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_817;
wire n_985;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_769;
wire n_927;
wire n_596;
wire n_951;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_303;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_624;
wire n_426;
wire n_725;
wire n_818;
wire n_844;
wire n_738;
wire n_979;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_828;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_939;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_950;
wire n_910;
wire n_460;
wire n_478;
wire n_482;
wire n_415;
wire n_703;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_823;
wire n_970;
wire n_822;
wire n_984;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_539;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_947;
wire n_924;
wire n_912;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_992;
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_223), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_262), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_196), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_283), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_97), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_56), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_11), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_51), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_71), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_26), .Y(n_299) );
BUFx10_ASAP7_75t_L g300 ( .A(n_275), .Y(n_300) );
CKINVDCx16_ASAP7_75t_R g301 ( .A(n_171), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_156), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_189), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_247), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_139), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_87), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_17), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_27), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_148), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_9), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_0), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_177), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_268), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_137), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_228), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_122), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_270), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_49), .Y(n_318) );
INVx2_ASAP7_75t_SL g319 ( .A(n_260), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g320 ( .A(n_233), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_230), .Y(n_321) );
INVxp33_ASAP7_75t_SL g322 ( .A(n_37), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_253), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_257), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_53), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_215), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_98), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_20), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_73), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_278), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_207), .Y(n_332) );
INVxp33_ASAP7_75t_L g333 ( .A(n_136), .Y(n_333) );
INVx1_ASAP7_75t_SL g334 ( .A(n_169), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_109), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_265), .B(n_54), .Y(n_336) );
INVxp67_ASAP7_75t_SL g337 ( .A(n_244), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_194), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_83), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_20), .Y(n_340) );
CKINVDCx16_ASAP7_75t_R g341 ( .A(n_204), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_68), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_96), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_106), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_197), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_128), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_168), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_93), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_229), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_214), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_37), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_75), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_184), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_282), .B(n_249), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_70), .Y(n_355) );
BUFx5_ASAP7_75t_L g356 ( .A(n_126), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_143), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_46), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_208), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_11), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_125), .Y(n_361) );
BUFx10_ASAP7_75t_L g362 ( .A(n_48), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_172), .Y(n_363) );
CKINVDCx14_ASAP7_75t_R g364 ( .A(n_138), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_85), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_69), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_72), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_199), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_32), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_124), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_81), .B(n_7), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_67), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_203), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_287), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_242), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_112), .Y(n_376) );
INVxp67_ASAP7_75t_L g377 ( .A(n_35), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_258), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_10), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_183), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_224), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_141), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_239), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_30), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_86), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_267), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_180), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_158), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_167), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_105), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_181), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_251), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_121), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_110), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_248), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_185), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_132), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_220), .Y(n_398) );
BUFx2_ASAP7_75t_L g399 ( .A(n_63), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_159), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_47), .Y(n_401) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_157), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_94), .Y(n_403) );
CKINVDCx16_ASAP7_75t_R g404 ( .A(n_111), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_95), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_213), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_161), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_192), .Y(n_408) );
BUFx10_ASAP7_75t_L g409 ( .A(n_288), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_142), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_225), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_274), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_32), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_108), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_107), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_123), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_279), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_52), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_62), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_113), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_209), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_218), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_285), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_178), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_256), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_43), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_59), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_166), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_236), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_211), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_263), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_116), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_77), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_165), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_264), .Y(n_435) );
BUFx2_ASAP7_75t_L g436 ( .A(n_328), .Y(n_436) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_361), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_328), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_333), .B(n_0), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_333), .B(n_1), .Y(n_440) );
OAI21x1_ASAP7_75t_L g441 ( .A1(n_297), .A2(n_55), .B(n_50), .Y(n_441) );
BUFx2_ASAP7_75t_L g442 ( .A(n_399), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_432), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_364), .B(n_1), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_319), .B(n_2), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_384), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_298), .B(n_2), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_356), .Y(n_448) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_361), .Y(n_449) );
OAI21x1_ASAP7_75t_L g450 ( .A1(n_324), .A2(n_58), .B(n_57), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_377), .A2(n_341), .B1(n_404), .B2(n_301), .Y(n_451) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_361), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_356), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_347), .B(n_3), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_364), .B(n_3), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_377), .B(n_4), .Y(n_456) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_361), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_322), .A2(n_6), .B1(n_4), .B2(n_5), .Y(n_458) );
AOI22xp5_ASAP7_75t_SL g459 ( .A1(n_426), .A2(n_8), .B1(n_5), .B2(n_6), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_370), .B(n_8), .Y(n_460) );
INVx4_ASAP7_75t_L g461 ( .A(n_290), .Y(n_461) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_385), .Y(n_462) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_385), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_307), .B(n_10), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_308), .B(n_12), .Y(n_465) );
BUFx8_ASAP7_75t_SL g466 ( .A(n_316), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_448), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_448), .B(n_356), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_453), .Y(n_469) );
BUFx4f_ASAP7_75t_L g470 ( .A(n_444), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_464), .Y(n_471) );
AND2x2_ASAP7_75t_SL g472 ( .A(n_444), .B(n_371), .Y(n_472) );
OAI22xp33_ASAP7_75t_SL g473 ( .A1(n_458), .A2(n_299), .B1(n_311), .B2(n_296), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_453), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_437), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_437), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_464), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_446), .Y(n_478) );
INVx5_ASAP7_75t_L g479 ( .A(n_437), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_439), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_437), .Y(n_481) );
OAI22xp33_ASAP7_75t_SL g482 ( .A1(n_451), .A2(n_329), .B1(n_379), .B2(n_340), .Y(n_482) );
OAI22xp33_ASAP7_75t_L g483 ( .A1(n_436), .A2(n_351), .B1(n_369), .B2(n_360), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_439), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_445), .B(n_356), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_440), .Y(n_486) );
INVx2_ASAP7_75t_SL g487 ( .A(n_436), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_449), .Y(n_488) );
INVx4_ASAP7_75t_L g489 ( .A(n_455), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_438), .B(n_356), .Y(n_490) );
NAND2xp33_ASAP7_75t_SL g491 ( .A(n_455), .B(n_320), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_478), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_489), .B(n_440), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_480), .B(n_441), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_478), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_487), .B(n_442), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_484), .B(n_441), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_467), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_467), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_489), .B(n_461), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_489), .B(n_461), .Y(n_501) );
NAND3xp33_ASAP7_75t_L g502 ( .A(n_486), .B(n_443), .C(n_456), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_471), .B(n_461), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_477), .B(n_447), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_472), .B(n_454), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_472), .B(n_460), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_470), .B(n_401), .Y(n_507) );
INVxp67_ASAP7_75t_L g508 ( .A(n_491), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_470), .B(n_450), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_490), .Y(n_510) );
NOR2xp67_ASAP7_75t_L g511 ( .A(n_490), .B(n_465), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_485), .B(n_300), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_485), .B(n_291), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_469), .B(n_450), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_483), .A2(n_346), .B1(n_357), .B2(n_348), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_474), .B(n_293), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_474), .B(n_294), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_468), .Y(n_518) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_468), .Y(n_519) );
BUFx3_ASAP7_75t_L g520 ( .A(n_479), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_482), .B(n_302), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_473), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_479), .B(n_305), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_479), .B(n_300), .Y(n_524) );
INVxp67_ASAP7_75t_L g525 ( .A(n_475), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_475), .B(n_362), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_476), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_505), .A2(n_310), .B(n_337), .C(n_292), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_506), .B(n_466), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_509), .A2(n_337), .B(n_295), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_508), .B(n_459), .Y(n_531) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_493), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_494), .A2(n_304), .B(n_303), .Y(n_533) );
O2A1O1Ixp33_ASAP7_75t_SL g534 ( .A1(n_494), .A2(n_354), .B(n_336), .C(n_309), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_522), .A2(n_387), .B1(n_388), .B2(n_378), .Y(n_535) );
NOR2x1p5_ASAP7_75t_SL g536 ( .A(n_518), .B(n_356), .Y(n_536) );
BUFx3_ASAP7_75t_L g537 ( .A(n_520), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_496), .B(n_413), .Y(n_538) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_497), .A2(n_317), .B(n_314), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_514), .A2(n_323), .B(n_321), .Y(n_540) );
INVx3_ASAP7_75t_L g541 ( .A(n_520), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_514), .A2(n_335), .B(n_326), .Y(n_542) );
BUFx2_ASAP7_75t_L g543 ( .A(n_515), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_526), .B(n_397), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_500), .B(n_306), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_502), .A2(n_339), .B(n_342), .C(n_338), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_507), .B(n_407), .Y(n_547) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_498), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_501), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_503), .A2(n_504), .B(n_510), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_511), .A2(n_349), .B(n_350), .C(n_343), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_526), .B(n_313), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_492), .B(n_315), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_495), .B(n_318), .Y(n_554) );
AOI21xp33_ASAP7_75t_L g555 ( .A1(n_512), .A2(n_521), .B(n_513), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_512), .B(n_325), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_516), .A2(n_368), .B(n_352), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_499), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_499), .A2(n_375), .B(n_380), .C(n_373), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_517), .A2(n_382), .B(n_381), .Y(n_560) );
OAI21x1_ASAP7_75t_L g561 ( .A1(n_523), .A2(n_390), .B(n_383), .Y(n_561) );
INVx2_ASAP7_75t_SL g562 ( .A(n_524), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_519), .B(n_409), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_519), .B(n_327), .Y(n_564) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_519), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_527), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_525), .B(n_391), .Y(n_567) );
O2A1O1Ixp5_ASAP7_75t_L g568 ( .A1(n_555), .A2(n_392), .B(n_400), .C(n_395), .Y(n_568) );
OAI21x1_ASAP7_75t_L g569 ( .A1(n_561), .A2(n_406), .B(n_403), .Y(n_569) );
NAND2x1p5_ASAP7_75t_L g570 ( .A(n_537), .B(n_358), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_550), .A2(n_412), .B(n_408), .Y(n_571) );
AND2x6_ASAP7_75t_L g572 ( .A(n_541), .B(n_416), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_558), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_535), .Y(n_574) );
OAI21x1_ASAP7_75t_L g575 ( .A1(n_540), .A2(n_420), .B(n_417), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_535), .B(n_13), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_532), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g578 ( .A1(n_555), .A2(n_423), .B(n_427), .C(n_421), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_531), .B(n_358), .Y(n_579) );
OAI21x1_ASAP7_75t_L g580 ( .A1(n_542), .A2(n_431), .B(n_429), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_533), .A2(n_435), .B(n_434), .Y(n_581) );
NAND2x1_ASAP7_75t_L g582 ( .A(n_548), .B(n_385), .Y(n_582) );
OAI21x1_ASAP7_75t_L g583 ( .A1(n_539), .A2(n_488), .B(n_481), .Y(n_583) );
AO31x2_ASAP7_75t_L g584 ( .A1(n_530), .A2(n_452), .A3(n_463), .B(n_457), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_539), .A2(n_334), .B(n_312), .Y(n_585) );
AO21x2_ASAP7_75t_L g586 ( .A1(n_534), .A2(n_402), .B(n_452), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_549), .B(n_358), .Y(n_587) );
NAND2x1_ASAP7_75t_L g588 ( .A(n_548), .B(n_402), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_544), .B(n_330), .Y(n_589) );
OAI22x1_ASAP7_75t_L g590 ( .A1(n_547), .A2(n_418), .B1(n_331), .B2(n_332), .Y(n_590) );
BUFx3_ASAP7_75t_L g591 ( .A(n_541), .Y(n_591) );
OAI21x1_ASAP7_75t_L g592 ( .A1(n_566), .A2(n_402), .B(n_61), .Y(n_592) );
AO31x2_ASAP7_75t_L g593 ( .A1(n_559), .A2(n_452), .A3(n_463), .B(n_457), .Y(n_593) );
AOI21xp33_ASAP7_75t_L g594 ( .A1(n_529), .A2(n_538), .B(n_528), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_548), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_553), .A2(n_345), .B(n_344), .Y(n_596) );
NOR2x1_ASAP7_75t_SL g597 ( .A(n_565), .B(n_365), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_554), .A2(n_355), .B(n_353), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_557), .A2(n_363), .B(n_359), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_552), .B(n_366), .Y(n_600) );
OAI21x1_ASAP7_75t_L g601 ( .A1(n_560), .A2(n_64), .B(n_60), .Y(n_601) );
AOI21xp33_ASAP7_75t_L g602 ( .A1(n_562), .A2(n_372), .B(n_367), .Y(n_602) );
INVx3_ASAP7_75t_SL g603 ( .A(n_564), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_545), .A2(n_376), .B(n_374), .Y(n_604) );
AO31x2_ASAP7_75t_L g605 ( .A1(n_551), .A2(n_546), .A3(n_567), .B(n_563), .Y(n_605) );
OAI21x1_ASAP7_75t_L g606 ( .A1(n_567), .A2(n_66), .B(n_65), .Y(n_606) );
AO31x2_ASAP7_75t_L g607 ( .A1(n_536), .A2(n_463), .A3(n_452), .B(n_457), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_565), .B(n_386), .Y(n_608) );
AOI21x1_ASAP7_75t_L g609 ( .A1(n_556), .A2(n_565), .B(n_463), .Y(n_609) );
A2O1A1Ixp33_ASAP7_75t_L g610 ( .A1(n_550), .A2(n_411), .B(n_463), .C(n_452), .Y(n_610) );
BUFx12f_ASAP7_75t_L g611 ( .A(n_543), .Y(n_611) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_573), .Y(n_612) );
NAND3xp33_ASAP7_75t_L g613 ( .A(n_610), .B(n_457), .C(n_449), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_574), .A2(n_393), .B1(n_394), .B2(n_389), .Y(n_614) );
AO21x2_ASAP7_75t_L g615 ( .A1(n_609), .A2(n_462), .B(n_449), .Y(n_615) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_594), .A2(n_424), .B1(n_398), .B2(n_433), .C(n_430), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_572), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_593), .Y(n_618) );
NOR2x1_ASAP7_75t_R g619 ( .A(n_611), .B(n_396), .Y(n_619) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_577), .Y(n_620) );
OAI21x1_ASAP7_75t_SL g621 ( .A1(n_597), .A2(n_14), .B(n_15), .Y(n_621) );
OA21x2_ASAP7_75t_L g622 ( .A1(n_592), .A2(n_410), .B(n_405), .Y(n_622) );
INVx3_ASAP7_75t_L g623 ( .A(n_591), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_578), .B(n_14), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g625 ( .A1(n_568), .A2(n_415), .B(n_414), .Y(n_625) );
OA21x2_ASAP7_75t_L g626 ( .A1(n_606), .A2(n_422), .B(n_419), .Y(n_626) );
BUFx2_ASAP7_75t_L g627 ( .A(n_572), .Y(n_627) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_570), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_576), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_571), .A2(n_462), .B(n_425), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_572), .Y(n_631) );
OAI21x1_ASAP7_75t_L g632 ( .A1(n_583), .A2(n_462), .B(n_76), .Y(n_632) );
OAI21x1_ASAP7_75t_L g633 ( .A1(n_569), .A2(n_78), .B(n_74), .Y(n_633) );
OAI21x1_ASAP7_75t_L g634 ( .A1(n_582), .A2(n_80), .B(n_79), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_587), .Y(n_635) );
OAI21x1_ASAP7_75t_L g636 ( .A1(n_588), .A2(n_84), .B(n_82), .Y(n_636) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_595), .Y(n_637) );
BUFx2_ASAP7_75t_R g638 ( .A(n_603), .Y(n_638) );
OAI21x1_ASAP7_75t_SL g639 ( .A1(n_597), .A2(n_16), .B(n_17), .Y(n_639) );
AO21x1_ASAP7_75t_L g640 ( .A1(n_579), .A2(n_18), .B(n_19), .Y(n_640) );
INVx8_ASAP7_75t_L g641 ( .A(n_590), .Y(n_641) );
OAI21x1_ASAP7_75t_L g642 ( .A1(n_601), .A2(n_89), .B(n_88), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_593), .Y(n_643) );
OA21x2_ASAP7_75t_L g644 ( .A1(n_575), .A2(n_428), .B(n_91), .Y(n_644) );
BUFx2_ASAP7_75t_SL g645 ( .A(n_595), .Y(n_645) );
OAI21x1_ASAP7_75t_L g646 ( .A1(n_580), .A2(n_92), .B(n_90), .Y(n_646) );
NAND2x1p5_ASAP7_75t_L g647 ( .A(n_608), .B(n_19), .Y(n_647) );
OAI21xp5_ASAP7_75t_L g648 ( .A1(n_581), .A2(n_21), .B(n_22), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_593), .Y(n_649) );
BUFx3_ASAP7_75t_L g650 ( .A(n_607), .Y(n_650) );
BUFx4f_ASAP7_75t_L g651 ( .A(n_602), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_589), .A2(n_23), .B1(n_24), .B2(n_25), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_584), .Y(n_653) );
INVx4_ASAP7_75t_L g654 ( .A(n_586), .Y(n_654) );
OAI21x1_ASAP7_75t_L g655 ( .A1(n_585), .A2(n_100), .B(n_99), .Y(n_655) );
OAI21x1_ASAP7_75t_L g656 ( .A1(n_596), .A2(n_102), .B(n_101), .Y(n_656) );
OAI21x1_ASAP7_75t_L g657 ( .A1(n_598), .A2(n_104), .B(n_103), .Y(n_657) );
OAI21x1_ASAP7_75t_L g658 ( .A1(n_607), .A2(n_115), .B(n_114), .Y(n_658) );
OAI21x1_ASAP7_75t_L g659 ( .A1(n_607), .A2(n_118), .B(n_117), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_600), .A2(n_23), .B1(n_24), .B2(n_25), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_599), .B(n_26), .Y(n_661) );
OAI21x1_ASAP7_75t_SL g662 ( .A1(n_604), .A2(n_27), .B(n_28), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_605), .Y(n_663) );
OAI21x1_ASAP7_75t_L g664 ( .A1(n_584), .A2(n_120), .B(n_119), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_605), .Y(n_665) );
OAI21x1_ASAP7_75t_SL g666 ( .A1(n_605), .A2(n_29), .B(n_30), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_574), .B(n_31), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_577), .Y(n_668) );
AO21x2_ASAP7_75t_L g669 ( .A1(n_653), .A2(n_31), .B(n_33), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_620), .Y(n_670) );
OAI21xp5_ASAP7_75t_L g671 ( .A1(n_624), .A2(n_33), .B(n_34), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_612), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_620), .Y(n_673) );
BUFx3_ASAP7_75t_L g674 ( .A(n_623), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_668), .Y(n_675) );
BUFx3_ASAP7_75t_L g676 ( .A(n_641), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_629), .Y(n_677) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_637), .Y(n_678) );
INVxp67_ASAP7_75t_SL g679 ( .A(n_650), .Y(n_679) );
OR2x6_ASAP7_75t_L g680 ( .A(n_645), .B(n_35), .Y(n_680) );
BUFx4f_ASAP7_75t_L g681 ( .A(n_641), .Y(n_681) );
OAI222xp33_ASAP7_75t_L g682 ( .A1(n_660), .A2(n_36), .B1(n_38), .B2(n_39), .C1(n_40), .C2(n_41), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_660), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_652), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_663), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_665), .Y(n_686) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_618), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_635), .B(n_38), .Y(n_688) );
OAI21x1_ASAP7_75t_L g689 ( .A1(n_632), .A2(n_649), .B(n_643), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_652), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_647), .Y(n_691) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_624), .A2(n_39), .B(n_40), .Y(n_692) );
INVx3_ASAP7_75t_L g693 ( .A(n_628), .Y(n_693) );
INVxp67_ASAP7_75t_L g694 ( .A(n_617), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_647), .Y(n_695) );
INVx1_ASAP7_75t_SL g696 ( .A(n_617), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_666), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_631), .A2(n_41), .B1(n_42), .B2(n_43), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_648), .Y(n_699) );
INVxp67_ASAP7_75t_R g700 ( .A(n_638), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_615), .A2(n_289), .B(n_212), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_648), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_640), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_662), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_661), .Y(n_705) );
INVx1_ASAP7_75t_SL g706 ( .A(n_631), .Y(n_706) );
AOI21x1_ASAP7_75t_L g707 ( .A1(n_644), .A2(n_44), .B(n_45), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_621), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_626), .B(n_44), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_639), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_633), .Y(n_711) );
BUFx2_ASAP7_75t_L g712 ( .A(n_619), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_651), .A2(n_46), .B1(n_47), .B2(n_127), .Y(n_713) );
AND2x4_ASAP7_75t_L g714 ( .A(n_646), .B(n_129), .Y(n_714) );
OA21x2_ASAP7_75t_L g715 ( .A1(n_613), .A2(n_130), .B(n_131), .Y(n_715) );
INVx8_ASAP7_75t_L g716 ( .A(n_638), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_622), .Y(n_717) );
OR2x2_ASAP7_75t_L g718 ( .A(n_614), .B(n_286), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_664), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_622), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_656), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_657), .Y(n_722) );
INVx3_ASAP7_75t_L g723 ( .A(n_644), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_658), .Y(n_724) );
INVx2_ASAP7_75t_SL g725 ( .A(n_619), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_614), .Y(n_726) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_654), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_626), .B(n_625), .Y(n_728) );
NAND2x1_ASAP7_75t_L g729 ( .A(n_654), .B(n_133), .Y(n_729) );
AO21x1_ASAP7_75t_SL g730 ( .A1(n_625), .A2(n_134), .B(n_135), .Y(n_730) );
OA21x2_ASAP7_75t_L g731 ( .A1(n_613), .A2(n_140), .B(n_144), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_630), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_634), .Y(n_733) );
AOI22xp33_ASAP7_75t_SL g734 ( .A1(n_659), .A2(n_145), .B1(n_146), .B2(n_147), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_636), .Y(n_735) );
OAI21x1_ASAP7_75t_L g736 ( .A1(n_642), .A2(n_149), .B(n_150), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_655), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_616), .B(n_151), .Y(n_738) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_615), .Y(n_739) );
OR2x2_ASAP7_75t_L g740 ( .A(n_630), .B(n_284), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_616), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_667), .B(n_152), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_629), .B(n_153), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_629), .B(n_154), .Y(n_744) );
OR2x6_ASAP7_75t_L g745 ( .A(n_627), .B(n_155), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_685), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_686), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_687), .Y(n_748) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_678), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_672), .B(n_160), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_675), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_677), .Y(n_752) );
INVxp67_ASAP7_75t_SL g753 ( .A(n_678), .Y(n_753) );
INVx2_ASAP7_75t_SL g754 ( .A(n_674), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_670), .Y(n_755) );
BUFx2_ASAP7_75t_L g756 ( .A(n_680), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_705), .A2(n_162), .B1(n_163), .B2(n_164), .Y(n_757) );
CKINVDCx6p67_ASAP7_75t_R g758 ( .A(n_716), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_687), .Y(n_759) );
INVx3_ASAP7_75t_L g760 ( .A(n_745), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_689), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_723), .Y(n_762) );
OR2x2_ASAP7_75t_L g763 ( .A(n_673), .B(n_280), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_683), .A2(n_170), .B1(n_173), .B2(n_174), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_684), .A2(n_175), .B1(n_176), .B2(n_179), .Y(n_765) );
AOI22xp33_ASAP7_75t_SL g766 ( .A1(n_726), .A2(n_182), .B1(n_186), .B2(n_187), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_723), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_688), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_690), .B(n_188), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_745), .A2(n_190), .B1(n_191), .B2(n_193), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_699), .B(n_195), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_702), .B(n_198), .Y(n_772) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_727), .Y(n_773) );
INVx2_ASAP7_75t_L g774 ( .A(n_669), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_703), .B(n_200), .Y(n_775) );
AND2x4_ASAP7_75t_L g776 ( .A(n_745), .B(n_201), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_743), .Y(n_777) );
OAI21xp5_ASAP7_75t_SL g778 ( .A1(n_712), .A2(n_202), .B(n_205), .Y(n_778) );
INVx2_ASAP7_75t_SL g779 ( .A(n_681), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_742), .B(n_206), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_743), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_744), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_708), .B(n_210), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_716), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_719), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_744), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_691), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_695), .Y(n_788) );
BUFx6f_ASAP7_75t_L g789 ( .A(n_693), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_724), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_739), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_725), .B(n_216), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_711), .Y(n_793) );
INVxp67_ASAP7_75t_L g794 ( .A(n_727), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_741), .A2(n_217), .B1(n_219), .B2(n_221), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_709), .Y(n_796) );
INVx3_ASAP7_75t_L g797 ( .A(n_696), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_671), .Y(n_798) );
AND2x4_ASAP7_75t_L g799 ( .A(n_679), .B(n_222), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_671), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_692), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_692), .Y(n_802) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_696), .Y(n_803) );
AND2x2_ASAP7_75t_L g804 ( .A(n_700), .B(n_226), .Y(n_804) );
INVx3_ASAP7_75t_L g805 ( .A(n_706), .Y(n_805) );
AND2x4_ASAP7_75t_L g806 ( .A(n_694), .B(n_227), .Y(n_806) );
BUFx4f_ASAP7_75t_SL g807 ( .A(n_676), .Y(n_807) );
INVx2_ASAP7_75t_L g808 ( .A(n_717), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_698), .B(n_231), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_720), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_738), .A2(n_232), .B1(n_234), .B2(n_235), .Y(n_811) );
AND2x4_ASAP7_75t_L g812 ( .A(n_694), .B(n_237), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_710), .Y(n_813) );
BUFx2_ASAP7_75t_L g814 ( .A(n_732), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_704), .Y(n_815) );
OR2x2_ASAP7_75t_L g816 ( .A(n_716), .B(n_277), .Y(n_816) );
AND2x2_ASAP7_75t_L g817 ( .A(n_698), .B(n_238), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_707), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_718), .A2(n_240), .B1(n_241), .B2(n_243), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_697), .Y(n_820) );
INVx2_ASAP7_75t_SL g821 ( .A(n_729), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_713), .B(n_245), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_730), .B(n_246), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_728), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_733), .Y(n_825) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_737), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_735), .Y(n_827) );
INVx4_ASAP7_75t_L g828 ( .A(n_714), .Y(n_828) );
INVxp67_ASAP7_75t_L g829 ( .A(n_740), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_721), .Y(n_830) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_773), .Y(n_831) );
OR2x2_ASAP7_75t_L g832 ( .A(n_814), .B(n_722), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_752), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_794), .B(n_734), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_794), .B(n_734), .Y(n_835) );
AND2x2_ASAP7_75t_L g836 ( .A(n_751), .B(n_731), .Y(n_836) );
AND2x4_ASAP7_75t_L g837 ( .A(n_828), .B(n_701), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_755), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_746), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_749), .B(n_701), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_756), .A2(n_715), .B1(n_682), .B2(n_736), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_749), .B(n_715), .Y(n_842) );
INVx2_ASAP7_75t_L g843 ( .A(n_746), .Y(n_843) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_748), .Y(n_844) );
AND2x4_ASAP7_75t_L g845 ( .A(n_828), .B(n_753), .Y(n_845) );
INVx2_ASAP7_75t_L g846 ( .A(n_747), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_787), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_788), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_796), .B(n_250), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_754), .B(n_252), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_798), .B(n_254), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_808), .Y(n_852) );
BUFx3_ASAP7_75t_L g853 ( .A(n_807), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_800), .B(n_255), .Y(n_854) );
AND2x4_ASAP7_75t_L g855 ( .A(n_760), .B(n_259), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_813), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_785), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_790), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_768), .B(n_261), .Y(n_859) );
AND2x4_ASAP7_75t_L g860 ( .A(n_760), .B(n_266), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_815), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_759), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_803), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_803), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_801), .B(n_269), .Y(n_865) );
AOI22xp33_ASAP7_75t_SL g866 ( .A1(n_776), .A2(n_271), .B1(n_272), .B2(n_273), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_820), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_802), .B(n_276), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_797), .B(n_805), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_797), .B(n_805), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_826), .Y(n_871) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_829), .A2(n_776), .B1(n_770), .B2(n_766), .Y(n_872) );
HB1xp67_ASAP7_75t_L g873 ( .A(n_791), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_830), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_777), .B(n_781), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_824), .B(n_782), .Y(n_876) );
NOR2x1p5_ASAP7_75t_L g877 ( .A(n_758), .B(n_816), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_786), .B(n_750), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_810), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_775), .B(n_774), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_775), .Y(n_881) );
AOI22xp33_ASAP7_75t_SL g882 ( .A1(n_799), .A2(n_770), .B1(n_817), .B2(n_809), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_766), .A2(n_778), .B1(n_819), .B2(n_763), .Y(n_883) );
AOI22xp33_ASAP7_75t_SL g884 ( .A1(n_784), .A2(n_780), .B1(n_812), .B2(n_806), .Y(n_884) );
INVx4_ASAP7_75t_L g885 ( .A(n_789), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_783), .Y(n_886) );
AND2x4_ASAP7_75t_L g887 ( .A(n_762), .B(n_767), .Y(n_887) );
CKINVDCx10_ASAP7_75t_R g888 ( .A(n_779), .Y(n_888) );
NOR2xp67_ASAP7_75t_L g889 ( .A(n_872), .B(n_804), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_833), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_875), .B(n_818), .Y(n_891) );
INVx4_ASAP7_75t_L g892 ( .A(n_853), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_869), .B(n_812), .Y(n_893) );
AND2x4_ASAP7_75t_L g894 ( .A(n_845), .B(n_821), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_870), .B(n_806), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_844), .Y(n_896) );
OR2x2_ASAP7_75t_L g897 ( .A(n_831), .B(n_827), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_838), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_847), .Y(n_899) );
OR2x2_ASAP7_75t_L g900 ( .A(n_844), .B(n_827), .Y(n_900) );
OR2x2_ASAP7_75t_L g901 ( .A(n_863), .B(n_825), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_848), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_856), .Y(n_903) );
OR2x2_ASAP7_75t_L g904 ( .A(n_864), .B(n_825), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_861), .Y(n_905) );
AND2x4_ASAP7_75t_L g906 ( .A(n_832), .B(n_793), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_876), .B(n_793), .Y(n_907) );
INVx2_ASAP7_75t_L g908 ( .A(n_873), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_876), .B(n_769), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_871), .B(n_761), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_873), .Y(n_911) );
INVx2_ASAP7_75t_L g912 ( .A(n_839), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_878), .B(n_823), .Y(n_913) );
BUFx2_ASAP7_75t_SL g914 ( .A(n_853), .Y(n_914) );
INVxp67_ASAP7_75t_SL g915 ( .A(n_842), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_867), .Y(n_916) );
OR2x2_ASAP7_75t_L g917 ( .A(n_862), .B(n_772), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_881), .B(n_772), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_843), .B(n_771), .Y(n_919) );
INVx2_ASAP7_75t_SL g920 ( .A(n_888), .Y(n_920) );
OR2x2_ASAP7_75t_L g921 ( .A(n_846), .B(n_792), .Y(n_921) );
OR2x2_ASAP7_75t_L g922 ( .A(n_846), .B(n_757), .Y(n_922) );
BUFx2_ASAP7_75t_L g923 ( .A(n_885), .Y(n_923) );
HB1xp67_ASAP7_75t_L g924 ( .A(n_852), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_890), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_898), .Y(n_926) );
AND2x4_ASAP7_75t_SL g927 ( .A(n_892), .B(n_850), .Y(n_927) );
OR2x6_ASAP7_75t_L g928 ( .A(n_914), .B(n_837), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_893), .B(n_887), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_899), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_895), .B(n_887), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_891), .B(n_835), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_891), .B(n_834), .Y(n_933) );
AOI21xp33_ASAP7_75t_SL g934 ( .A1(n_920), .A2(n_883), .B(n_884), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_902), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_903), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_905), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_889), .B(n_886), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_916), .B(n_882), .Y(n_939) );
OR2x6_ASAP7_75t_L g940 ( .A(n_894), .B(n_877), .Y(n_940) );
OR2x2_ASAP7_75t_L g941 ( .A(n_896), .B(n_879), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_915), .B(n_874), .Y(n_942) );
OR2x2_ASAP7_75t_L g943 ( .A(n_908), .B(n_879), .Y(n_943) );
NOR2x1_ASAP7_75t_L g944 ( .A(n_923), .B(n_885), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_915), .B(n_840), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_907), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_907), .Y(n_947) );
OR2x2_ASAP7_75t_L g948 ( .A(n_911), .B(n_880), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_942), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_946), .B(n_913), .Y(n_950) );
NAND3xp33_ASAP7_75t_L g951 ( .A(n_934), .B(n_866), .C(n_841), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_942), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_947), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_925), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_926), .Y(n_955) );
AOI22xp5_ASAP7_75t_L g956 ( .A1(n_939), .A2(n_940), .B1(n_932), .B2(n_933), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g957 ( .A1(n_940), .A2(n_841), .B1(n_909), .B2(n_921), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_930), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_945), .B(n_906), .Y(n_959) );
INVx3_ASAP7_75t_L g960 ( .A(n_940), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_935), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_938), .B(n_906), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_936), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_937), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_960), .A2(n_944), .B1(n_928), .B2(n_927), .Y(n_965) );
AO22x1_ASAP7_75t_L g966 ( .A1(n_957), .A2(n_855), .B1(n_860), .B2(n_931), .Y(n_966) );
OA22x2_ASAP7_75t_L g967 ( .A1(n_956), .A2(n_929), .B1(n_860), .B2(n_855), .Y(n_967) );
OA21x2_ASAP7_75t_L g968 ( .A1(n_951), .A2(n_949), .B(n_952), .Y(n_968) );
INVx1_ASAP7_75t_SL g969 ( .A(n_950), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_953), .Y(n_970) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_951), .A2(n_943), .B1(n_941), .B2(n_948), .Y(n_971) );
INVx2_ASAP7_75t_SL g972 ( .A(n_959), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_954), .Y(n_973) );
AOI211xp5_ASAP7_75t_L g974 ( .A1(n_965), .A2(n_964), .B(n_963), .C(n_961), .Y(n_974) );
AOI221x1_ASAP7_75t_L g975 ( .A1(n_971), .A2(n_958), .B1(n_955), .B2(n_962), .C(n_849), .Y(n_975) );
OAI222xp33_ASAP7_75t_L g976 ( .A1(n_967), .A2(n_918), .B1(n_922), .B2(n_917), .C1(n_904), .C2(n_901), .Y(n_976) );
NAND3xp33_ASAP7_75t_L g977 ( .A(n_968), .B(n_757), .C(n_764), .Y(n_977) );
AOI21xp5_ASAP7_75t_L g978 ( .A1(n_966), .A2(n_924), .B(n_910), .Y(n_978) );
NOR2xp33_ASAP7_75t_L g979 ( .A(n_969), .B(n_897), .Y(n_979) );
NAND3xp33_ASAP7_75t_SL g980 ( .A(n_974), .B(n_970), .C(n_973), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_979), .Y(n_981) );
NOR2xp33_ASAP7_75t_SL g982 ( .A(n_976), .B(n_972), .Y(n_982) );
NAND4xp25_ASAP7_75t_L g983 ( .A(n_977), .B(n_811), .C(n_765), .D(n_764), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_981), .Y(n_984) );
NOR2x1_ASAP7_75t_L g985 ( .A(n_980), .B(n_978), .Y(n_985) );
NAND4xp75_ASAP7_75t_L g986 ( .A(n_982), .B(n_975), .C(n_822), .D(n_859), .Y(n_986) );
NOR2x1_ASAP7_75t_L g987 ( .A(n_985), .B(n_983), .Y(n_987) );
INVx2_ASAP7_75t_SL g988 ( .A(n_984), .Y(n_988) );
NOR2x1_ASAP7_75t_L g989 ( .A(n_987), .B(n_986), .Y(n_989) );
NOR2xp67_ASAP7_75t_L g990 ( .A(n_988), .B(n_849), .Y(n_990) );
INVxp33_ASAP7_75t_L g991 ( .A(n_989), .Y(n_991) );
AO22x2_ASAP7_75t_L g992 ( .A1(n_991), .A2(n_990), .B1(n_868), .B2(n_851), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_992), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_993), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g995 ( .A1(n_994), .A2(n_795), .B1(n_854), .B2(n_865), .Y(n_995) );
OR2x6_ASAP7_75t_L g996 ( .A(n_995), .B(n_900), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_996), .B(n_912), .Y(n_997) );
OR2x6_ASAP7_75t_L g998 ( .A(n_997), .B(n_919), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g999 ( .A1(n_998), .A2(n_836), .B1(n_858), .B2(n_857), .Y(n_999) );
endmodule