module fake_jpeg_18008_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_1),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_63),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_0),
.Y(n_73)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_56),
.Y(n_77)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_65),
.A2(n_49),
.B1(n_45),
.B2(n_61),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_79),
.B1(n_74),
.B2(n_83),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_84),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_31),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_29),
.B(n_39),
.C(n_37),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_78),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_45),
.B1(n_61),
.B2(n_56),
.Y(n_79)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_47),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_97),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_90),
.A2(n_96),
.B1(n_102),
.B2(n_6),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_52),
.B(n_3),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_6),
.C(n_7),
.Y(n_111)
);

AOI22x1_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_48),
.B1(n_57),
.B2(n_62),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_54),
.B1(n_58),
.B2(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_62),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_53),
.B1(n_60),
.B2(n_46),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_50),
.B1(n_57),
.B2(n_5),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_78),
.B1(n_4),
.B2(n_5),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

AND2x4_ASAP7_75t_SL g105 ( 
.A(n_94),
.B(n_2),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_109),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_21),
.C(n_42),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_113),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_102),
.B1(n_98),
.B2(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_7),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_115),
.A2(n_105),
.B(n_108),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_107),
.B1(n_105),
.B2(n_114),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_120),
.A2(n_122),
.B1(n_112),
.B2(n_95),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_115),
.A2(n_111),
.B(n_96),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_117),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_116),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_125),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_118),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_128),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_121),
.B1(n_23),
.B2(n_27),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_20),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_130),
.B(n_126),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_132),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_134),
.A2(n_129),
.B1(n_133),
.B2(n_28),
.Y(n_135)
);

OAI21x1_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_22),
.B(n_43),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_129),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_13),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_103),
.C(n_19),
.Y(n_140)
);

AOI322xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_12),
.A3(n_32),
.B1(n_30),
.B2(n_36),
.C1(n_11),
.C2(n_10),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_8),
.B(n_9),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_9),
.Y(n_143)
);


endmodule