module real_jpeg_22963_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_0),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_0),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_0),
.A2(n_59),
.B1(n_62),
.B2(n_67),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_0),
.A2(n_39),
.B1(n_41),
.B2(n_59),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_0),
.A2(n_26),
.B1(n_33),
.B2(n_59),
.Y(n_209)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_2),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_2),
.B(n_61),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_2),
.B(n_39),
.C(n_83),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_2),
.A2(n_62),
.B1(n_67),
.B2(n_171),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_2),
.B(n_125),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_2),
.A2(n_39),
.B1(n_41),
.B2(n_171),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_2),
.B(n_26),
.C(n_44),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_2),
.A2(n_25),
.B(n_258),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_3),
.A2(n_39),
.B1(n_41),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_3),
.A2(n_26),
.B1(n_33),
.B2(n_48),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_3),
.A2(n_48),
.B1(n_62),
.B2(n_67),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_5),
.A2(n_75),
.B1(n_77),
.B2(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_5),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_5),
.A2(n_62),
.B1(n_67),
.B2(n_147),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_5),
.A2(n_39),
.B1(n_41),
.B2(n_147),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_5),
.A2(n_26),
.B1(n_33),
.B2(n_147),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_8),
.A2(n_57),
.B1(n_77),
.B2(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_8),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_8),
.A2(n_62),
.B1(n_67),
.B2(n_110),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_8),
.A2(n_39),
.B1(n_41),
.B2(n_110),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_8),
.A2(n_26),
.B1(n_33),
.B2(n_110),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_11),
.A2(n_62),
.B1(n_67),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_11),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_11),
.A2(n_39),
.B1(n_41),
.B2(n_87),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_11),
.A2(n_57),
.B1(n_58),
.B2(n_87),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_11),
.A2(n_26),
.B1(n_33),
.B2(n_87),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_13),
.A2(n_38),
.B1(n_62),
.B2(n_67),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_13),
.A2(n_26),
.B1(n_33),
.B2(n_38),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_14),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_14),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_15),
.A2(n_58),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_15),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_15),
.A2(n_62),
.B1(n_67),
.B2(n_72),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_15),
.A2(n_39),
.B1(n_41),
.B2(n_72),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_15),
.A2(n_26),
.B1(n_33),
.B2(n_72),
.Y(n_228)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_16),
.Y(n_100)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_16),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_137),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_135),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_114),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_21),
.B(n_114),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_78),
.C(n_94),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_22),
.A2(n_78),
.B1(n_79),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_22),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_23),
.A2(n_24),
.B(n_52),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_24),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_24),
.A2(n_35),
.B1(n_36),
.B2(n_51),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B(n_32),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_25),
.A2(n_32),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_25),
.A2(n_99),
.B1(n_100),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_25),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_25),
.A2(n_100),
.B1(n_176),
.B2(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_25),
.B(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_25),
.A2(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_26),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_26),
.A2(n_33),
.B1(n_44),
.B2(n_45),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_28),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_28),
.Y(n_281)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_30),
.A2(n_226),
.B(n_227),
.Y(n_225)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_33),
.B(n_285),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_42),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_37),
.A2(n_42),
.B1(n_49),
.B2(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_39),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_39),
.A2(n_41),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_39),
.B(n_266),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_42),
.A2(n_49),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_42),
.B(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_42),
.A2(n_49),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_46),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_46),
.A2(n_90),
.B1(n_104),
.B2(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_46),
.A2(n_157),
.B(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_46),
.A2(n_196),
.B(n_231),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_46),
.B(n_171),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_49),
.B(n_197),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_60),
.B(n_68),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_54),
.A2(n_60),
.B1(n_111),
.B2(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp33_ASAP7_75t_SL g170 ( 
.A(n_56),
.B(n_171),
.Y(n_170)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_SL g199 ( 
.A1(n_58),
.A2(n_170),
.B(n_171),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_70),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_60),
.A2(n_68),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_61),
.A2(n_73),
.B1(n_109),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_61)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_67),
.B1(n_83),
.B2(n_84),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_62),
.A2(n_66),
.B(n_170),
.C(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_62),
.B(n_224),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_66),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_SL g172 ( 
.A(n_65),
.B(n_67),
.C(n_77),
.Y(n_172)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_73),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_73),
.A2(n_113),
.B(n_199),
.Y(n_198)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_89),
.B(n_93),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_89),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_88),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_81),
.A2(n_164),
.B(n_166),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_81),
.A2(n_166),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_82),
.A2(n_106),
.B(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_82),
.A2(n_150),
.B(n_205),
.Y(n_204)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_88),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_90),
.A2(n_245),
.B(n_246),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_90),
.A2(n_246),
.B(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_92),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_94),
.A2(n_95),
.B1(n_315),
.B2(n_317),
.Y(n_314)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_105),
.C(n_107),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_96),
.A2(n_97),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_98),
.A2(n_101),
.B1(n_102),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_98),
.Y(n_159)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_100),
.Y(n_177)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_100),
.Y(n_287)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_105),
.B(n_107),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B(n_112),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_132),
.B2(n_134),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_128),
.B1(n_129),
.B2(n_131),
.Y(n_121)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_124),
.A2(n_125),
.B1(n_165),
.B2(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_125),
.B(n_151),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_132),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_313),
.B(n_319),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_185),
.B(n_312),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_178),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_140),
.B(n_178),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_158),
.C(n_160),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_141),
.A2(n_142),
.B1(n_158),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_152),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_148),
.C(n_152),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_153),
.B(n_156),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_174),
.B1(n_175),
.B2(n_177),
.Y(n_173)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_158),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_160),
.B(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.C(n_167),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_163),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_167),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_173),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_168),
.A2(n_169),
.B1(n_173),
.B2(n_202),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_171),
.B(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_174),
.A2(n_270),
.B1(n_272),
.B2(n_274),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_184),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_180),
.B(n_181),
.C(n_184),
.Y(n_318)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_216),
.B(n_306),
.C(n_311),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_210),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_210),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_200),
.C(n_203),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_188),
.A2(n_189),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_198),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_194),
.C(n_198),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_193),
.Y(n_205)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_203),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.C(n_208),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_211),
.B(n_214),
.C(n_215),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_299),
.B(n_305),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_247),
.B(n_298),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_236),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_221),
.B(n_236),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_229),
.C(n_233),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_222),
.B(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_225),
.Y(n_243)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_227),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_228),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_229),
.A2(n_233),
.B1(n_234),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_229),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_232),
.Y(n_245)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_241),
.B2(n_242),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_237),
.B(n_243),
.C(n_244),
.Y(n_304)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_292),
.B(n_297),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_267),
.B(n_291),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_261),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_261),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_256),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_252),
.B(n_255),
.C(n_256),
.Y(n_296)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_277),
.B(n_290),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_275),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_275),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_281),
.B(n_282),
.Y(n_280)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_283),
.B(n_289),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_280),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_288),
.Y(n_283)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_296),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_304),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_304),
.Y(n_305)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_318),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_318),
.Y(n_319)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_315),
.Y(n_317)
);


endmodule