module real_jpeg_27208_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_200;
wire n_48;
wire n_56;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_0),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_0),
.A2(n_23),
.B1(n_26),
.B2(n_45),
.Y(n_53)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_1),
.B(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_1),
.B(n_184),
.Y(n_189)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_1),
.Y(n_200)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_4),
.A2(n_23),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_4),
.A2(n_33),
.B1(n_42),
.B2(n_43),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_4),
.A2(n_6),
.B1(n_33),
.B2(n_64),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_4),
.A2(n_33),
.B1(n_68),
.B2(n_69),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_5),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_5),
.A2(n_25),
.B1(n_42),
.B2(n_43),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_5),
.A2(n_25),
.B1(n_68),
.B2(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_5),
.B(n_64),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_5),
.A2(n_64),
.B(n_107),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_5),
.A2(n_10),
.B(n_43),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_5),
.B(n_93),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_5),
.A2(n_7),
.B(n_23),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_5),
.B(n_85),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_6),
.A2(n_8),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_8),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_8),
.A2(n_65),
.B1(n_68),
.B2(n_69),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_65),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_8),
.A2(n_23),
.B1(n_26),
.B2(n_65),
.Y(n_184)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_131),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_130),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_112),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_16),
.B(n_112),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_89),
.B2(n_111),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_50),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_29),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_21),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_22),
.A2(n_27),
.B(n_35),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_22),
.B(n_35),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_23),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_23),
.A2(n_26),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_25),
.A2(n_69),
.B(n_82),
.C(n_140),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_25),
.A2(n_39),
.B(n_43),
.C(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_25),
.B(n_37),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_25),
.B(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_26),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_27),
.B(n_32),
.Y(n_54)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_27),
.Y(n_110)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_29),
.A2(n_53),
.B(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_30),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_53),
.B(n_54),
.Y(n_52)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_35),
.B(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B(n_46),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_37),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_49),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_38),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_38),
.B(n_58),
.Y(n_165)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_42),
.A2(n_43),
.B1(n_83),
.B2(n_84),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_46),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_47),
.B(n_150),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_59),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_52),
.B(n_55),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_54),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_54),
.B(n_183),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_56),
.B(n_166),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_57),
.B(n_149),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_58),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_76),
.B2(n_77),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_72),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_62),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_63),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_66),
.B(n_67),
.C(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_66)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_71),
.Y(n_105)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_80),
.B(n_81),
.C(n_85),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_69),
.B(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_69),
.A2(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_74),
.B(n_120),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_86),
.B(n_87),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_79),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_79),
.B(n_88),
.Y(n_146)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_85),
.B(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_85),
.B(n_129),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_98),
.C(n_103),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_91),
.B1(n_98),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_101),
.B(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_103),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_104),
.B(n_109),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.C(n_117),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_113),
.B(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_116),
.B(n_117),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.C(n_125),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_118),
.B(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_126),
.Y(n_214)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_227),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_223),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_210),
.B(n_222),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_168),
.B(n_209),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_151),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_137),
.B(n_151),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_144),
.C(n_147),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_138),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_139),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_142),
.Y(n_167)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_207)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_162),
.B2(n_163),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_152),
.B(n_164),
.C(n_167),
.Y(n_211)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_154),
.B(n_157),
.C(n_160),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_189),
.Y(n_197)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_204),
.B(n_208),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_185),
.B(n_203),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_171),
.B(n_176),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_174),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_182),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_181),
.C(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_192),
.B(n_202),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_187),
.B(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_196),
.B(n_201),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_194),
.B(n_195),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_205),
.B(n_206),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_211),
.B(n_212),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_215),
.B1(n_216),
.B2(n_221),
.Y(n_212)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_220),
.C(n_221),
.Y(n_224)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_225),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);


endmodule