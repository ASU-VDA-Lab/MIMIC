module fake_jpeg_26936_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_59),
.Y(n_88)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_45),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_95),
.B(n_50),
.Y(n_105)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_74),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_19),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_76),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_28),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_44),
.B1(n_48),
.B2(n_17),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_91),
.B1(n_52),
.B2(n_60),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_34),
.B1(n_17),
.B2(n_18),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_47),
.C(n_46),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_25),
.C(n_39),
.Y(n_113)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_86),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_30),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_34),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_71),
.Y(n_102)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_44),
.B1(n_17),
.B2(n_40),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_66),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

CKINVDCx12_ASAP7_75t_R g93 ( 
.A(n_61),
.Y(n_93)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_34),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_56),
.A2(n_18),
.B1(n_35),
.B2(n_28),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_85),
.B1(n_97),
.B2(n_35),
.Y(n_126)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_78),
.A2(n_44),
.B1(n_55),
.B2(n_52),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_99),
.A2(n_90),
.B1(n_80),
.B2(n_84),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_107),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_66),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_91),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_55),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_18),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_87),
.B1(n_22),
.B2(n_35),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_24),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_77),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_25),
.C(n_77),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_25),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_116),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_29),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_69),
.A2(n_35),
.B1(n_22),
.B2(n_27),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_31),
.B1(n_32),
.B2(n_85),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_73),
.B(n_29),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_116),
.Y(n_148)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_100),
.B(n_30),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_131),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_132),
.A2(n_36),
.B1(n_32),
.B2(n_83),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_137),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_143),
.B(n_108),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_127),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_145),
.B1(n_154),
.B2(n_123),
.Y(n_157)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_102),
.B(n_26),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_144),
.Y(n_172)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_77),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_148),
.Y(n_179)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

BUFx12_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_114),
.B(n_26),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_21),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_104),
.A2(n_36),
.B1(n_26),
.B2(n_31),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_108),
.C(n_109),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_124),
.B1(n_122),
.B2(n_113),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_156),
.A2(n_171),
.B1(n_176),
.B2(n_183),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_157),
.A2(n_159),
.B(n_169),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_100),
.A3(n_103),
.B1(n_105),
.B2(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_161),
.B(n_177),
.C(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_162),
.B(n_163),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_120),
.B1(n_111),
.B2(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_164),
.B(n_173),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_143),
.B(n_134),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_130),
.A2(n_112),
.B1(n_125),
.B2(n_119),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g174 ( 
.A1(n_135),
.A2(n_115),
.B(n_101),
.Y(n_174)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_112),
.B1(n_123),
.B2(n_115),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_175),
.A2(n_186),
.B1(n_142),
.B2(n_149),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_136),
.A2(n_98),
.B1(n_21),
.B2(n_25),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_101),
.C(n_98),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_140),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_178),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_151),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_181),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_141),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_145),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_83),
.C(n_94),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_33),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_147),
.A2(n_42),
.B1(n_33),
.B2(n_25),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_151),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_161),
.C(n_177),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_193),
.Y(n_241)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_133),
.Y(n_195)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_181),
.B(n_128),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_196),
.Y(n_239)
);

NOR2x1_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_134),
.Y(n_197)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_198),
.B(n_206),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_144),
.Y(n_199)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_200),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_154),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_209),
.B(n_215),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_216),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_167),
.B(n_137),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_153),
.Y(n_207)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_162),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_129),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_164),
.B(n_143),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_211),
.Y(n_221)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_213),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_170),
.B(n_148),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_170),
.B(n_132),
.Y(n_214)
);

INVxp33_ASAP7_75t_SL g234 ( 
.A(n_214),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_166),
.B(n_150),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_149),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_217),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_219),
.B(n_197),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_173),
.C(n_159),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_198),
.C(n_215),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_193),
.A2(n_169),
.B1(n_174),
.B2(n_166),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_222),
.A2(n_227),
.B1(n_232),
.B2(n_200),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_188),
.A2(n_174),
.B1(n_183),
.B2(n_178),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_225),
.A2(n_229),
.B1(n_211),
.B2(n_205),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_189),
.A2(n_182),
.B1(n_160),
.B2(n_180),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_188),
.A2(n_186),
.B1(n_160),
.B2(n_142),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_210),
.A2(n_150),
.B(n_24),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_231),
.A2(n_235),
.B(n_237),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_189),
.A2(n_150),
.B1(n_72),
.B2(n_33),
.Y(n_232)
);

NAND2x1_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_94),
.Y(n_235)
);

OAI22x1_ASAP7_75t_L g237 ( 
.A1(n_197),
.A2(n_94),
.B1(n_24),
.B2(n_2),
.Y(n_237)
);

AOI21xp33_ASAP7_75t_L g238 ( 
.A1(n_194),
.A2(n_8),
.B(n_15),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_238),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_239),
.B(n_192),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_245),
.B(n_252),
.Y(n_279)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_256),
.B1(n_222),
.B2(n_233),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_220),
.B(n_190),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_248),
.B(n_264),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_194),
.Y(n_249)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_233),
.A2(n_212),
.B(n_210),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_208),
.Y(n_251)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_251),
.Y(n_284)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

AO22x1_ASAP7_75t_L g282 ( 
.A1(n_254),
.A2(n_229),
.B1(n_218),
.B2(n_224),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_199),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_258),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_204),
.B1(n_218),
.B2(n_205),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_195),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_261),
.C(n_263),
.Y(n_267)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_202),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_262),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_235),
.A2(n_201),
.B1(n_187),
.B2(n_204),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_227),
.B(n_207),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_265),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_201),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_242),
.C(n_228),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_221),
.C(n_242),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_275),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_278),
.B1(n_283),
.B2(n_254),
.Y(n_288)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_261),
.C(n_253),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_235),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_231),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_236),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_247),
.A2(n_232),
.B1(n_237),
.B2(n_243),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_246),
.Y(n_280)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_282),
.B(n_265),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_260),
.A2(n_243),
.B1(n_187),
.B2(n_226),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_279),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_294),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_284),
.B(n_271),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_282),
.B1(n_281),
.B2(n_274),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_266),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_289),
.B(n_297),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_293),
.C(n_300),
.Y(n_306)
);

INVxp33_ASAP7_75t_SL g291 ( 
.A(n_280),
.Y(n_291)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_262),
.C(n_249),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_277),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_270),
.A2(n_253),
.B(n_224),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_296),
.A2(n_274),
.B1(n_9),
.B2(n_10),
.Y(n_305)
);

OAI21xp33_ASAP7_75t_L g297 ( 
.A1(n_275),
.A2(n_250),
.B(n_236),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_298),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_299),
.B(n_6),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_217),
.C(n_236),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_308),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_307),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_292),
.A2(n_7),
.B1(n_15),
.B2(n_13),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_7),
.B1(n_15),
.B2(n_13),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_6),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_300),
.C(n_290),
.Y(n_314)
);

XNOR2x1_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_313),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_0),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_297),
.B1(n_293),
.B2(n_289),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_10),
.B1(n_11),
.B2(n_2),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_309),
.A2(n_285),
.B(n_9),
.Y(n_316)
);

AOI21xp33_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_321),
.B(n_311),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_16),
.C(n_5),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_319),
.C(n_313),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_13),
.C(n_12),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_301),
.A2(n_10),
.B(n_11),
.Y(n_321)
);

OAI21x1_ASAP7_75t_L g323 ( 
.A1(n_317),
.A2(n_312),
.B(n_311),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_325),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_324),
.A2(n_322),
.B(n_3),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_317),
.A2(n_304),
.B1(n_310),
.B2(n_11),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_327),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_329),
.C(n_1),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_320),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_330),
.A2(n_331),
.B(n_328),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

BUFx12f_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_332),
.B(n_333),
.C(n_325),
.Y(n_337)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_337),
.Y(n_338)
);

OAI211xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_336),
.B(n_3),
.C(n_4),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_3),
.Y(n_340)
);


endmodule