module fake_jpeg_15961_n_152 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_2),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_21),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_71),
.Y(n_72)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_1),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_53),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_61),
.B1(n_49),
.B2(n_58),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_83),
.B1(n_84),
.B2(n_57),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_61),
.B1(n_49),
.B2(n_55),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_44),
.B1(n_60),
.B2(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_50),
.B1(n_47),
.B2(n_56),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_92),
.Y(n_114)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_83),
.B(n_84),
.C(n_42),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_1),
.Y(n_94)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_2),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_3),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_4),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_72),
.B(n_62),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_4),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_5),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_48),
.C(n_54),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_106),
.A2(n_42),
.B1(n_57),
.B2(n_8),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_93),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_113),
.A2(n_94),
.B1(n_9),
.B2(n_10),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_114),
.A2(n_105),
.B1(n_91),
.B2(n_102),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_120),
.B1(n_121),
.B2(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_123),
.B(n_115),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_124),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_115),
.B(n_116),
.C(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_116),
.Y(n_129)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_132),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_136),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_134),
.A2(n_128),
.B1(n_130),
.B2(n_132),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_126),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_133),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_138),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_133),
.B(n_123),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_111),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_32),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_93),
.C(n_13),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_SL g146 ( 
.A(n_145),
.B(n_31),
.C(n_15),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_146),
.A2(n_33),
.B(n_16),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_34),
.C(n_18),
.Y(n_148)
);

OAI321xp33_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_35),
.A3(n_19),
.B1(n_22),
.B2(n_25),
.C(n_26),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_37),
.B(n_28),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_38),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_107),
.B1(n_29),
.B2(n_30),
.Y(n_152)
);


endmodule