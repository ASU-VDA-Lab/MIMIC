module fake_jpeg_11294_n_238 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_238);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_238;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_18),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

CKINVDCx9p33_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_23),
.A2(n_27),
.B1(n_20),
.B2(n_31),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_34),
.B1(n_20),
.B2(n_31),
.Y(n_74)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_34),
.B1(n_32),
.B2(n_28),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_62),
.B1(n_75),
.B2(n_80),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_20),
.B1(n_27),
.B2(n_31),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_61),
.A2(n_26),
.B1(n_22),
.B2(n_25),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_34),
.B1(n_32),
.B2(n_28),
.Y(n_62)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_71),
.B(n_79),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_44),
.B1(n_51),
.B2(n_52),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_28),
.B1(n_27),
.B2(n_29),
.Y(n_75)
);

NOR2x1_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_30),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_12),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_39),
.C(n_43),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_53),
.A2(n_28),
.B1(n_21),
.B2(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_17),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_30),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_86),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_88),
.B(n_99),
.Y(n_135)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_89),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_104),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_91),
.A2(n_92),
.B1(n_108),
.B2(n_72),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_26),
.B1(n_22),
.B2(n_45),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_102),
.B1(n_56),
.B2(n_67),
.Y(n_125)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_75),
.A2(n_25),
.B1(n_54),
.B2(n_36),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_2),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_114),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_65),
.A2(n_66),
.B1(n_64),
.B2(n_69),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_56),
.A2(n_50),
.B1(n_3),
.B2(n_5),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_13),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_111),
.B(n_116),
.Y(n_131)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_78),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_2),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_13),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_69),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_64),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_136),
.B1(n_113),
.B2(n_104),
.Y(n_146)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_73),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_127),
.B(n_7),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_129),
.B1(n_112),
.B2(n_115),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_57),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_106),
.C(n_95),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_78),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_134),
.B(n_106),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_90),
.A2(n_85),
.B1(n_86),
.B2(n_6),
.Y(n_136)
);

OAI31xp33_ASAP7_75t_L g137 ( 
.A1(n_88),
.A2(n_2),
.A3(n_3),
.B(n_6),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_7),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_142),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_91),
.B1(n_94),
.B2(n_126),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_129),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_151),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_133),
.A2(n_108),
.B1(n_102),
.B2(n_110),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_95),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_161),
.C(n_119),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_105),
.Y(n_152)
);

XNOR2x1_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_156),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_135),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_89),
.Y(n_157)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_158),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_87),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_101),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_107),
.Y(n_162)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_163),
.Y(n_171)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_166),
.A2(n_145),
.B1(n_148),
.B2(n_157),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_162),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_167),
.B(n_177),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_152),
.A2(n_137),
.B(n_136),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_164),
.B(n_161),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_151),
.A2(n_131),
.B(n_132),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_174),
.A2(n_181),
.B(n_144),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_158),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_170),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_143),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_120),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_132),
.B(n_138),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_124),
.C(n_139),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_156),
.C(n_154),
.Y(n_187)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_142),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_186),
.B(n_193),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_198),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_188),
.A2(n_196),
.B(n_166),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_180),
.B1(n_183),
.B2(n_178),
.Y(n_207)
);

OAI321xp33_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_148),
.A3(n_155),
.B1(n_165),
.B2(n_139),
.C(n_124),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_195),
.A3(n_192),
.B1(n_173),
.B2(n_172),
.C1(n_191),
.C2(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_194),
.Y(n_201)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

AOI221xp5_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_120),
.B1(n_144),
.B2(n_9),
.C(n_11),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_123),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_199),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_209),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_198),
.B(n_170),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_208),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_210),
.B1(n_188),
.B2(n_196),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_187),
.B(n_182),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_197),
.A2(n_182),
.B(n_174),
.C(n_168),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_201),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_213),
.Y(n_223)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_190),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_214),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_215),
.B(n_218),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_185),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_217),
.A2(n_203),
.B(n_8),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_189),
.C(n_173),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_171),
.C(n_93),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_219),
.B(n_208),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_214),
.A2(n_202),
.B1(n_207),
.B2(n_205),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_217),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_224),
.B(n_212),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_SL g230 ( 
.A1(n_225),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_230)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_223),
.B(n_219),
.CI(n_218),
.CON(n_226),
.SN(n_226)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_229),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_228),
.Y(n_234)
);

A2O1A1O1Ixp25_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_216),
.B(n_212),
.C(n_9),
.D(n_11),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_230),
.A2(n_222),
.B(n_220),
.Y(n_231)
);

OAI21x1_ASAP7_75t_L g236 ( 
.A1(n_231),
.A2(n_232),
.B(n_11),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_93),
.B(n_96),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_230),
.C(n_96),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_236),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_234),
.Y(n_238)
);


endmodule