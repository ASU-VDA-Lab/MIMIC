module fake_netlist_1_1995_n_610 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_610);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_610;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g75 ( .A(n_53), .Y(n_75) );
CKINVDCx20_ASAP7_75t_R g76 ( .A(n_3), .Y(n_76) );
INVx2_ASAP7_75t_SL g77 ( .A(n_18), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_23), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_54), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_16), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_36), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_41), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_42), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_21), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_64), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_45), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_63), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_72), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_65), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_5), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_7), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_34), .Y(n_92) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_21), .Y(n_93) );
INVxp67_ASAP7_75t_L g94 ( .A(n_19), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_47), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_46), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_40), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_17), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_19), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_16), .Y(n_100) );
BUFx2_ASAP7_75t_L g101 ( .A(n_58), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_73), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_9), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_4), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_4), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_27), .Y(n_106) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_14), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_44), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_1), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_24), .Y(n_110) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_5), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_61), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_59), .Y(n_113) );
INVxp33_ASAP7_75t_L g114 ( .A(n_31), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_3), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_0), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_29), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_17), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_75), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_75), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_79), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_79), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_81), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_81), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_87), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_87), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_83), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_101), .B(n_0), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_89), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_89), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_95), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_92), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_110), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_95), .Y(n_134) );
BUFx2_ASAP7_75t_L g135 ( .A(n_111), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_96), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_101), .B(n_1), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_96), .Y(n_138) );
INVx4_ASAP7_75t_L g139 ( .A(n_112), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_109), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_97), .Y(n_141) );
AND2x2_ASAP7_75t_SL g142 ( .A(n_97), .B(n_106), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_106), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_108), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_108), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_117), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_117), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_112), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_105), .B(n_2), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_109), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_114), .B(n_2), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_84), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_84), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_93), .Y(n_154) );
OR2x2_ASAP7_75t_L g155 ( .A(n_107), .B(n_6), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_93), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_94), .B(n_6), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_135), .B(n_100), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_120), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_120), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_120), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_128), .B(n_77), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_123), .Y(n_163) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_123), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_128), .B(n_77), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
NOR2xp33_ASAP7_75t_SL g168 ( .A(n_142), .B(n_86), .Y(n_168) );
OAI22xp5_ASAP7_75t_L g169 ( .A1(n_142), .A2(n_118), .B1(n_116), .B2(n_91), .Y(n_169) );
NAND2x1p5_ASAP7_75t_L g170 ( .A(n_128), .B(n_118), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_123), .Y(n_171) );
INVxp67_ASAP7_75t_SL g172 ( .A(n_155), .Y(n_172) );
INVxp67_ASAP7_75t_SL g173 ( .A(n_155), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_154), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_140), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_142), .B(n_116), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_148), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_150), .B(n_102), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_119), .B(n_113), .Y(n_180) );
INVx5_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_154), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_134), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_119), .B(n_78), .Y(n_184) );
INVxp67_ASAP7_75t_L g185 ( .A(n_151), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_127), .Y(n_186) );
AND2x6_ASAP7_75t_L g187 ( .A(n_151), .B(n_93), .Y(n_187) );
NAND2x1p5_ASAP7_75t_L g188 ( .A(n_121), .B(n_91), .Y(n_188) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_121), .A2(n_85), .B(n_88), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_134), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_148), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_154), .Y(n_192) );
CKINVDCx16_ASAP7_75t_R g193 ( .A(n_137), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_139), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_138), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_122), .B(n_82), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_138), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_138), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_147), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_147), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_147), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_131), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_131), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_154), .Y(n_204) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_122), .A2(n_98), .B(n_104), .Y(n_205) );
INVx4_ASAP7_75t_L g206 ( .A(n_187), .Y(n_206) );
INVx4_ASAP7_75t_SL g207 ( .A(n_187), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_159), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_172), .B(n_124), .Y(n_209) );
BUFx2_ASAP7_75t_L g210 ( .A(n_164), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_168), .A2(n_130), .B1(n_124), .B2(n_125), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_159), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_173), .B(n_125), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_161), .Y(n_214) );
NAND2xp33_ASAP7_75t_SL g215 ( .A(n_167), .B(n_132), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_186), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_185), .B(n_126), .Y(n_217) );
INVx1_ASAP7_75t_SL g218 ( .A(n_193), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_176), .B(n_167), .Y(n_219) );
INVx1_ASAP7_75t_SL g220 ( .A(n_175), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_167), .B(n_126), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_161), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_163), .Y(n_223) );
INVx2_ASAP7_75t_SL g224 ( .A(n_187), .Y(n_224) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_170), .Y(n_225) );
BUFx2_ASAP7_75t_L g226 ( .A(n_187), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_163), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_170), .B(n_129), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_170), .B(n_129), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_177), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_171), .Y(n_231) );
NOR3xp33_ASAP7_75t_SL g232 ( .A(n_186), .B(n_133), .C(n_149), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_162), .B(n_130), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_177), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_191), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_176), .B(n_136), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_162), .B(n_136), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_188), .B(n_141), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_191), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_160), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_162), .B(n_141), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_160), .Y(n_242) );
BUFx2_ASAP7_75t_L g243 ( .A(n_187), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_171), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_166), .B(n_143), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_166), .B(n_144), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_169), .A2(n_157), .B1(n_143), .B2(n_144), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_166), .A2(n_145), .B1(n_146), .B2(n_98), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_187), .Y(n_249) );
BUFx2_ASAP7_75t_L g250 ( .A(n_187), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_178), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_188), .B(n_184), .Y(n_252) );
INVx4_ASAP7_75t_L g253 ( .A(n_181), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_178), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_183), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_183), .Y(n_256) );
NOR2x1_ASAP7_75t_L g257 ( .A(n_205), .B(n_145), .Y(n_257) );
BUFx4f_ASAP7_75t_L g258 ( .A(n_188), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_190), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_196), .B(n_139), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_190), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_180), .B(n_139), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_158), .A2(n_146), .B1(n_80), .B2(n_90), .Y(n_263) );
NOR3xp33_ASAP7_75t_SL g264 ( .A(n_179), .B(n_115), .C(n_104), .Y(n_264) );
BUFx3_ASAP7_75t_L g265 ( .A(n_258), .Y(n_265) );
AOI211xp5_ASAP7_75t_L g266 ( .A1(n_218), .A2(n_103), .B(n_80), .C(n_99), .Y(n_266) );
INVx1_ASAP7_75t_SL g267 ( .A(n_210), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_210), .B(n_205), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_258), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_220), .B(n_205), .Y(n_270) );
INVx1_ASAP7_75t_SL g271 ( .A(n_238), .Y(n_271) );
OA21x2_ASAP7_75t_L g272 ( .A1(n_208), .A2(n_199), .B(n_201), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_238), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_236), .B(n_209), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_219), .B(n_202), .Y(n_275) );
AOI22xp33_ASAP7_75t_SL g276 ( .A1(n_216), .A2(n_76), .B1(n_189), .B2(n_99), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_258), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_211), .A2(n_197), .B1(n_201), .B2(n_200), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_246), .Y(n_279) );
INVx5_ASAP7_75t_L g280 ( .A(n_206), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_225), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_234), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_216), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_246), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_246), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_236), .B(n_202), .Y(n_286) );
OAI221xp5_ASAP7_75t_L g287 ( .A1(n_264), .A2(n_203), .B1(n_90), .B2(n_103), .C(n_197), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_232), .Y(n_288) );
OAI21xp5_ASAP7_75t_L g289 ( .A1(n_257), .A2(n_189), .B(n_194), .Y(n_289) );
NAND2x1p5_ASAP7_75t_L g290 ( .A(n_206), .B(n_198), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_213), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_219), .Y(n_292) );
INVx3_ASAP7_75t_SL g293 ( .A(n_207), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_217), .B(n_203), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_221), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_251), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_219), .A2(n_189), .B1(n_200), .B2(n_199), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_252), .B(n_194), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_263), .B(n_189), .Y(n_299) );
BUFx3_ASAP7_75t_L g300 ( .A(n_234), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_251), .Y(n_301) );
AOI222xp33_ASAP7_75t_L g302 ( .A1(n_233), .A2(n_152), .B1(n_153), .B2(n_195), .C1(n_160), .C2(n_165), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_255), .B(n_165), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_253), .Y(n_304) );
INVx4_ASAP7_75t_L g305 ( .A(n_206), .Y(n_305) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_237), .A2(n_152), .B1(n_153), .B2(n_195), .C(n_165), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_211), .A2(n_198), .B1(n_148), .B2(n_181), .Y(n_307) );
OR2x6_ASAP7_75t_L g308 ( .A(n_249), .B(n_93), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_228), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_229), .B(n_198), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_249), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_226), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_226), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_241), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_245), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_243), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_255), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_272), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_291), .B(n_248), .Y(n_319) );
CKINVDCx16_ASAP7_75t_R g320 ( .A(n_267), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_265), .B(n_207), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_294), .A2(n_248), .B1(n_214), .B2(n_244), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_305), .Y(n_323) );
OAI22xp33_ASAP7_75t_L g324 ( .A1(n_271), .A2(n_247), .B1(n_227), .B2(n_208), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_289), .A2(n_260), .B(n_257), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_SL g326 ( .A1(n_296), .A2(n_214), .B(n_223), .C(n_222), .Y(n_326) );
INVx5_ASAP7_75t_L g327 ( .A(n_308), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_272), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_272), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_283), .Y(n_330) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_287), .A2(n_231), .B(n_227), .C(n_223), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_314), .B(n_212), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_315), .B(n_212), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_273), .B(n_256), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_276), .A2(n_215), .B1(n_222), .B2(n_254), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_274), .B(n_256), .Y(n_336) );
NAND3xp33_ASAP7_75t_L g337 ( .A(n_266), .B(n_234), .C(n_235), .Y(n_337) );
XOR2xp5_ASAP7_75t_L g338 ( .A(n_283), .B(n_243), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_309), .B(n_259), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_292), .A2(n_268), .B1(n_275), .B2(n_270), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_308), .Y(n_341) );
AOI22xp33_ASAP7_75t_SL g342 ( .A1(n_268), .A2(n_254), .B1(n_244), .B2(n_231), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_280), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_270), .A2(n_295), .B1(n_302), .B2(n_292), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_296), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_275), .B(n_259), .Y(n_346) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_299), .A2(n_261), .B(n_230), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_265), .B(n_207), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_275), .A2(n_240), .B1(n_242), .B2(n_250), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_294), .B(n_261), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_279), .A2(n_240), .B1(n_242), .B2(n_250), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_343), .Y(n_352) );
OAI221xp5_ASAP7_75t_SL g353 ( .A1(n_335), .A2(n_299), .B1(n_286), .B2(n_306), .C(n_297), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_345), .Y(n_354) );
OAI221xp5_ASAP7_75t_L g355 ( .A1(n_344), .A2(n_285), .B1(n_284), .B2(n_288), .C(n_281), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_318), .Y(n_356) );
OAI221xp5_ASAP7_75t_L g357 ( .A1(n_344), .A2(n_288), .B1(n_269), .B2(n_278), .C(n_298), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_319), .B(n_269), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_324), .A2(n_93), .B1(n_307), .B2(n_303), .C(n_317), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_322), .A2(n_317), .B1(n_301), .B2(n_308), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_350), .B(n_301), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_324), .A2(n_303), .B1(n_93), .B2(n_312), .Y(n_362) );
OAI221xp5_ASAP7_75t_L g363 ( .A1(n_335), .A2(n_277), .B1(n_310), .B2(n_240), .C(n_242), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_343), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g365 ( .A1(n_325), .A2(n_239), .B(n_230), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_318), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_345), .Y(n_367) );
OAI21x1_ASAP7_75t_L g368 ( .A1(n_347), .A2(n_290), .B(n_304), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_343), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_318), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_340), .B(n_277), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_329), .Y(n_372) );
OA21x2_ASAP7_75t_L g373 ( .A1(n_347), .A2(n_156), .B(n_239), .Y(n_373) );
A2O1A1Ixp33_ASAP7_75t_L g374 ( .A1(n_331), .A2(n_304), .B(n_313), .C(n_224), .Y(n_374) );
OAI22xp5_ASAP7_75t_SL g375 ( .A1(n_320), .A2(n_308), .B1(n_312), .B2(n_316), .Y(n_375) );
AOI222xp33_ASAP7_75t_L g376 ( .A1(n_322), .A2(n_316), .B1(n_207), .B2(n_313), .C1(n_304), .C2(n_305), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_329), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_350), .A2(n_300), .B1(n_235), .B2(n_234), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_329), .Y(n_379) );
OAI321xp33_ASAP7_75t_L g380 ( .A1(n_355), .A2(n_337), .A3(n_319), .B1(n_328), .B2(n_331), .C(n_332), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_356), .Y(n_381) );
OAI33xp33_ASAP7_75t_L g382 ( .A1(n_360), .A2(n_337), .A3(n_156), .B1(n_328), .B2(n_332), .B3(n_333), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_368), .A2(n_347), .B(n_325), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_354), .B(n_336), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_355), .A2(n_342), .B1(n_336), .B2(n_320), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_361), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_361), .Y(n_387) );
INVx4_ASAP7_75t_L g388 ( .A(n_352), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_354), .B(n_342), .Y(n_389) );
NOR3xp33_ASAP7_75t_L g390 ( .A(n_357), .B(n_333), .C(n_346), .Y(n_390) );
OAI221xp5_ASAP7_75t_SL g391 ( .A1(n_362), .A2(n_338), .B1(n_346), .B2(n_334), .C(n_339), .Y(n_391) );
OAI221xp5_ASAP7_75t_L g392 ( .A1(n_357), .A2(n_359), .B1(n_362), .B2(n_353), .C(n_363), .Y(n_392) );
NAND2xp33_ASAP7_75t_R g393 ( .A(n_373), .B(n_341), .Y(n_393) );
NOR3xp33_ASAP7_75t_SL g394 ( .A(n_358), .B(n_330), .C(n_262), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_359), .A2(n_334), .B1(n_339), .B2(n_338), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_367), .B(n_341), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_370), .B(n_323), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_352), .B(n_323), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_352), .B(n_323), .Y(n_399) );
AND2x2_ASAP7_75t_SL g400 ( .A(n_379), .B(n_321), .Y(n_400) );
AO22x1_ASAP7_75t_L g401 ( .A1(n_360), .A2(n_370), .B1(n_379), .B2(n_377), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_356), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_356), .Y(n_403) );
AOI222xp33_ASAP7_75t_L g404 ( .A1(n_375), .A2(n_327), .B1(n_323), .B2(n_349), .C1(n_348), .C2(n_321), .Y(n_404) );
OR2x6_ASAP7_75t_L g405 ( .A(n_375), .B(n_321), .Y(n_405) );
AND2x4_ASAP7_75t_SL g406 ( .A(n_369), .B(n_321), .Y(n_406) );
A2O1A1Ixp33_ASAP7_75t_L g407 ( .A1(n_363), .A2(n_327), .B(n_351), .C(n_348), .Y(n_407) );
AOI31xp33_ASAP7_75t_L g408 ( .A1(n_371), .A2(n_348), .A3(n_326), .B(n_290), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_366), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_358), .B(n_348), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_402), .B(n_366), .Y(n_411) );
INVx2_ASAP7_75t_SL g412 ( .A(n_388), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_381), .B(n_366), .Y(n_413) );
OAI21xp33_ASAP7_75t_L g414 ( .A1(n_391), .A2(n_353), .B(n_376), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_384), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_384), .B(n_372), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_381), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_392), .A2(n_371), .B1(n_376), .B2(n_369), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_381), .Y(n_419) );
INVx2_ASAP7_75t_SL g420 ( .A(n_388), .Y(n_420) );
OAI211xp5_ASAP7_75t_L g421 ( .A1(n_385), .A2(n_371), .B(n_378), .C(n_364), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_403), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_386), .B(n_372), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_403), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_403), .B(n_372), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_409), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_387), .B(n_377), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_409), .B(n_377), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_409), .B(n_373), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_388), .B(n_368), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_397), .B(n_373), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_397), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_389), .Y(n_433) );
NOR3xp33_ASAP7_75t_L g434 ( .A(n_391), .B(n_364), .C(n_369), .Y(n_434) );
NOR3xp33_ASAP7_75t_L g435 ( .A(n_380), .B(n_364), .C(n_369), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_388), .B(n_368), .Y(n_436) );
OAI21xp5_ASAP7_75t_SL g437 ( .A1(n_408), .A2(n_378), .B(n_374), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_389), .B(n_373), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_396), .B(n_373), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_396), .B(n_365), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_401), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_400), .B(n_365), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_400), .B(n_7), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_400), .B(n_8), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_392), .A2(n_154), .B1(n_224), .B2(n_182), .C(n_192), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_390), .B(n_8), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_395), .A2(n_327), .B1(n_300), .B2(n_282), .Y(n_447) );
NOR2xp33_ASAP7_75t_SL g448 ( .A(n_382), .B(n_327), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_398), .B(n_9), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_398), .B(n_10), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_398), .B(n_10), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_401), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_398), .B(n_11), .Y(n_453) );
AND2x4_ASAP7_75t_SL g454 ( .A(n_449), .B(n_405), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_414), .A2(n_408), .B1(n_405), .B2(n_407), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_415), .B(n_405), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_433), .B(n_383), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_433), .B(n_405), .Y(n_458) );
NAND2xp33_ASAP7_75t_R g459 ( .A(n_430), .B(n_394), .Y(n_459) );
OAI31xp33_ASAP7_75t_L g460 ( .A1(n_414), .A2(n_446), .A3(n_444), .B(n_443), .Y(n_460) );
NAND4xp25_ASAP7_75t_L g461 ( .A(n_418), .B(n_404), .C(n_410), .D(n_393), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_431), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_438), .B(n_383), .Y(n_463) );
NAND2xp33_ASAP7_75t_R g464 ( .A(n_430), .B(n_11), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_450), .B(n_399), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_438), .B(n_406), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_432), .B(n_416), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_432), .B(n_406), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_439), .B(n_406), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_431), .B(n_12), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_423), .Y(n_471) );
INVx2_ASAP7_75t_SL g472 ( .A(n_412), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_427), .B(n_12), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_411), .B(n_154), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_429), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_425), .B(n_13), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_425), .B(n_13), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_425), .B(n_14), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_440), .B(n_15), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_451), .B(n_15), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_440), .B(n_18), .Y(n_481) );
NAND4xp25_ASAP7_75t_L g482 ( .A(n_443), .B(n_20), .C(n_305), .D(n_253), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_417), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_434), .A2(n_327), .B1(n_282), .B2(n_235), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_420), .B(n_327), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_417), .B(n_20), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_425), .Y(n_487) );
NOR2xp33_ASAP7_75t_R g488 ( .A(n_420), .B(n_327), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_430), .A2(n_282), .B(n_280), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_419), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_453), .B(n_282), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_430), .B(n_22), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_453), .Y(n_493) );
AND2x4_ASAP7_75t_L g494 ( .A(n_436), .B(n_25), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_422), .Y(n_495) );
OAI33xp33_ASAP7_75t_L g496 ( .A1(n_441), .A2(n_26), .A3(n_28), .B1(n_30), .B2(n_32), .B3(n_33), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_422), .Y(n_497) );
NAND5xp2_ASAP7_75t_SL g498 ( .A(n_444), .B(n_35), .C(n_37), .D(n_38), .E(n_39), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_424), .B(n_235), .Y(n_499) );
OAI31xp33_ASAP7_75t_L g500 ( .A1(n_482), .A2(n_421), .A3(n_437), .B(n_436), .Y(n_500) );
INVxp67_ASAP7_75t_L g501 ( .A(n_462), .Y(n_501) );
OAI21xp33_ASAP7_75t_L g502 ( .A1(n_455), .A2(n_452), .B(n_441), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_471), .B(n_413), .Y(n_503) );
BUFx2_ASAP7_75t_SL g504 ( .A(n_472), .Y(n_504) );
OA22x2_ASAP7_75t_L g505 ( .A1(n_454), .A2(n_436), .B1(n_452), .B2(n_442), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_483), .Y(n_506) );
INVxp67_ASAP7_75t_L g507 ( .A(n_464), .Y(n_507) );
AOI221xp5_ASAP7_75t_L g508 ( .A1(n_460), .A2(n_447), .B1(n_435), .B2(n_442), .C(n_424), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_475), .B(n_428), .Y(n_509) );
INVx2_ASAP7_75t_SL g510 ( .A(n_488), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_490), .Y(n_511) );
NOR2xp33_ASAP7_75t_SL g512 ( .A(n_492), .B(n_436), .Y(n_512) );
OAI21xp33_ASAP7_75t_SL g513 ( .A1(n_485), .A2(n_426), .B(n_413), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_495), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_467), .B(n_426), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_456), .B(n_448), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_469), .B(n_43), .Y(n_517) );
OAI21xp33_ASAP7_75t_SL g518 ( .A1(n_461), .A2(n_445), .B(n_311), .Y(n_518) );
NAND2x1p5_ASAP7_75t_L g519 ( .A(n_492), .B(n_280), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_493), .B(n_48), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_455), .A2(n_293), .B1(n_280), .B2(n_311), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_474), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_497), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_486), .Y(n_524) );
OAI31xp33_ASAP7_75t_L g525 ( .A1(n_480), .A2(n_49), .A3(n_50), .B(n_51), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_459), .A2(n_234), .B1(n_293), .B2(n_280), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_470), .A2(n_181), .B1(n_55), .B2(n_56), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_474), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_476), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_457), .B(n_52), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_466), .B(n_57), .Y(n_531) );
AOI322xp5_ASAP7_75t_L g532 ( .A1(n_479), .A2(n_60), .A3(n_62), .B1(n_66), .B2(n_67), .C1(n_68), .C2(n_69), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_465), .B(n_70), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_457), .B(n_71), .Y(n_534) );
INVxp67_ASAP7_75t_SL g535 ( .A(n_463), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_479), .B(n_74), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_458), .B(n_174), .Y(n_537) );
AOI222xp33_ASAP7_75t_L g538 ( .A1(n_481), .A2(n_174), .B1(n_182), .B2(n_192), .C1(n_204), .C2(n_181), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_477), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_487), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_478), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_494), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_466), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_468), .A2(n_174), .B1(n_182), .B2(n_192), .Y(n_544) );
AOI322xp5_ASAP7_75t_L g545 ( .A1(n_463), .A2(n_174), .A3(n_181), .B1(n_182), .B2(n_192), .C1(n_204), .C2(n_484), .Y(n_545) );
OAI221xp5_ASAP7_75t_L g546 ( .A1(n_507), .A2(n_473), .B1(n_468), .B2(n_491), .C(n_489), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_501), .B(n_499), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_535), .B(n_499), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_506), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_504), .Y(n_550) );
INVx4_ASAP7_75t_L g551 ( .A(n_519), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_543), .B(n_174), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_511), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_510), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_514), .Y(n_555) );
INVx1_ASAP7_75t_SL g556 ( .A(n_542), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_524), .B(n_496), .Y(n_557) );
XOR2x2_ASAP7_75t_L g558 ( .A(n_505), .B(n_498), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_523), .Y(n_559) );
NAND2xp33_ASAP7_75t_L g560 ( .A(n_519), .B(n_192), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_540), .Y(n_561) );
NAND4xp25_ASAP7_75t_SL g562 ( .A(n_513), .B(n_181), .C(n_204), .D(n_500), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_515), .Y(n_563) );
INVx2_ASAP7_75t_SL g564 ( .A(n_505), .Y(n_564) );
AND2x2_ASAP7_75t_SL g565 ( .A(n_512), .B(n_508), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_503), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_509), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_529), .B(n_539), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_522), .B(n_541), .Y(n_569) );
A2O1A1Ixp33_ASAP7_75t_SL g570 ( .A1(n_525), .A2(n_520), .B(n_527), .C(n_536), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_522), .B(n_528), .Y(n_571) );
O2A1O1Ixp5_ASAP7_75t_L g572 ( .A1(n_527), .A2(n_521), .B(n_517), .C(n_534), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_537), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_502), .B(n_516), .Y(n_574) );
NOR3xp33_ASAP7_75t_SL g575 ( .A(n_518), .B(n_521), .C(n_534), .Y(n_575) );
AOI21x1_ASAP7_75t_L g576 ( .A1(n_558), .A2(n_530), .B(n_533), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_549), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_564), .A2(n_531), .B1(n_526), .B2(n_544), .Y(n_578) );
AO221x1_ASAP7_75t_L g579 ( .A1(n_554), .A2(n_532), .B1(n_538), .B2(n_545), .C(n_564), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_569), .B(n_538), .Y(n_580) );
XNOR2x1_ASAP7_75t_L g581 ( .A(n_550), .B(n_558), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_565), .A2(n_575), .B1(n_562), .B2(n_546), .Y(n_582) );
INVx1_ASAP7_75t_SL g583 ( .A(n_556), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_551), .B(n_572), .Y(n_584) );
BUFx3_ASAP7_75t_L g585 ( .A(n_551), .Y(n_585) );
INVxp67_ASAP7_75t_L g586 ( .A(n_568), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_563), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_553), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_561), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_566), .B(n_567), .Y(n_590) );
AOI222xp33_ASAP7_75t_L g591 ( .A1(n_579), .A2(n_574), .B1(n_557), .B2(n_548), .C1(n_547), .C2(n_559), .Y(n_591) );
OAI322xp33_ASAP7_75t_SL g592 ( .A1(n_584), .A2(n_555), .A3(n_573), .B1(n_561), .B2(n_570), .C1(n_571), .C2(n_560), .Y(n_592) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_580), .B(n_552), .C(n_578), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_587), .B(n_590), .Y(n_594) );
INVx5_ASAP7_75t_L g595 ( .A(n_585), .Y(n_595) );
NOR3xp33_ASAP7_75t_L g596 ( .A(n_576), .B(n_585), .C(n_588), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_577), .A2(n_579), .B1(n_565), .B2(n_582), .Y(n_597) );
NOR3x2_ASAP7_75t_L g598 ( .A(n_589), .B(n_581), .C(n_579), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_579), .A2(n_584), .B1(n_587), .B2(n_586), .C(n_590), .Y(n_599) );
AO22x2_ASAP7_75t_L g600 ( .A1(n_581), .A2(n_584), .B1(n_564), .B2(n_583), .Y(n_600) );
AOI211xp5_ASAP7_75t_SL g601 ( .A1(n_582), .A2(n_507), .B(n_578), .C(n_560), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_595), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_599), .A2(n_597), .B1(n_601), .B2(n_591), .C(n_596), .Y(n_603) );
NOR2x1p5_ASAP7_75t_L g604 ( .A(n_593), .B(n_594), .Y(n_604) );
XNOR2xp5_ASAP7_75t_L g605 ( .A(n_603), .B(n_598), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_602), .B(n_595), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_605), .Y(n_607) );
INVx2_ASAP7_75t_SL g608 ( .A(n_607), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_608), .A2(n_600), .B1(n_606), .B2(n_604), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_609), .A2(n_600), .B(n_592), .Y(n_610) );
endmodule