module fake_jpeg_19006_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_6),
.B(n_1),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx11_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_24),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_18),
.B(n_17),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_17),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_23),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_24),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_20),
.A2(n_13),
.B1(n_15),
.B2(n_12),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_10),
.B1(n_9),
.B2(n_13),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_21),
.B1(n_12),
.B2(n_22),
.Y(n_35)
);

OAI32xp33_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_26),
.A3(n_14),
.B1(n_9),
.B2(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_24),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_22),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_32),
.B(n_33),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_43),
.B(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_22),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_37),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_8),
.B(n_3),
.Y(n_53)
);

NOR3xp33_ASAP7_75t_SL g48 ( 
.A(n_46),
.B(n_41),
.C(n_14),
.Y(n_48)
);

AOI322xp5_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_50),
.A3(n_7),
.B1(n_8),
.B2(n_17),
.C1(n_10),
.C2(n_4),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_52),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_3),
.B(n_4),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_50),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_21),
.B1(n_4),
.B2(n_5),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_58),
.A2(n_57),
.B1(n_55),
.B2(n_21),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_0),
.B(n_58),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_0),
.Y(n_61)
);


endmodule