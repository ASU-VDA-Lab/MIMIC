module fake_jpeg_14443_n_645 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_645);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_645;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_538;
wire n_47;
wire n_625;
wire n_312;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_14),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVxp33_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_27),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_62),
.B(n_63),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_19),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_27),
.B(n_14),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_67),
.B(n_72),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_68),
.Y(n_177)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g191 ( 
.A(n_69),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_71),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_31),
.B(n_13),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_73),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_13),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_74),
.B(n_81),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_75),
.Y(n_174)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_77),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

BUFx24_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g132 ( 
.A(n_79),
.Y(n_132)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_46),
.B(n_1),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_83),
.Y(n_178)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_85),
.B(n_88),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_86),
.Y(n_193)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_87),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_21),
.B(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_89),
.B(n_91),
.Y(n_212)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_90),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_19),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_19),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_92),
.B(n_95),
.Y(n_214)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_93),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_94),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_45),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_96),
.Y(n_195)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_21),
.B(n_54),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_99),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_25),
.B(n_3),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_101),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_45),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_102),
.B(n_103),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_45),
.Y(n_103)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_104),
.Y(n_197)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g203 ( 
.A(n_105),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_106),
.Y(n_196)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_38),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_108),
.Y(n_209)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g208 ( 
.A(n_109),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_44),
.B(n_3),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_110),
.B(n_120),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_111),
.Y(n_216)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_38),
.Y(n_112)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_112),
.Y(n_207)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_29),
.B(n_3),
.Y(n_114)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_23),
.Y(n_115)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_28),
.Y(n_117)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_45),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_118),
.Y(n_210)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_29),
.Y(n_119)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_41),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_37),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_37),
.Y(n_122)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_30),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_37),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_22),
.Y(n_126)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_126),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_32),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_127),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_32),
.Y(n_128)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_42),
.Y(n_129)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_42),
.Y(n_130)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_70),
.A2(n_49),
.B1(n_28),
.B2(n_48),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_138),
.A2(n_52),
.B1(n_104),
.B2(n_39),
.Y(n_240)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_149),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_68),
.A2(n_32),
.B1(n_47),
.B2(n_55),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_151),
.A2(n_117),
.B1(n_128),
.B2(n_127),
.Y(n_235)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_153),
.Y(n_238)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_65),
.Y(n_156)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_156),
.Y(n_262)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

INVx11_ASAP7_75t_L g246 ( 
.A(n_158),
.Y(n_246)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_160),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_79),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_163),
.B(n_190),
.Y(n_218)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_88),
.B(n_61),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_164),
.B(n_9),
.Y(n_291)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_165),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_61),
.C(n_58),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_168),
.B(n_24),
.C(n_22),
.Y(n_245)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_170),
.Y(n_237)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_173),
.Y(n_266)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_94),
.Y(n_175)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_175),
.Y(n_268)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_180),
.Y(n_282)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_109),
.Y(n_181)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_181),
.Y(n_283)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_64),
.Y(n_182)
);

INVx5_ASAP7_75t_SL g251 ( 
.A(n_182),
.Y(n_251)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_115),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_183),
.Y(n_242)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_76),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_93),
.B(n_58),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_192),
.B(n_50),
.Y(n_258)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_83),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_198),
.Y(n_232)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_87),
.Y(n_202)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

INVx11_ASAP7_75t_L g204 ( 
.A(n_80),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_204),
.Y(n_263)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_121),
.Y(n_215)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g219 ( 
.A(n_143),
.B(n_66),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_219),
.B(n_245),
.Y(n_296)
);

AO22x2_ASAP7_75t_L g222 ( 
.A1(n_132),
.A2(n_101),
.B1(n_77),
.B2(n_75),
.Y(n_222)
);

AO22x1_ASAP7_75t_SL g300 ( 
.A1(n_222),
.A2(n_131),
.B1(n_139),
.B2(n_211),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_186),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_223),
.B(n_227),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_141),
.Y(n_224)
);

INVx5_ASAP7_75t_L g342 ( 
.A(n_224),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_122),
.B1(n_86),
.B2(n_73),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_225),
.A2(n_240),
.B1(n_252),
.B2(n_275),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_141),
.Y(n_226)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_226),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_150),
.B(n_50),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_169),
.Y(n_228)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_228),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_157),
.B(n_148),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_230),
.B(n_233),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_167),
.B(n_111),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_167),
.B(n_71),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_234),
.B(n_236),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_235),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_214),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_157),
.B(n_34),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_241),
.B(n_247),
.Y(n_332)
);

CKINVDCx12_ASAP7_75t_R g243 ( 
.A(n_191),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_243),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_206),
.A2(n_34),
.B1(n_57),
.B2(n_56),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_244),
.A2(n_292),
.B1(n_133),
.B2(n_189),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_214),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_164),
.B(n_55),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_248),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_138),
.A2(n_39),
.B1(n_57),
.B2(n_56),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_166),
.Y(n_253)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_253),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_203),
.A2(n_55),
.B1(n_47),
.B2(n_24),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_254),
.A2(n_277),
.B1(n_132),
.B2(n_144),
.Y(n_297)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_166),
.Y(n_255)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_255),
.Y(n_309)
);

BUFx2_ASAP7_75t_SL g256 ( 
.A(n_201),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_256),
.Y(n_299)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_205),
.Y(n_257)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_257),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_258),
.B(n_259),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_187),
.B(n_53),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_210),
.B(n_53),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_260),
.B(n_261),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_146),
.B(n_40),
.Y(n_261)
);

BUFx2_ASAP7_75t_SL g264 ( 
.A(n_209),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_264),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_169),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_265),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_174),
.Y(n_267)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_267),
.Y(n_340)
);

AND2x2_ASAP7_75t_SL g269 ( 
.A(n_164),
.B(n_55),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_291),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_197),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_270),
.B(n_272),
.Y(n_345)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_205),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_271),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_187),
.B(n_212),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_212),
.B(n_40),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_273),
.B(n_274),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_188),
.B(n_125),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_172),
.A2(n_69),
.B1(n_4),
.B2(n_5),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_174),
.Y(n_276)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_203),
.A2(n_69),
.B1(n_4),
.B2(n_5),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_206),
.B(n_3),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_278),
.B(n_279),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_146),
.B(n_6),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_136),
.B(n_6),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_280),
.B(n_288),
.Y(n_351)
);

AO22x1_ASAP7_75t_L g281 ( 
.A1(n_197),
.A2(n_147),
.B1(n_161),
.B2(n_145),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_281),
.A2(n_135),
.B(n_159),
.Y(n_335)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_155),
.Y(n_284)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_142),
.Y(n_285)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_285),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_134),
.A2(n_199),
.B1(n_208),
.B2(n_193),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_286),
.A2(n_200),
.B1(n_196),
.B2(n_162),
.Y(n_311)
);

O2A1O1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_209),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_287)
);

O2A1O1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_287),
.A2(n_144),
.B(n_176),
.C(n_177),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_172),
.B(n_8),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_140),
.B(n_9),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_289),
.B(n_290),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_171),
.B(n_9),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_151),
.A2(n_10),
.B1(n_11),
.B2(n_208),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_152),
.B(n_10),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_293),
.A2(n_211),
.B1(n_195),
.B2(n_217),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_297),
.Y(n_366)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_298),
.Y(n_357)
);

OAI21xp33_ASAP7_75t_SL g359 ( 
.A1(n_300),
.A2(n_320),
.B(n_222),
.Y(n_359)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_301),
.Y(n_363)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_302),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_232),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_303),
.B(n_306),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_218),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_184),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_308),
.B(n_336),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_311),
.A2(n_246),
.B1(n_265),
.B2(n_224),
.Y(n_367)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_268),
.Y(n_313)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_313),
.Y(n_394)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_316),
.Y(n_396)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_282),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_317),
.Y(n_365)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_239),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_321),
.B(n_324),
.Y(n_381)
);

NAND2x1_ASAP7_75t_SL g322 ( 
.A(n_281),
.B(n_269),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_322),
.A2(n_335),
.B(n_346),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_251),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_323),
.B(n_285),
.Y(n_385)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_239),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_249),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_326),
.B(n_329),
.Y(n_393)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_249),
.Y(n_328)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_328),
.Y(n_373)
);

OAI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_240),
.A2(n_200),
.B1(n_179),
.B2(n_178),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_333),
.A2(n_348),
.B1(n_292),
.B2(n_251),
.Y(n_360)
);

NOR2x1p5_ASAP7_75t_L g334 ( 
.A(n_222),
.B(n_137),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_334),
.B(n_222),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_248),
.B(n_207),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_291),
.B(n_154),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_291),
.C(n_219),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_343),
.A2(n_254),
.B1(n_286),
.B2(n_277),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_219),
.B(n_216),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_235),
.A2(n_176),
.B1(n_216),
.B2(n_245),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_220),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_350),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_354),
.B(n_338),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_356),
.B(n_400),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_299),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_358),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g406 ( 
.A1(n_359),
.A2(n_367),
.B1(n_399),
.B2(n_346),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_360),
.A2(n_366),
.B(n_361),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_322),
.B(n_274),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_368),
.Y(n_403)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_327),
.Y(n_362)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_362),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_346),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_364),
.B(n_369),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_296),
.B(n_221),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_325),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_370),
.Y(n_407)
);

INVx13_ASAP7_75t_L g371 ( 
.A(n_341),
.Y(n_371)
);

INVx3_ASAP7_75t_SL g414 ( 
.A(n_371),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_315),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_374),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_330),
.A2(n_263),
.B1(n_267),
.B2(n_226),
.Y(n_374)
);

INVx6_ASAP7_75t_L g376 ( 
.A(n_342),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_376),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_296),
.B(n_221),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_378),
.B(n_380),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_330),
.A2(n_276),
.B1(n_228),
.B2(n_242),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_296),
.B(n_229),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_382),
.B(n_383),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_238),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_305),
.B(n_262),
.C(n_266),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_308),
.C(n_305),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_385),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_311),
.A2(n_284),
.B1(n_246),
.B2(n_253),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_386),
.A2(n_397),
.B1(n_353),
.B2(n_337),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_332),
.B(n_266),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_387),
.B(n_391),
.Y(n_402)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_327),
.Y(n_388)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_388),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_331),
.B(n_250),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_389),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_345),
.B(n_250),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_310),
.B(n_242),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_392),
.B(n_398),
.Y(n_405)
);

INVx8_ASAP7_75t_L g395 ( 
.A(n_342),
.Y(n_395)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_395),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_353),
.A2(n_255),
.B1(n_257),
.B2(n_271),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_339),
.B(n_220),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_343),
.A2(n_334),
.B1(n_344),
.B2(n_335),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_305),
.A2(n_287),
.B(n_237),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_360),
.A2(n_334),
.B1(n_300),
.B2(n_344),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_404),
.A2(n_416),
.B1(n_429),
.B2(n_436),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_406),
.A2(n_377),
.B(n_384),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_408),
.A2(n_421),
.B(n_432),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_409),
.B(n_415),
.C(n_420),
.Y(n_442)
);

OA22x2_ASAP7_75t_L g411 ( 
.A1(n_356),
.A2(n_300),
.B1(n_320),
.B2(n_314),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_411),
.B(n_380),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_382),
.A2(n_351),
.B1(n_349),
.B2(n_308),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_368),
.B(n_336),
.C(n_307),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_355),
.A2(n_336),
.B(n_347),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_372),
.B(n_317),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_422),
.Y(n_475)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_357),
.Y(n_424)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_424),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_378),
.B(n_304),
.C(n_328),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_425),
.B(n_426),
.C(n_390),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_354),
.B(n_231),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_381),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_427),
.B(n_430),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_428),
.B(n_373),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_366),
.A2(n_295),
.B1(n_340),
.B2(n_318),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_375),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_355),
.A2(n_337),
.B(n_237),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_392),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_433),
.B(n_439),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_369),
.A2(n_295),
.B1(n_340),
.B2(n_319),
.Y(n_436)
);

HAxp5_ASAP7_75t_SL g438 ( 
.A(n_364),
.B(n_294),
.CON(n_438),
.SN(n_438)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_438),
.B(n_400),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_383),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_407),
.A2(n_393),
.B1(n_399),
.B2(n_370),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_440),
.A2(n_462),
.B1(n_470),
.B2(n_421),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_422),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_443),
.B(n_444),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_402),
.Y(n_444)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_446),
.B(n_450),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_433),
.B(n_387),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_448),
.B(n_449),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_398),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_402),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_451),
.B(n_468),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_419),
.A2(n_377),
.B(n_358),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_452),
.B(n_455),
.Y(n_504)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_424),
.Y(n_454)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_454),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_412),
.B(n_377),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_456),
.B(n_459),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_457),
.A2(n_471),
.B(n_411),
.Y(n_507)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_423),
.Y(n_458)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_458),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_426),
.B(n_363),
.C(n_357),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_439),
.B(n_394),
.Y(n_460)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_460),
.Y(n_488)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_436),
.Y(n_461)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_461),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_407),
.A2(n_374),
.B1(n_390),
.B2(n_394),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_410),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_463),
.B(n_444),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_415),
.B(n_363),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_464),
.B(n_420),
.Y(n_494)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_410),
.Y(n_465)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_465),
.Y(n_503)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_413),
.Y(n_466)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_466),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_404),
.A2(n_395),
.B1(n_376),
.B2(n_388),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_467),
.A2(n_469),
.B1(n_414),
.B2(n_417),
.Y(n_501)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_413),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_434),
.A2(n_362),
.B1(n_396),
.B2(n_379),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_419),
.A2(n_318),
.B1(n_319),
.B2(n_396),
.Y(n_470)
);

INVx13_ASAP7_75t_L g472 ( 
.A(n_414),
.Y(n_472)
);

BUFx4f_ASAP7_75t_SL g505 ( 
.A(n_472),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_405),
.B(n_379),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_473),
.B(n_401),
.Y(n_498)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_478),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_471),
.A2(n_452),
.B(n_447),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_479),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_460),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_480),
.B(n_507),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_427),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_481),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_464),
.B(n_409),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_483),
.B(n_494),
.Y(n_514)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_458),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_486),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_405),
.Y(n_487)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_487),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_445),
.B(n_434),
.Y(n_490)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_490),
.Y(n_533)
);

NOR3xp33_ASAP7_75t_SL g491 ( 
.A(n_448),
.B(n_437),
.C(n_403),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_491),
.B(n_492),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_474),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_469),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_493),
.B(n_500),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_463),
.B(n_465),
.Y(n_495)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_495),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_457),
.A2(n_419),
.B1(n_403),
.B2(n_411),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_496),
.A2(n_462),
.B1(n_446),
.B2(n_411),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_497),
.A2(n_441),
.B1(n_443),
.B2(n_447),
.Y(n_510)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_498),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_455),
.B(n_418),
.Y(n_500)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_501),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_442),
.B(n_437),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_502),
.B(n_453),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_459),
.B(n_416),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_509),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_510),
.A2(n_513),
.B1(n_517),
.B2(n_488),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_480),
.B(n_495),
.Y(n_512)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_512),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_485),
.A2(n_441),
.B1(n_467),
.B2(n_461),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_497),
.A2(n_473),
.B1(n_440),
.B2(n_450),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_442),
.C(n_456),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_519),
.B(n_523),
.C(n_529),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_477),
.B(n_475),
.Y(n_520)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_520),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_425),
.C(n_471),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_477),
.B(n_470),
.Y(n_525)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_525),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_482),
.B(n_468),
.Y(n_526)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_526),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_482),
.B(n_466),
.Y(n_527)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_527),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_502),
.B(n_432),
.C(n_428),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_531),
.A2(n_504),
.B1(n_538),
.B2(n_539),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_494),
.B(n_454),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_532),
.B(n_535),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_534),
.B(n_539),
.C(n_499),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_483),
.B(n_453),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_489),
.B(n_417),
.C(n_411),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_511),
.B(n_479),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_540),
.A2(n_525),
.B(n_512),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_514),
.B(n_489),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_541),
.B(n_549),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_SL g542 ( 
.A(n_535),
.B(n_496),
.Y(n_542)
);

MAJx2_ASAP7_75t_L g573 ( 
.A(n_542),
.B(n_550),
.C(n_555),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_544),
.A2(n_429),
.B1(n_414),
.B2(n_431),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_546),
.A2(n_554),
.B1(n_531),
.B2(n_560),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_519),
.B(n_490),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_547),
.B(n_563),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_514),
.B(n_504),
.Y(n_549)
);

XNOR2x1_ASAP7_75t_SL g550 ( 
.A(n_529),
.B(n_491),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_516),
.B(n_484),
.Y(n_551)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_551),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_522),
.B(n_484),
.Y(n_552)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_552),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_517),
.A2(n_488),
.B1(n_485),
.B2(n_499),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_521),
.B(n_500),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_556),
.B(n_557),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_523),
.B(n_503),
.C(n_507),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_537),
.A2(n_503),
.B1(n_498),
.B2(n_476),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_558),
.A2(n_536),
.B1(n_524),
.B2(n_518),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_515),
.B(n_486),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_561),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_SL g562 ( 
.A(n_534),
.B(n_508),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_562),
.B(n_533),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_532),
.B(n_508),
.C(n_476),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_553),
.B(n_537),
.Y(n_565)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_565),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_548),
.B(n_528),
.C(n_538),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_566),
.B(n_577),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_540),
.Y(n_567)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_567),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_570),
.A2(n_579),
.B1(n_505),
.B2(n_472),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_563),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_571),
.B(n_555),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_572),
.B(n_542),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_545),
.B(n_520),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_574),
.Y(n_595)
);

NAND2xp33_ASAP7_75t_SL g575 ( 
.A(n_559),
.B(n_511),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_575),
.A2(n_576),
.B(n_578),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_548),
.B(n_530),
.C(n_526),
.Y(n_577)
);

AOI21x1_ASAP7_75t_L g578 ( 
.A1(n_564),
.A2(n_527),
.B(n_530),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_554),
.A2(n_557),
.B(n_540),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_580),
.A2(n_541),
.B(n_550),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_582),
.A2(n_567),
.B1(n_580),
.B2(n_565),
.Y(n_588)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_586),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_588),
.B(n_574),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_583),
.B(n_549),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g610 ( 
.A(n_590),
.B(n_602),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_591),
.B(n_601),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_592),
.B(n_596),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_585),
.B(n_562),
.Y(n_593)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_593),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_566),
.B(n_577),
.C(n_568),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_594),
.B(n_596),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_569),
.B(n_543),
.C(n_435),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_584),
.A2(n_505),
.B1(n_431),
.B2(n_435),
.Y(n_599)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_599),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_569),
.B(n_373),
.C(n_365),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_600),
.B(n_603),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_581),
.B(n_365),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_573),
.B(n_570),
.Y(n_603)
);

CKINVDCx14_ASAP7_75t_R g607 ( 
.A(n_593),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_607),
.B(n_613),
.Y(n_619)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_608),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_612),
.B(n_600),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_587),
.B(n_573),
.C(n_576),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_594),
.B(n_575),
.C(n_578),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_615),
.B(n_617),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_SL g616 ( 
.A1(n_591),
.A2(n_582),
.B(n_505),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_616),
.A2(n_589),
.B(n_601),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_586),
.B(n_365),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_SL g618 ( 
.A1(n_608),
.A2(n_597),
.B1(n_605),
.B2(n_611),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_618),
.B(n_621),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_604),
.B(n_595),
.Y(n_620)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_620),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_610),
.B(n_614),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_612),
.B(n_603),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_622),
.B(n_624),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_626),
.B(n_627),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_613),
.B(n_588),
.Y(n_627)
);

AOI322xp5_ASAP7_75t_L g628 ( 
.A1(n_623),
.A2(n_606),
.A3(n_615),
.B1(n_598),
.B2(n_589),
.C1(n_609),
.C2(n_472),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_628),
.B(n_625),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_619),
.A2(n_609),
.B(n_592),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_SL g637 ( 
.A(n_629),
.B(n_632),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_627),
.A2(n_294),
.B(n_309),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_635),
.A2(n_636),
.B(n_638),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_630),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_SL g638 ( 
.A(n_634),
.B(n_624),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_637),
.B(n_631),
.C(n_633),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_640),
.B(n_630),
.C(n_309),
.Y(n_641)
);

MAJx2_ASAP7_75t_L g642 ( 
.A(n_641),
.B(n_639),
.C(n_371),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_642),
.B(n_312),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_643),
.B(n_302),
.C(n_316),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_644),
.B(n_312),
.C(n_231),
.Y(n_645)
);


endmodule