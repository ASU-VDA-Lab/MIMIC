module fake_jpeg_3686_n_487 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_487);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_487;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_SL g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_8),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_48),
.B(n_39),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_51),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_17),
.B(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_63),
.Y(n_101)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_8),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_54),
.B(n_67),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_55),
.Y(n_141)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_29),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_18),
.B(n_14),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_25),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_88),
.Y(n_117)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_25),
.B(n_7),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_90),
.Y(n_151)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_94),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_21),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_25),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_21),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_38),
.B1(n_40),
.B2(n_34),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_98),
.A2(n_111),
.B1(n_127),
.B2(n_129),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_38),
.B1(n_32),
.B2(n_40),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_131),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_69),
.A2(n_22),
.B1(n_26),
.B2(n_34),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_128),
.B(n_137),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_43),
.A2(n_26),
.B1(n_22),
.B2(n_32),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_58),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_48),
.B(n_35),
.Y(n_137)
);

INVx6_ASAP7_75t_SL g139 ( 
.A(n_90),
.Y(n_139)
);

CKINVDCx12_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_72),
.B(n_39),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_143),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_74),
.B(n_35),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_79),
.B(n_31),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_86),
.Y(n_176)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_155),
.Y(n_213)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_156),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_89),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_157),
.Y(n_207)
);

BUFx12_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_L g159 ( 
.A1(n_98),
.A2(n_84),
.B1(n_76),
.B2(n_75),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_166),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_105),
.A2(n_31),
.B1(n_23),
.B2(n_18),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_108),
.A2(n_46),
.B1(n_50),
.B2(n_55),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_162),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_101),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_174),
.Y(n_202)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_110),
.A2(n_45),
.B1(n_66),
.B2(n_61),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_99),
.Y(n_167)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_71),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_169),
.B(n_190),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_125),
.A2(n_60),
.B1(n_68),
.B2(n_82),
.Y(n_173)
);

OAI22x1_ASAP7_75t_L g215 ( 
.A1(n_173),
.A2(n_153),
.B1(n_130),
.B2(n_144),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_116),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_178),
.Y(n_218)
);

NOR4xp25_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_11),
.C(n_14),
.D(n_2),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g214 ( 
.A(n_177),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_100),
.B(n_97),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_182),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_112),
.B(n_59),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_192),
.Y(n_227)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_107),
.Y(n_185)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_103),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_103),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_129),
.B(n_0),
.Y(n_190)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_109),
.Y(n_191)
);

INVx5_ASAP7_75t_SL g222 ( 
.A(n_191),
.Y(n_222)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_197),
.Y(n_212)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_102),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_133),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_118),
.B(n_0),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_145),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_121),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_198),
.A2(n_141),
.B1(n_120),
.B2(n_132),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_204),
.B(n_162),
.Y(n_240)
);

NAND2x1p5_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_96),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_208),
.B(n_190),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g209 ( 
.A(n_157),
.B(n_138),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_217),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

OAI32xp33_ASAP7_75t_L g216 ( 
.A1(n_169),
.A2(n_148),
.A3(n_142),
.B1(n_152),
.B2(n_127),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_180),
.A2(n_146),
.B(n_153),
.Y(n_217)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_225),
.Y(n_232)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_233),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_236),
.Y(n_262)
);

INVx13_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_235),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_226),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_211),
.A2(n_173),
.B1(n_196),
.B2(n_171),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_237),
.A2(n_239),
.B1(n_244),
.B2(n_254),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_217),
.A2(n_181),
.B1(n_159),
.B2(n_175),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_242),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_172),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_211),
.A2(n_144),
.B1(n_106),
.B2(n_130),
.Y(n_244)
);

INVx13_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_245),
.Y(n_260)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_179),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_208),
.C(n_209),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_192),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_250),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_185),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_202),
.B(n_194),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_253),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_214),
.B(n_195),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_207),
.A2(n_147),
.B1(n_106),
.B2(n_141),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_227),
.B(n_198),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_257),
.Y(n_272)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_216),
.A2(n_147),
.B1(n_133),
.B2(n_132),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_221),
.Y(n_258)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_261),
.B(n_234),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_209),
.C(n_200),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_282),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_200),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_269),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_249),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_208),
.Y(n_273)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_241),
.A2(n_231),
.B1(n_215),
.B2(n_212),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_276),
.A2(n_281),
.B1(n_283),
.B2(n_238),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_251),
.A2(n_219),
.B(n_229),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_277),
.A2(n_271),
.B(n_259),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_238),
.A2(n_239),
.B1(n_244),
.B2(n_232),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_278),
.A2(n_274),
.B1(n_238),
.B2(n_272),
.Y(n_291)
);

OA21x2_ASAP7_75t_L g280 ( 
.A1(n_257),
.A2(n_219),
.B(n_229),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_280),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_251),
.A2(n_224),
.B1(n_168),
.B2(n_223),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_255),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_251),
.A2(n_224),
.B1(n_199),
.B2(n_186),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_277),
.A2(n_251),
.B(n_250),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_287),
.A2(n_290),
.B(n_310),
.Y(n_317)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_266),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_299),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_291),
.A2(n_297),
.B1(n_301),
.B2(n_303),
.Y(n_330)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_265),
.Y(n_318)
);

AND2x6_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_234),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_294),
.B(n_280),
.Y(n_338)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_295),
.Y(n_326)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_279),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_296),
.Y(n_332)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_270),
.B(n_242),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_305),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_274),
.A2(n_232),
.B1(n_252),
.B2(n_243),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_274),
.A2(n_246),
.B1(n_236),
.B2(n_256),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_306),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_270),
.B(n_220),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_272),
.A2(n_254),
.B1(n_256),
.B2(n_258),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_307),
.A2(n_278),
.B1(n_269),
.B2(n_266),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_263),
.B(n_264),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_247),
.Y(n_331)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_281),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_280),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_273),
.A2(n_170),
.B(n_191),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_SL g311 ( 
.A(n_265),
.B(n_245),
.C(n_233),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_311),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_289),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_312),
.B(n_315),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_314),
.A2(n_291),
.B1(n_309),
.B2(n_297),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_286),
.B(n_263),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_318),
.B(n_310),
.Y(n_340)
);

A2O1A1O1Ixp25_ASAP7_75t_L g319 ( 
.A1(n_286),
.A2(n_262),
.B(n_261),
.C(n_264),
.D(n_267),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_319),
.A2(n_323),
.B(n_235),
.Y(n_354)
);

AO22x1_ASAP7_75t_L g320 ( 
.A1(n_285),
.A2(n_276),
.B1(n_283),
.B2(n_280),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_320),
.B(n_321),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_285),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_290),
.B(n_267),
.Y(n_322)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_322),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_287),
.A2(n_262),
.B(n_280),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_303),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_329),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_288),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_331),
.A2(n_337),
.B1(n_268),
.B2(n_210),
.Y(n_350)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_333),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_302),
.B(n_261),
.Y(n_335)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_335),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_220),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_336),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_302),
.B(n_260),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_338),
.B(n_213),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_260),
.Y(n_339)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_339),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_340),
.B(n_353),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_341),
.A2(n_360),
.B1(n_329),
.B2(n_332),
.Y(n_380)
);

AND2x2_ASAP7_75t_SL g342 ( 
.A(n_322),
.B(n_311),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_342),
.B(n_317),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_304),
.C(n_299),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_343),
.B(n_351),
.C(n_364),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_335),
.B(n_294),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_346),
.B(n_165),
.Y(n_390)
);

AO22x1_ASAP7_75t_L g347 ( 
.A1(n_333),
.A2(n_292),
.B1(n_296),
.B2(n_295),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_347),
.A2(n_358),
.B(n_312),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_330),
.A2(n_307),
.B1(n_305),
.B2(n_275),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_349),
.A2(n_356),
.B1(n_320),
.B2(n_314),
.Y(n_374)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_350),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_268),
.C(n_210),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_337),
.B(n_203),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_354),
.B(n_315),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_330),
.A2(n_201),
.B1(n_205),
.B2(n_233),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_317),
.A2(n_235),
.B(n_245),
.Y(n_358)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_316),
.Y(n_361)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_361),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_338),
.A2(n_201),
.B1(n_205),
.B2(n_253),
.Y(n_363)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_363),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_323),
.B(n_203),
.C(n_193),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_328),
.B(n_213),
.Y(n_365)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_365),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_366),
.Y(n_398)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_368),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_343),
.B(n_339),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_371),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_346),
.B(n_327),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_374),
.A2(n_379),
.B1(n_382),
.B2(n_341),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_327),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_375),
.B(n_351),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_358),
.A2(n_319),
.B(n_316),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_377),
.B(n_381),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_378),
.B(n_385),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_345),
.A2(n_320),
.B1(n_325),
.B2(n_321),
.Y(n_379)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_380),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_359),
.A2(n_332),
.B1(n_326),
.B2(n_324),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_345),
.A2(n_326),
.B1(n_324),
.B2(n_313),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_352),
.B(n_313),
.C(n_206),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_384),
.B(n_353),
.C(n_364),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_340),
.B(n_352),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_348),
.Y(n_386)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_386),
.Y(n_395)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_348),
.Y(n_387)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_387),
.Y(n_404)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_388),
.Y(n_406)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_389),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_SL g394 ( 
.A(n_390),
.B(n_342),
.C(n_344),
.Y(n_394)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_391),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_383),
.B(n_344),
.C(n_342),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_393),
.B(n_184),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_394),
.B(n_376),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_369),
.B(n_355),
.Y(n_397)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_397),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_368),
.A2(n_362),
.B(n_357),
.Y(n_399)
);

MAJx2_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_375),
.C(n_390),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_379),
.A2(n_362),
.B(n_357),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_400),
.A2(n_408),
.B(n_119),
.Y(n_424)
);

INVxp33_ASAP7_75t_L g427 ( 
.A(n_403),
.Y(n_427)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_405),
.Y(n_421)
);

BUFx12_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_407),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_347),
.Y(n_408)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_384),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_155),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_373),
.B(n_349),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_356),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_402),
.A2(n_372),
.B1(n_367),
.B2(n_374),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_414),
.B(n_417),
.Y(n_440)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_415),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_383),
.C(n_385),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_SL g443 ( 
.A(n_418),
.B(n_430),
.Y(n_443)
);

FAx1_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_371),
.CI(n_370),
.CON(n_419),
.SN(n_419)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_419),
.A2(n_400),
.B(n_401),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_422),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_393),
.B(n_376),
.C(n_151),
.Y(n_422)
);

AOI221xp5_ASAP7_75t_L g444 ( 
.A1(n_423),
.A2(n_428),
.B1(n_406),
.B2(n_395),
.C(n_394),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_424),
.A2(n_119),
.B1(n_138),
.B2(n_120),
.Y(n_445)
);

BUFx24_ASAP7_75t_SL g425 ( 
.A(n_398),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_425),
.B(n_396),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_188),
.C(n_167),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_426),
.B(n_397),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_410),
.B(n_164),
.C(n_114),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_435),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_421),
.Y(n_433)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_433),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_417),
.B(n_410),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_418),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_413),
.B(n_392),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_436),
.B(n_439),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_429),
.B(n_403),
.C(n_402),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_437),
.B(n_441),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_438),
.A2(n_419),
.B(n_407),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_416),
.B(n_404),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_427),
.A2(n_409),
.B1(n_408),
.B2(n_401),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_444),
.A2(n_57),
.B1(n_158),
.B2(n_3),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_445),
.B(n_430),
.Y(n_449)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_449),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_427),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_453),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_452),
.B(n_13),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_434),
.B(n_419),
.C(n_415),
.Y(n_453)
);

AOI221xp5_ASAP7_75t_L g466 ( 
.A1(n_454),
.A2(n_458),
.B1(n_9),
.B2(n_13),
.C(n_0),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_438),
.C(n_443),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_455),
.B(n_457),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_432),
.A2(n_407),
.B(n_158),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_456),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_442),
.A2(n_146),
.B(n_85),
.Y(n_457)
);

AOI322xp5_ASAP7_75t_L g460 ( 
.A1(n_450),
.A2(n_441),
.A3(n_445),
.B1(n_27),
.B2(n_5),
.C1(n_7),
.C2(n_9),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_460),
.B(n_461),
.Y(n_470)
);

AOI322xp5_ASAP7_75t_L g461 ( 
.A1(n_446),
.A2(n_27),
.A3(n_11),
.B1(n_3),
.B2(n_7),
.C1(n_9),
.C2(n_14),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_3),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_465),
.Y(n_472)
);

AOI322xp5_ASAP7_75t_L g465 ( 
.A1(n_447),
.A2(n_27),
.A3(n_3),
.B1(n_9),
.B2(n_12),
.C1(n_13),
.C2(n_1),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_466),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_467),
.B(n_0),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_462),
.Y(n_471)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_471),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_473),
.B(n_474),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_468),
.B(n_455),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_459),
.A2(n_453),
.B(n_456),
.Y(n_475)
);

AOI21x1_ASAP7_75t_L g480 ( 
.A1(n_475),
.A2(n_0),
.B(n_1),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_470),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_477),
.B(n_479),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_472),
.A2(n_463),
.B(n_459),
.Y(n_479)
);

NAND3xp33_ASAP7_75t_L g483 ( 
.A(n_480),
.B(n_1),
.C(n_27),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_478),
.B(n_469),
.Y(n_482)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_482),
.A2(n_483),
.B(n_476),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_484),
.A2(n_481),
.B(n_1),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_485),
.B(n_1),
.Y(n_486)
);

BUFx24_ASAP7_75t_SL g487 ( 
.A(n_486),
.Y(n_487)
);


endmodule