module real_jpeg_15201_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_457),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_0),
.B(n_458),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_1),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_82)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_1),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_1),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_167)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_1),
.A2(n_37),
.A3(n_184),
.B1(n_185),
.B2(n_188),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_1),
.A2(n_194),
.B1(n_195),
.B2(n_198),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_1),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_1),
.B(n_154),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_1),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_1),
.B(n_310),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_3),
.A2(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_3),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_3),
.A2(n_108),
.B1(n_149),
.B2(n_214),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_3),
.A2(n_108),
.B1(n_225),
.B2(n_228),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_3),
.A2(n_108),
.B1(n_238),
.B2(n_241),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_4),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_4),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_4),
.Y(n_130)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_4),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_4),
.Y(n_263)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_5),
.A2(n_143),
.B1(n_144),
.B2(n_148),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_6),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_6),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_6),
.Y(n_247)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_6),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_7),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_8),
.Y(n_125)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_8),
.Y(n_140)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_8),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_8),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_9),
.A2(n_22),
.B1(n_133),
.B2(n_136),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_9),
.A2(n_22),
.B1(n_359),
.B2(n_363),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_10),
.Y(n_79)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_10),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_10),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_12),
.Y(n_115)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_12),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_12),
.Y(n_197)
);

BUFx4f_ASAP7_75t_L g362 ( 
.A(n_12),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_13),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_13),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_174),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_173),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_155),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_19),
.B(n_155),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g459 ( 
.A(n_19),
.Y(n_459)
);

FAx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_56),
.CI(n_102),
.CON(n_19),
.SN(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_21),
.A2(n_142),
.B1(n_153),
.B2(n_154),
.Y(n_141)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_25),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_26),
.Y(n_147)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_26),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_26),
.Y(n_338)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_32),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_46),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_35),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g212 ( 
.A1(n_35),
.A2(n_46),
.B1(n_167),
.B2(n_213),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g305 ( 
.A1(n_35),
.A2(n_46),
.B1(n_167),
.B2(n_213),
.Y(n_305)
);

AO21x1_ASAP7_75t_L g404 ( 
.A1(n_35),
.A2(n_46),
.B(n_167),
.Y(n_404)
);

NAND2x1p5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_46),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_41),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_46),
.Y(n_154)
);

OA22x2_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_52),
.B2(n_54),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_51),
.Y(n_256)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_72),
.B(n_80),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_63),
.B1(n_65),
.B2(n_71),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g342 ( 
.A(n_62),
.Y(n_342)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_63),
.A2(n_64),
.B1(n_353),
.B2(n_356),
.Y(n_352)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_71),
.A2(n_190),
.B1(n_374),
.B2(n_375),
.Y(n_373)
);

OAI21x1_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_93),
.B(n_98),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_82),
.B1(n_92),
.B2(n_104),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_72),
.A2(n_82),
.B1(n_92),
.B2(n_104),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_72),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_72),
.B(n_92),
.Y(n_384)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_90),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_81),
.B(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_86),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_86),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_86),
.B(n_223),
.Y(n_222)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_93),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_100),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_109),
.C(n_141),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_103),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_103),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_103),
.B(n_212),
.C(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_103),
.A2(n_158),
.B1(n_212),
.B2(n_230),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_103),
.B(n_305),
.C(n_412),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_103),
.A2(n_158),
.B1(n_305),
.B2(n_311),
.Y(n_420)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_109),
.B(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_109),
.B(n_165),
.Y(n_444)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_132),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_111),
.Y(n_289)
);

AOI21x1_ASAP7_75t_SL g321 ( 
.A1(n_111),
.A2(n_322),
.B(n_324),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_111),
.A2(n_373),
.B(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_122),
.Y(n_121)
);

AO22x2_ASAP7_75t_L g216 ( 
.A1(n_112),
.A2(n_121),
.B1(n_217),
.B2(n_224),
.Y(n_216)
);

AO22x1_ASAP7_75t_L g234 ( 
.A1(n_112),
.A2(n_121),
.B1(n_217),
.B2(n_224),
.Y(n_234)
);

AO22x2_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_119),
.Y(n_112)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_114),
.Y(n_205)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_115),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_116),
.Y(n_357)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_118),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_120),
.Y(n_378)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_121),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_126),
.B1(n_128),
.B2(n_131),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_124),
.Y(n_229)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_125),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_132),
.A2(n_289),
.B1(n_372),
.B2(n_378),
.Y(n_371)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_140),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_153),
.B1(n_154),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_143),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_144),
.A2(n_330),
.B1(n_339),
.B2(n_343),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx2_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_161),
.C(n_163),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_L g441 ( 
.A1(n_156),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.Y(n_441)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_164),
.C(n_165),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_161),
.B(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_161),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_161),
.B(n_230),
.C(n_321),
.Y(n_426)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_162),
.B(n_404),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_162),
.B(n_444),
.Y(n_443)
);

XOR2x2_ASAP7_75t_L g440 ( 
.A(n_163),
.B(n_441),
.Y(n_440)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_171),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_171),
.B(n_340),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_438),
.B(n_454),
.Y(n_175)
);

AO221x1_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_345),
.B1(n_347),
.B2(n_431),
.C(n_437),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_315),
.B(n_344),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_298),
.B(n_314),
.Y(n_178)
);

OAI21x1_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_249),
.B(n_297),
.Y(n_179)
);

NOR2xp67_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_232),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_181),
.B(n_232),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_211),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_182),
.B(n_216),
.C(n_230),
.Y(n_313)
);

XOR2x2_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_191),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_183),
.B(n_191),
.Y(n_301)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_201),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g235 ( 
.A1(n_192),
.A2(n_236),
.B1(n_237),
.B2(n_244),
.Y(n_235)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_193),
.B(n_202),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_218),
.B(n_222),
.Y(n_217)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_197),
.Y(n_240)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_197),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_197),
.Y(n_363)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_201),
.B(n_358),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_206),
.Y(n_201)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI32xp33_ASAP7_75t_L g252 ( 
.A1(n_205),
.A2(n_222),
.A3(n_253),
.B1(n_257),
.B2(n_261),
.Y(n_252)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_207),
.Y(n_281)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_216),
.B1(n_230),
.B2(n_231),
.Y(n_211)
);

INVx3_ASAP7_75t_SL g230 ( 
.A(n_212),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_212),
.A2(n_230),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_216),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_216),
.A2(n_231),
.B1(n_252),
.B2(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_216),
.B(n_398),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_216),
.A2(n_231),
.B1(n_398),
.B2(n_424),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_217),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_217),
.B(n_323),
.Y(n_389)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.C(n_248),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_233),
.A2(n_234),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_233),
.B(n_301),
.C(n_303),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_233),
.A2(n_234),
.B1(n_351),
.B2(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_248),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_234),
.B(n_351),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_235),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_235),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_235),
.B(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_235),
.B(n_287),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_235),
.A2(n_268),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_236),
.A2(n_352),
.B1(n_358),
.B2(n_364),
.Y(n_351)
);

OA21x2_ASAP7_75t_L g282 ( 
.A1(n_237),
.A2(n_283),
.B(n_285),
.Y(n_282)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_243),
.Y(n_355)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_247),
.Y(n_284)
);

AOI21x1_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_271),
.B(n_296),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_267),
.Y(n_250)
);

NOR2xp67_ASAP7_75t_SL g296 ( 
.A(n_251),
.B(n_267),
.Y(n_296)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_252),
.Y(n_294)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_268),
.B(n_329),
.Y(n_412)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_291),
.B(n_295),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_286),
.B(n_290),
.Y(n_272)
);

NOR2x1_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_282),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_280),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_282),
.A2(n_292),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_282),
.B(n_305),
.C(n_309),
.Y(n_326)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_285),
.A2(n_352),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp33_ASAP7_75t_SL g295 ( 
.A(n_292),
.B(n_293),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_313),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_313),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_303),
.B1(n_304),
.B2(n_312),
.Y(n_299)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_301),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_311),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_305),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_305),
.A2(n_371),
.B(n_379),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_305),
.B(n_371),
.Y(n_379)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_317),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_325),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_318),
.B(n_326),
.C(n_327),
.Y(n_417)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_335),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_415),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_405),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_390),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_R g437 ( 
.A(n_348),
.B(n_390),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_369),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_349),
.B(n_370),
.C(n_450),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_350),
.B(n_393),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_351),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_368),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_380),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_379),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_379),
.A2(n_443),
.B1(n_445),
.B2(n_453),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_380),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_387),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_385),
.B2(n_386),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_382),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_382),
.A2(n_385),
.B1(n_388),
.B2(n_395),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_382),
.A2(n_386),
.B(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_383),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_385),
.B(n_388),
.Y(n_387)
);

INVxp33_ASAP7_75t_L g447 ( 
.A(n_387),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_388),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_394),
.C(n_396),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_394),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_396),
.B(n_414),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_402),
.C(n_403),
.Y(n_396)
);

XNOR2x1_ASAP7_75t_L g407 ( 
.A(n_397),
.B(n_408),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_398),
.Y(n_424)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_405),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_413),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_406),
.B(n_413),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_409),
.C(n_411),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_407),
.B(n_409),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_429),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_412),
.B(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_427),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_417),
.B(n_418),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_421),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_423),
.C(n_425),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_423),
.B1(n_425),
.B2(n_426),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_427),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_430),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_428),
.B(n_430),
.Y(n_432)
);

A2O1A1Ixp33_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_433),
.B(n_435),
.C(n_436),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_448),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_439),
.A2(n_455),
.B(n_456),
.Y(n_454)
);

NOR2xp67_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_442),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_442),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_445),
.C(n_446),
.Y(n_442)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_443),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_446),
.B(n_452),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_451),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_449),
.B(n_451),
.Y(n_455)
);


endmodule