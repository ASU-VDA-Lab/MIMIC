module real_aes_1990_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_826, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_826;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_626;
wire n_400;
wire n_539;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g226 ( .A(n_0), .B(n_148), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_1), .B(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g141 ( .A(n_2), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_3), .B(n_154), .Y(n_167) );
NAND2xp33_ASAP7_75t_SL g218 ( .A(n_4), .B(n_152), .Y(n_218) );
INVx1_ASAP7_75t_L g199 ( .A(n_5), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_6), .B(n_172), .Y(n_545) );
OAI22xp5_ASAP7_75t_SL g114 ( .A1(n_7), .A2(n_115), .B1(n_116), .B2(n_118), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_7), .Y(n_115) );
INVx1_ASAP7_75t_L g525 ( .A(n_8), .Y(n_525) );
CKINVDCx16_ASAP7_75t_R g790 ( .A(n_9), .Y(n_790) );
AND2x2_ASAP7_75t_L g165 ( .A(n_10), .B(n_158), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_11), .Y(n_492) );
INVx2_ASAP7_75t_L g159 ( .A(n_12), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_13), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g124 ( .A(n_14), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_14), .B(n_27), .Y(n_721) );
INVx1_ASAP7_75t_L g553 ( .A(n_15), .Y(n_553) );
OAI22xp5_ASAP7_75t_SL g806 ( .A1(n_16), .A2(n_27), .B1(n_775), .B2(n_807), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_16), .Y(n_807) );
AOI221x1_ASAP7_75t_L g212 ( .A1(n_17), .A2(n_136), .B1(n_213), .B2(n_215), .C(n_217), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_18), .B(n_154), .Y(n_187) );
INVx1_ASAP7_75t_L g109 ( .A(n_19), .Y(n_109) );
INVx1_ASAP7_75t_L g551 ( .A(n_20), .Y(n_551) );
INVx1_ASAP7_75t_SL g474 ( .A(n_21), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_22), .B(n_155), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_23), .A2(n_136), .B(n_169), .Y(n_168) );
AOI221xp5_ASAP7_75t_SL g179 ( .A1(n_24), .A2(n_40), .B1(n_136), .B2(n_154), .C(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_25), .B(n_148), .Y(n_170) );
AOI33xp33_ASAP7_75t_L g511 ( .A1(n_26), .A2(n_53), .A3(n_202), .B1(n_208), .B2(n_512), .B3(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g775 ( .A(n_27), .Y(n_775) );
INVx1_ASAP7_75t_L g485 ( .A(n_28), .Y(n_485) );
OR2x2_ASAP7_75t_L g160 ( .A(n_29), .B(n_93), .Y(n_160) );
OA21x2_ASAP7_75t_L g193 ( .A1(n_29), .A2(n_93), .B(n_159), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_30), .B(n_144), .Y(n_191) );
INVxp67_ASAP7_75t_L g211 ( .A(n_31), .Y(n_211) );
AND2x2_ASAP7_75t_L g242 ( .A(n_32), .B(n_157), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_33), .B(n_200), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_34), .A2(n_136), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_35), .B(n_144), .Y(n_181) );
AND2x2_ASAP7_75t_L g137 ( .A(n_36), .B(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g152 ( .A(n_36), .B(n_141), .Y(n_152) );
INVx1_ASAP7_75t_L g207 ( .A(n_36), .Y(n_207) );
OR2x6_ASAP7_75t_L g107 ( .A(n_37), .B(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_38), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_39), .B(n_200), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_41), .A2(n_172), .B1(n_216), .B2(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_42), .B(n_543), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_43), .A2(n_83), .B1(n_136), .B2(n_205), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_44), .B(n_155), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_45), .B(n_148), .Y(n_240) );
INVx1_ASAP7_75t_L g781 ( .A(n_46), .Y(n_781) );
XNOR2xp5_ASAP7_75t_L g809 ( .A(n_47), .B(n_87), .Y(n_809) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_48), .B(n_192), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_49), .B(n_155), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_50), .Y(n_538) );
AND2x2_ASAP7_75t_L g229 ( .A(n_51), .B(n_157), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_52), .B(n_157), .Y(n_183) );
XOR2xp5_ASAP7_75t_L g801 ( .A(n_52), .B(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g818 ( .A(n_52), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_54), .B(n_155), .Y(n_503) );
INVx1_ASAP7_75t_L g140 ( .A(n_55), .Y(n_140) );
INVx1_ASAP7_75t_L g150 ( .A(n_55), .Y(n_150) );
AND2x2_ASAP7_75t_L g504 ( .A(n_56), .B(n_157), .Y(n_504) );
AOI221xp5_ASAP7_75t_L g523 ( .A1(n_57), .A2(n_76), .B1(n_200), .B2(n_205), .C(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_58), .B(n_200), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_59), .B(n_154), .Y(n_241) );
OAI22xp5_ASAP7_75t_SL g113 ( .A1(n_60), .A2(n_114), .B1(n_119), .B2(n_120), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_60), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_61), .B(n_216), .Y(n_494) );
AOI21xp5_ASAP7_75t_SL g463 ( .A1(n_62), .A2(n_205), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g161 ( .A(n_63), .B(n_157), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_64), .B(n_144), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_65), .B(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_SL g194 ( .A(n_66), .B(n_158), .Y(n_194) );
INVx1_ASAP7_75t_L g548 ( .A(n_67), .Y(n_548) );
XNOR2xp5_ASAP7_75t_L g116 ( .A(n_68), .B(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_69), .A2(n_136), .B(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g502 ( .A(n_70), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_71), .B(n_144), .Y(n_171) );
AND2x2_ASAP7_75t_SL g279 ( .A(n_72), .B(n_192), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_73), .A2(n_205), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g138 ( .A(n_74), .Y(n_138) );
INVx1_ASAP7_75t_L g146 ( .A(n_74), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_75), .B(n_200), .Y(n_514) );
AND2x2_ASAP7_75t_L g476 ( .A(n_77), .B(n_215), .Y(n_476) );
INVx1_ASAP7_75t_L g549 ( .A(n_78), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_79), .A2(n_205), .B(n_473), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_80), .A2(n_205), .B(n_275), .C(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_81), .B(n_154), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_82), .A2(n_86), .B1(n_154), .B2(n_200), .Y(n_277) );
INVx1_ASAP7_75t_L g110 ( .A(n_84), .Y(n_110) );
AND2x2_ASAP7_75t_SL g461 ( .A(n_85), .B(n_215), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_88), .A2(n_205), .B1(n_509), .B2(n_510), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_89), .B(n_148), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_90), .B(n_148), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g815 ( .A(n_91), .B(n_816), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_92), .A2(n_136), .B(n_142), .Y(n_135) );
INVx1_ASAP7_75t_L g465 ( .A(n_94), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_95), .B(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g515 ( .A(n_96), .B(n_215), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_97), .A2(n_483), .B(n_484), .C(n_486), .Y(n_482) );
INVxp67_ASAP7_75t_L g214 ( .A(n_98), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_99), .B(n_154), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_100), .B(n_144), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_101), .A2(n_136), .B(n_189), .Y(n_188) );
BUFx2_ASAP7_75t_L g791 ( .A(n_102), .Y(n_791) );
BUFx2_ASAP7_75t_SL g822 ( .A(n_102), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_103), .B(n_155), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_783), .B1(n_794), .B2(n_796), .C(n_817), .Y(n_104) );
OAI31xp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_111), .A3(n_777), .B(n_779), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_106), .B(n_124), .Y(n_793) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g782 ( .A(n_107), .B(n_124), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_112), .B(n_121), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_113), .B(n_778), .Y(n_777) );
INVxp33_ASAP7_75t_L g120 ( .A(n_114), .Y(n_120) );
INVx1_ASAP7_75t_L g118 ( .A(n_116), .Y(n_118) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g778 ( .A(n_122), .Y(n_778) );
OAI21x1_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_125), .B(n_451), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g776 ( .A(n_124), .Y(n_776) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_390), .Y(n_125) );
NOR3xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_283), .C(n_334), .Y(n_126) );
OAI211xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_173), .B(n_230), .C(n_261), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_162), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_132), .B(n_235), .Y(n_398) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g243 ( .A(n_133), .B(n_164), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_133), .B(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g260 ( .A(n_133), .B(n_250), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_133), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g297 ( .A(n_133), .B(n_273), .Y(n_297) );
INVx2_ASAP7_75t_L g323 ( .A(n_133), .Y(n_323) );
AND2x4_ASAP7_75t_L g332 ( .A(n_133), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g437 ( .A(n_133), .B(n_304), .Y(n_437) );
AO21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_156), .B(n_161), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_153), .Y(n_134) );
AND2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
BUFx3_ASAP7_75t_L g204 ( .A(n_137), .Y(n_204) );
AND2x6_ASAP7_75t_L g148 ( .A(n_138), .B(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g209 ( .A(n_138), .Y(n_209) );
AND2x4_ASAP7_75t_L g205 ( .A(n_139), .B(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x4_ASAP7_75t_L g144 ( .A(n_140), .B(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g202 ( .A(n_140), .Y(n_202) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_141), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_147), .B(n_151), .Y(n_142) );
INVxp67_ASAP7_75t_L g554 ( .A(n_144), .Y(n_554) );
AND2x4_ASAP7_75t_L g155 ( .A(n_145), .B(n_149), .Y(n_155) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVxp67_ASAP7_75t_L g552 ( .A(n_148), .Y(n_552) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_151), .A2(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_151), .A2(n_181), .B(n_182), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_151), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_151), .A2(n_226), .B(n_227), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_151), .A2(n_239), .B(n_240), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g464 ( .A1(n_151), .A2(n_465), .B(n_466), .C(n_467), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_SL g473 ( .A1(n_151), .A2(n_466), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_151), .A2(n_466), .B(n_502), .C(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g509 ( .A(n_151), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_SL g524 ( .A1(n_151), .A2(n_466), .B(n_525), .C(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_151), .A2(n_541), .B(n_542), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_151), .B(n_172), .Y(n_555) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x4_ASAP7_75t_L g154 ( .A(n_152), .B(n_155), .Y(n_154) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_152), .Y(n_486) );
INVx1_ASAP7_75t_L g219 ( .A(n_155), .Y(n_219) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_156), .A2(n_236), .B(n_242), .Y(n_235) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_156), .A2(n_236), .B(n_242), .Y(n_250) );
AO21x2_ASAP7_75t_L g469 ( .A1(n_156), .A2(n_470), .B(n_476), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_157), .Y(n_156) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_157), .A2(n_179), .B(n_183), .Y(n_178) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_159), .B(n_160), .Y(n_158) );
AND2x4_ASAP7_75t_L g172 ( .A(n_159), .B(n_160), .Y(n_172) );
AND2x2_ASAP7_75t_L g321 ( .A(n_162), .B(n_322), .Y(n_321) );
OAI32xp33_ASAP7_75t_L g404 ( .A1(n_162), .A2(n_326), .A3(n_330), .B1(n_337), .B2(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_162), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g258 ( .A(n_163), .B(n_259), .Y(n_258) );
NAND3xp33_ASAP7_75t_L g331 ( .A(n_163), .B(n_253), .C(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g357 ( .A(n_163), .B(n_260), .Y(n_357) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_164), .Y(n_247) );
INVx5_ASAP7_75t_L g282 ( .A(n_164), .Y(n_282) );
AND2x4_ASAP7_75t_L g338 ( .A(n_164), .B(n_250), .Y(n_338) );
OR2x2_ASAP7_75t_L g353 ( .A(n_164), .B(n_273), .Y(n_353) );
OR2x2_ASAP7_75t_L g379 ( .A(n_164), .B(n_235), .Y(n_379) );
AND2x2_ASAP7_75t_L g387 ( .A(n_164), .B(n_333), .Y(n_387) );
AND2x4_ASAP7_75t_SL g412 ( .A(n_164), .B(n_332), .Y(n_412) );
OR2x6_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_172), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_172), .B(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_172), .B(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_172), .B(n_214), .Y(n_213) );
NOR3xp33_ASAP7_75t_L g217 ( .A(n_172), .B(n_218), .C(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_172), .A2(n_463), .B(n_468), .Y(n_462) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_174), .B(n_332), .Y(n_408) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_184), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_175), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
OR2x6_ASAP7_75t_SL g232 ( .A(n_176), .B(n_233), .Y(n_232) );
INVxp67_ASAP7_75t_SL g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g257 ( .A(n_177), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_177), .B(n_292), .Y(n_310) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_177), .Y(n_448) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g265 ( .A(n_178), .Y(n_265) );
AND2x2_ASAP7_75t_L g290 ( .A(n_178), .B(n_221), .Y(n_290) );
INVx2_ASAP7_75t_L g318 ( .A(n_178), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_178), .B(n_185), .Y(n_359) );
BUFx3_ASAP7_75t_L g383 ( .A(n_178), .Y(n_383) );
OR2x2_ASAP7_75t_L g395 ( .A(n_178), .B(n_185), .Y(n_395) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_178), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_184), .A2(n_426), .B1(n_429), .B2(n_430), .Y(n_425) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_195), .Y(n_184) );
INVx1_ASAP7_75t_L g253 ( .A(n_185), .Y(n_253) );
OR2x2_ASAP7_75t_L g264 ( .A(n_185), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g271 ( .A(n_185), .Y(n_271) );
AND2x4_ASAP7_75t_SL g288 ( .A(n_185), .B(n_196), .Y(n_288) );
AND2x4_ASAP7_75t_L g293 ( .A(n_185), .B(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g302 ( .A(n_185), .Y(n_302) );
OR2x2_ASAP7_75t_L g308 ( .A(n_185), .B(n_196), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_185), .B(n_310), .Y(n_309) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_185), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_185), .B(n_290), .Y(n_424) );
OR2x2_ASAP7_75t_L g440 ( .A(n_185), .B(n_343), .Y(n_440) );
OR2x6_ASAP7_75t_L g185 ( .A(n_186), .B(n_194), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_192), .Y(n_186) );
INVx2_ASAP7_75t_SL g275 ( .A(n_192), .Y(n_275) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_192), .A2(n_523), .B(n_527), .Y(n_522) );
BUFx4f_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx3_ASAP7_75t_L g216 ( .A(n_193), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_195), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g266 ( .A(n_195), .Y(n_266) );
AND2x2_ASAP7_75t_SL g373 ( .A(n_195), .B(n_257), .Y(n_373) );
AND2x4_ASAP7_75t_L g195 ( .A(n_196), .B(n_220), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_196), .B(n_221), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_196), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_196), .B(n_265), .Y(n_269) );
INVx3_ASAP7_75t_L g294 ( .A(n_196), .Y(n_294) );
INVx1_ASAP7_75t_L g327 ( .A(n_196), .Y(n_327) );
AND2x2_ASAP7_75t_L g407 ( .A(n_196), .B(n_271), .Y(n_407) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_212), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_200), .B1(n_205), .B2(n_210), .Y(n_197) );
INVx1_ASAP7_75t_L g495 ( .A(n_200), .Y(n_495) );
AND2x4_ASAP7_75t_L g200 ( .A(n_201), .B(n_204), .Y(n_200) );
INVx1_ASAP7_75t_L g536 ( .A(n_201), .Y(n_536) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
OR2x6_ASAP7_75t_L g466 ( .A(n_202), .B(n_209), .Y(n_466) );
INVxp33_ASAP7_75t_L g512 ( .A(n_202), .Y(n_512) );
INVx1_ASAP7_75t_L g537 ( .A(n_204), .Y(n_537) );
INVxp67_ASAP7_75t_L g493 ( .A(n_205), .Y(n_493) );
NOR2x1p5_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
INVx1_ASAP7_75t_L g513 ( .A(n_208), .Y(n_513) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_215), .A2(n_482), .B1(n_487), .B2(n_488), .Y(n_481) );
INVx3_ASAP7_75t_L g488 ( .A(n_215), .Y(n_488) );
INVx4_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AOI21x1_ASAP7_75t_L g222 ( .A1(n_216), .A2(n_223), .B(n_229), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_216), .B(n_491), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_219), .B(n_485), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_219), .A2(n_466), .B1(n_548), .B2(n_549), .Y(n_547) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_221), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g292 ( .A(n_221), .Y(n_292) );
AND2x2_ASAP7_75t_L g317 ( .A(n_221), .B(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g343 ( .A(n_221), .B(n_265), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_221), .B(n_294), .Y(n_360) );
INVx1_ASAP7_75t_L g366 ( .A(n_221), .Y(n_366) );
INVx3_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_228), .Y(n_223) );
AOI222xp33_ASAP7_75t_SL g230 ( .A1(n_231), .A2(n_234), .B1(n_244), .B2(n_251), .C1(n_254), .C2(n_258), .Y(n_230) );
CKINVDCx16_ASAP7_75t_R g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_243), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_235), .B(n_304), .Y(n_355) );
AND2x4_ASAP7_75t_L g371 ( .A(n_235), .B(n_282), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_241), .Y(n_236) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_246), .B(n_248), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g296 ( .A(n_247), .B(n_297), .Y(n_296) );
AOI222xp33_ASAP7_75t_L g261 ( .A1(n_248), .A2(n_262), .B1(n_267), .B2(n_272), .C1(n_280), .C2(n_826), .Y(n_261) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g400 ( .A(n_249), .B(n_304), .Y(n_400) );
OR2x2_ASAP7_75t_L g443 ( .A(n_249), .B(n_349), .Y(n_443) );
AND2x2_ASAP7_75t_L g272 ( .A(n_250), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g333 ( .A(n_250), .Y(n_333) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_250), .Y(n_348) );
O2A1O1Ixp33_ASAP7_75t_L g361 ( .A1(n_251), .A2(n_362), .B(n_367), .C(n_368), .Y(n_361) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g389 ( .A(n_253), .Y(n_389) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g319 ( .A(n_258), .Y(n_319) );
AND2x2_ASAP7_75t_L g303 ( .A(n_259), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g312 ( .A(n_259), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OAI31xp33_ASAP7_75t_L g354 ( .A1(n_262), .A2(n_280), .A3(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
A2O1A1Ixp33_ASAP7_75t_L g356 ( .A1(n_263), .A2(n_313), .B(n_357), .C(n_358), .Y(n_356) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
OR2x2_ASAP7_75t_L g345 ( .A(n_264), .B(n_294), .Y(n_345) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
BUFx2_ASAP7_75t_L g313 ( .A(n_273), .Y(n_313) );
AND2x2_ASAP7_75t_L g322 ( .A(n_273), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_274), .Y(n_304) );
AOI21x1_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B(n_279), .Y(n_274) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_275), .A2(n_507), .B(n_515), .Y(n_506) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_275), .A2(n_507), .B(n_515), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_282), .B(n_339), .Y(n_431) );
OAI211xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_295), .B(n_298), .C(n_320), .Y(n_283) );
INVxp33_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_286), .B(n_291), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g324 ( .A(n_288), .B(n_317), .Y(n_324) );
OR2x2_ASAP7_75t_L g300 ( .A(n_289), .B(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g330 ( .A(n_289), .B(n_304), .Y(n_330) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g406 ( .A(n_290), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g429 ( .A(n_291), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_293), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_293), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g441 ( .A(n_293), .B(n_317), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_293), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g384 ( .A(n_294), .B(n_366), .Y(n_384) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AOI322xp5_ASAP7_75t_L g438 ( .A1(n_297), .A2(n_317), .A3(n_371), .B1(n_396), .B2(n_439), .C1(n_441), .C2(n_442), .Y(n_438) );
AOI211xp5_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_303), .B(n_305), .C(n_314), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_301), .B(n_329), .Y(n_351) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g316 ( .A(n_302), .B(n_317), .Y(n_316) );
NOR2x1p5_ASAP7_75t_L g382 ( .A(n_302), .B(n_383), .Y(n_382) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_302), .Y(n_415) );
O2A1O1Ixp33_ASAP7_75t_L g320 ( .A1(n_303), .A2(n_321), .B(n_324), .C(n_325), .Y(n_320) );
AND2x4_ASAP7_75t_L g339 ( .A(n_304), .B(n_323), .Y(n_339) );
INVx2_ASAP7_75t_L g349 ( .A(n_304), .Y(n_349) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_304), .B(n_338), .Y(n_369) );
AND2x2_ASAP7_75t_L g411 ( .A(n_304), .B(n_412), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_304), .B(n_428), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_304), .B(n_332), .Y(n_450) );
AOI21xp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_309), .B(n_311), .Y(n_305) );
AND2x2_ASAP7_75t_L g401 ( .A(n_307), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g329 ( .A(n_310), .Y(n_329) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_319), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_322), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g416 ( .A(n_322), .Y(n_416) );
O2A1O1Ixp33_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_328), .B(n_330), .C(n_331), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_329), .Y(n_413) );
INVx3_ASAP7_75t_SL g428 ( .A(n_332), .Y(n_428) );
NAND5xp2_ASAP7_75t_L g334 ( .A(n_335), .B(n_354), .C(n_361), .D(n_374), .E(n_385), .Y(n_334) );
AOI222xp33_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_340), .B1(n_344), .B2(n_346), .C1(n_350), .C2(n_352), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_337), .A2(n_418), .B1(n_422), .B2(n_423), .Y(n_417) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g367 ( .A(n_338), .B(n_339), .Y(n_367) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_348), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_349), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g386 ( .A(n_349), .B(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g397 ( .A(n_349), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g427 ( .A(n_353), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g375 ( .A(n_360), .Y(n_375) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI21xp33_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B(n_372), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_371), .A2(n_375), .B1(n_376), .B2(n_380), .Y(n_374) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_371), .Y(n_422) );
INVx2_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g388 ( .A(n_373), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g393 ( .A(n_375), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVx1_ASAP7_75t_SL g421 ( .A(n_384), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
NOR3xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_409), .C(n_432), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_392), .B(n_408), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_396), .B1(n_399), .B2(n_401), .C(n_404), .Y(n_392) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g433 ( .A(n_395), .B(n_421), .Y(n_433) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
OAI321xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_413), .A3(n_414), .B1(n_416), .B2(n_417), .C(n_425), .Y(n_409) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_423), .A2(n_445), .B1(n_449), .B2(n_450), .Y(n_444) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI211xp5_ASAP7_75t_SL g432 ( .A1(n_433), .A2(n_434), .B(n_438), .C(n_444), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVxp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NOR2x1_ASAP7_75t_L g451 ( .A(n_452), .B(n_772), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_722), .Y(n_452) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_662), .B(n_721), .Y(n_453) );
NOR3xp33_ASAP7_75t_L g772 ( .A(n_454), .B(n_723), .C(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g812 ( .A(n_454), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_626), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_567), .C(n_596), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_457), .B(n_556), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_477), .B1(n_516), .B2(n_528), .Y(n_457) );
NAND2x1_ASAP7_75t_L g758 ( .A(n_458), .B(n_557), .Y(n_758) );
INVx2_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_469), .Y(n_459) );
INVx2_ASAP7_75t_L g530 ( .A(n_460), .Y(n_530) );
INVx4_ASAP7_75t_L g572 ( .A(n_460), .Y(n_572) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_460), .Y(n_592) );
AND2x4_ASAP7_75t_L g603 ( .A(n_460), .B(n_571), .Y(n_603) );
AND2x2_ASAP7_75t_L g609 ( .A(n_460), .B(n_533), .Y(n_609) );
NOR2x1_ASAP7_75t_SL g682 ( .A(n_460), .B(n_544), .Y(n_682) );
OR2x6_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVxp67_ASAP7_75t_L g483 ( .A(n_466), .Y(n_483) );
INVx2_ASAP7_75t_L g543 ( .A(n_466), .Y(n_543) );
INVx2_ASAP7_75t_L g575 ( .A(n_469), .Y(n_575) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_469), .Y(n_589) );
INVx1_ASAP7_75t_L g600 ( .A(n_469), .Y(n_600) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_469), .Y(n_612) );
AND2x2_ASAP7_75t_L g644 ( .A(n_469), .B(n_544), .Y(n_644) );
INVx1_ASAP7_75t_L g670 ( .A(n_469), .Y(n_670) );
AND2x2_ASAP7_75t_L g732 ( .A(n_469), .B(n_560), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_496), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g625 ( .A(n_479), .B(n_564), .Y(n_625) );
INVx2_ASAP7_75t_L g667 ( .A(n_479), .Y(n_667) );
AND2x2_ASAP7_75t_L g769 ( .A(n_479), .B(n_496), .Y(n_769) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_480), .B(n_519), .Y(n_563) );
INVx2_ASAP7_75t_L g584 ( .A(n_480), .Y(n_584) );
AND2x4_ASAP7_75t_L g606 ( .A(n_480), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g641 ( .A(n_480), .Y(n_641) );
AND2x2_ASAP7_75t_L g765 ( .A(n_480), .B(n_522), .Y(n_765) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_489), .Y(n_480) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_488), .A2(n_498), .B(n_504), .Y(n_497) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_488), .A2(n_498), .B(n_504), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_493), .B1(n_494), .B2(n_495), .Y(n_489) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g739 ( .A(n_496), .Y(n_739) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_505), .Y(n_496) );
NOR2xp67_ASAP7_75t_L g614 ( .A(n_497), .B(n_584), .Y(n_614) );
AND2x2_ASAP7_75t_L g619 ( .A(n_497), .B(n_584), .Y(n_619) );
INVx2_ASAP7_75t_L g632 ( .A(n_497), .Y(n_632) );
NOR2x1_ASAP7_75t_L g697 ( .A(n_497), .B(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
AND2x4_ASAP7_75t_L g605 ( .A(n_505), .B(n_518), .Y(n_605) );
AND2x2_ASAP7_75t_L g620 ( .A(n_505), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g675 ( .A(n_505), .Y(n_675) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_506), .B(n_522), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_506), .B(n_519), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_508), .B(n_514), .Y(n_507) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVxp33_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
INVx3_ASAP7_75t_L g581 ( .A(n_518), .Y(n_581) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_519), .Y(n_579) );
AND2x2_ASAP7_75t_L g693 ( .A(n_519), .B(n_694), .Y(n_693) );
INVx3_ASAP7_75t_L g636 ( .A(n_520), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_520), .B(n_675), .Y(n_716) );
BUFx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g583 ( .A(n_521), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x4_ASAP7_75t_L g564 ( .A(n_522), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g607 ( .A(n_522), .Y(n_607) );
INVxp67_ASAP7_75t_L g621 ( .A(n_522), .Y(n_621) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_522), .Y(n_694) );
INVx1_ASAP7_75t_L g698 ( .A(n_522), .Y(n_698) );
INVx1_ASAP7_75t_L g676 ( .A(n_528), .Y(n_676) );
NOR2x1_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
NOR2x1_ASAP7_75t_L g653 ( .A(n_529), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g718 ( .A(n_530), .B(n_559), .Y(n_718) );
OR2x2_ASAP7_75t_L g770 ( .A(n_531), .B(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g669 ( .A(n_532), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g705 ( .A(n_532), .B(n_592), .Y(n_705) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_544), .Y(n_532) );
AND2x4_ASAP7_75t_L g559 ( .A(n_533), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g571 ( .A(n_533), .Y(n_571) );
INVx2_ASAP7_75t_L g588 ( .A(n_533), .Y(n_588) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_533), .Y(n_714) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_539), .Y(n_533) );
NOR3xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .C(n_538), .Y(n_535) );
INVx3_ASAP7_75t_L g560 ( .A(n_544), .Y(n_560) );
INVx2_ASAP7_75t_L g654 ( .A(n_544), .Y(n_654) );
AND2x4_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_550), .B(n_555), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_552), .B1(n_553), .B2(n_554), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_561), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_558), .B(n_634), .Y(n_651) );
NOR2x1_ASAP7_75t_L g743 ( .A(n_558), .B(n_572), .Y(n_743) );
INVx4_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_559), .B(n_634), .Y(n_720) );
AND2x2_ASAP7_75t_L g587 ( .A(n_560), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g601 ( .A(n_560), .Y(n_601) );
AOI22xp5_ASAP7_75t_SL g649 ( .A1(n_561), .A2(n_650), .B1(n_651), .B2(n_652), .Y(n_649) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
NAND2x1p5_ASAP7_75t_L g646 ( .A(n_562), .B(n_620), .Y(n_646) );
INVx2_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g754 ( .A(n_563), .B(n_595), .Y(n_754) );
AND2x2_ASAP7_75t_L g577 ( .A(n_564), .B(n_578), .Y(n_577) );
AND2x4_ASAP7_75t_L g613 ( .A(n_564), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g756 ( .A(n_564), .B(n_667), .Y(n_756) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x4_ASAP7_75t_L g631 ( .A(n_566), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g657 ( .A(n_566), .Y(n_657) );
AND2x2_ASAP7_75t_L g692 ( .A(n_566), .B(n_584), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_576), .B1(n_580), .B2(n_585), .C(n_590), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .Y(n_569) );
INVx1_ASAP7_75t_L g648 ( .A(n_570), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_570), .B(n_644), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_570), .B(n_732), .Y(n_731) );
AND2x4_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NOR2xp67_ASAP7_75t_SL g616 ( .A(n_572), .B(n_617), .Y(n_616) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_572), .Y(n_629) );
AND2x4_ASAP7_75t_SL g713 ( .A(n_572), .B(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g760 ( .A(n_572), .B(n_761), .Y(n_760) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx3_ASAP7_75t_L g634 ( .A(n_574), .Y(n_634) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_575), .Y(n_771) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AOI221x1_ASAP7_75t_L g724 ( .A1(n_577), .A2(n_725), .B1(n_727), .B2(n_728), .C(n_730), .Y(n_724) );
AND2x2_ASAP7_75t_L g650 ( .A(n_578), .B(n_606), .Y(n_650) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AND2x2_ASAP7_75t_L g593 ( .A(n_581), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_581), .B(n_583), .Y(n_767) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
AND2x2_ASAP7_75t_SL g591 ( .A(n_587), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_587), .B(n_600), .Y(n_617) );
INVx2_ASAP7_75t_L g624 ( .A(n_587), .Y(n_624) );
INVx1_ASAP7_75t_L g686 ( .A(n_588), .Y(n_686) );
BUFx2_ASAP7_75t_L g706 ( .A(n_589), .Y(n_706) );
NAND2xp33_ASAP7_75t_SL g590 ( .A(n_591), .B(n_593), .Y(n_590) );
OR2x6_ASAP7_75t_L g623 ( .A(n_592), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g752 ( .A(n_592), .B(n_644), .Y(n_752) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_615), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_604), .B1(n_608), .B2(n_613), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .Y(n_598) );
AND2x2_ASAP7_75t_SL g661 ( .A(n_599), .B(n_603), .Y(n_661) );
AND2x4_ASAP7_75t_L g727 ( .A(n_599), .B(n_685), .Y(n_727) );
AND2x4_ASAP7_75t_SL g599 ( .A(n_600), .B(n_601), .Y(n_599) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_600), .Y(n_742) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_603), .B(n_643), .Y(n_642) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_603), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_603), .B(n_634), .Y(n_726) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
AND2x2_ASAP7_75t_L g747 ( .A(n_605), .B(n_666), .Y(n_747) );
INVx3_ASAP7_75t_L g658 ( .A(n_606), .Y(n_658) );
AND2x2_ASAP7_75t_L g679 ( .A(n_606), .B(n_631), .Y(n_679) );
NAND2x1_ASAP7_75t_SL g750 ( .A(n_606), .B(n_657), .Y(n_750) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_618), .B1(n_622), .B2(n_625), .Y(n_615) );
BUFx2_ASAP7_75t_L g671 ( .A(n_617), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_618), .A2(n_709), .B1(n_718), .B2(n_719), .Y(n_717) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
NAND2x1p5_ASAP7_75t_L g674 ( .A(n_619), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g639 ( .A(n_620), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND3xp33_ASAP7_75t_L g703 ( .A(n_624), .B(n_704), .C(n_706), .Y(n_703) );
INVx1_ASAP7_75t_L g659 ( .A(n_625), .Y(n_659) );
AOI211x1_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_635), .B(n_637), .C(n_655), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g737 ( .A(n_630), .B(n_718), .Y(n_737) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_631), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g709 ( .A(n_631), .B(n_667), .Y(n_709) );
AND2x2_ASAP7_75t_L g764 ( .A(n_631), .B(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g687 ( .A(n_634), .Y(n_687) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g729 ( .A(n_636), .B(n_674), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_649), .Y(n_637) );
AOI22xp5_ASAP7_75t_SL g638 ( .A1(n_639), .A2(n_642), .B1(n_645), .B2(n_647), .Y(n_638) );
BUFx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g702 ( .A(n_641), .B(n_697), .Y(n_702) );
INVx1_ASAP7_75t_SL g744 ( .A(n_641), .Y(n_744) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_SL g712 ( .A(n_644), .B(n_713), .Y(n_712) );
INVx3_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVxp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g748 ( .A(n_653), .B(n_670), .Y(n_748) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_659), .B(n_660), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_657), .B(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g672 ( .A(n_658), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVxp67_ASAP7_75t_SL g814 ( .A(n_662), .Y(n_814) );
NAND3x1_ASAP7_75t_L g662 ( .A(n_663), .B(n_699), .C(n_707), .Y(n_662) );
NAND4xp25_ASAP7_75t_L g773 ( .A(n_663), .B(n_699), .C(n_707), .D(n_774), .Y(n_773) );
NOR2x1_ASAP7_75t_L g663 ( .A(n_664), .B(n_677), .Y(n_663) );
OAI222xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_668), .B1(n_671), .B2(n_672), .C1(n_674), .C2(n_676), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OAI21xp5_ASAP7_75t_SL g751 ( .A1(n_669), .A2(n_752), .B(n_753), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g734 ( .A(n_670), .B(n_685), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_673), .A2(n_731), .B1(n_733), .B2(n_734), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_688), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_679), .B(n_680), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_681), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_687), .Y(n_683) );
INVx2_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_685), .B(n_687), .Y(n_690) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B1(n_695), .B2(n_696), .Y(n_688) );
AND2x4_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
AND2x2_ASAP7_75t_L g696 ( .A(n_692), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_700), .B(n_703), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g733 ( .A(n_702), .Y(n_733) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_717), .Y(n_707) );
AOI22xp5_ASAP7_75t_SL g708 ( .A1(n_709), .A2(n_710), .B1(n_712), .B2(n_715), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp33_ASAP7_75t_L g722 ( .A(n_721), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g813 ( .A(n_723), .Y(n_813) );
NAND3x1_ASAP7_75t_L g723 ( .A(n_724), .B(n_735), .C(n_755), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_727), .A2(n_747), .B1(n_748), .B2(n_749), .Y(n_746) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g761 ( .A(n_732), .Y(n_761) );
NOR2x1_ASAP7_75t_L g735 ( .A(n_736), .B(n_745), .Y(n_735) );
AOI21xp5_ASAP7_75t_SL g736 ( .A1(n_737), .A2(n_738), .B(n_744), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_751), .Y(n_745) );
INVx2_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_750), .B(n_763), .Y(n_762) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
AOI221xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B1(n_759), .B2(n_762), .C(n_766), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVxp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_768), .B(n_770), .Y(n_766) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_780), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_782), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_784), .Y(n_783) );
INVx2_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
AND2x2_ASAP7_75t_L g785 ( .A(n_786), .B(n_792), .Y(n_785) );
INVxp67_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NAND2xp5_ASAP7_75t_SL g787 ( .A(n_788), .B(n_791), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
OR2x2_ASAP7_75t_SL g795 ( .A(n_789), .B(n_791), .Y(n_795) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_789), .A2(n_820), .B(n_823), .Y(n_819) );
INVx1_ASAP7_75t_SL g816 ( .A(n_792), .Y(n_816) );
BUFx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
BUFx3_ASAP7_75t_L g800 ( .A(n_793), .Y(n_800) );
BUFx2_ASAP7_75t_L g824 ( .A(n_793), .Y(n_824) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
OAI21xp33_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_801), .B(n_815), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_798), .Y(n_797) );
CKINVDCx11_ASAP7_75t_R g798 ( .A(n_799), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_800), .Y(n_799) );
AOI22xp33_ASAP7_75t_SL g802 ( .A1(n_803), .A2(n_804), .B1(n_810), .B2(n_811), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_806), .B1(n_808), .B2(n_809), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
AND3x2_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .C(n_814), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .Y(n_817) );
CKINVDCx11_ASAP7_75t_R g820 ( .A(n_821), .Y(n_820) );
CKINVDCx8_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
endmodule