module fake_jpeg_9669_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_23),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_16),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_10),
.B1(n_9),
.B2(n_17),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_27),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_10),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_10),
.B(n_17),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_43),
.B(n_12),
.Y(n_51)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_11),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_41),
.B(n_42),
.Y(n_44)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_32),
.B1(n_13),
.B2(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_45),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_13),
.B1(n_16),
.B2(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_32),
.C(n_21),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_49),
.C(n_29),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_12),
.B(n_19),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_51),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_56),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_48),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_29),
.C(n_50),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_36),
.B1(n_52),
.B2(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_59),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_0),
.C(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_62),
.B(n_53),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_53),
.C(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_67),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_68),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_55),
.B1(n_62),
.B2(n_64),
.Y(n_71)
);

AOI322xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_29),
.A3(n_50),
.B1(n_5),
.B2(n_7),
.C1(n_3),
.C2(n_0),
.Y(n_73)
);

AO21x1_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_5),
.B(n_7),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_72),
.A2(n_73),
.B(n_71),
.Y(n_75)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_75),
.B(n_70),
.Y(n_76)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_2),
.B(n_3),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_2),
.Y(n_78)
);


endmodule