module fake_ibex_2025_n_958 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_958);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_958;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_328;
wire n_372;
wire n_293;
wire n_341;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_947;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_375;
wire n_340;
wire n_317;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_470;
wire n_276;
wire n_339;
wire n_259;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_918;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_444;
wire n_200;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_894;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_379;
wire n_320;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_450;
wire n_302;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_874;
wire n_890;
wire n_816;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_565;
wire n_424;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_298;
wire n_231;
wire n_202;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g185 ( 
.A(n_76),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_179),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_31),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_127),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_102),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_69),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_29),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_5),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_134),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_130),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_131),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_29),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_98),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_15),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_90),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_119),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_2),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_82),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_120),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_51),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_61),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_14),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_31),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_114),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_21),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_91),
.Y(n_218)
);

INVx4_ASAP7_75t_R g219 ( 
.A(n_115),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_148),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_25),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_22),
.Y(n_222)
);

NOR2xp67_ASAP7_75t_L g223 ( 
.A(n_180),
.B(n_43),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_168),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_56),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_107),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_64),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_41),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_5),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_73),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_93),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_101),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_62),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_8),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_151),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_156),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_172),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_97),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_111),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_74),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_11),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_22),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_65),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_75),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_146),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_10),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_94),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_171),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_23),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_175),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_33),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_123),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_135),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_42),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_92),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_144),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_78),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_67),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_176),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_174),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_55),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_169),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_153),
.Y(n_264)
);

INVxp33_ASAP7_75t_SL g265 ( 
.A(n_104),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_L g266 ( 
.A(n_66),
.B(n_14),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_57),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_34),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_1),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_125),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_52),
.B(n_161),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_173),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_37),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_100),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_87),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_18),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_126),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_40),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_11),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_41),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_42),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_117),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_54),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_124),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_59),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_12),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_20),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_77),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_45),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_23),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_154),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_13),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_181),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_159),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_116),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_86),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_121),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_106),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_88),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_53),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_89),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_166),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_132),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_133),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_68),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_145),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_139),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_8),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_143),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_186),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_229),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_216),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_247),
.B(n_0),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_0),
.Y(n_314)
);

BUFx8_ASAP7_75t_L g315 ( 
.A(n_213),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_255),
.B(n_1),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_216),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_186),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_229),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_250),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_250),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_257),
.Y(n_322)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_230),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_249),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_249),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_298),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_186),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_298),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_257),
.Y(n_329)
);

OA21x2_ASAP7_75t_L g330 ( 
.A1(n_185),
.A2(n_99),
.B(n_178),
.Y(n_330)
);

AND2x4_ASAP7_75t_L g331 ( 
.A(n_255),
.B(n_3),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_258),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_273),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_286),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_258),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_273),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_234),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_263),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_239),
.B(n_3),
.Y(n_339)
);

BUFx12f_ASAP7_75t_L g340 ( 
.A(n_216),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_263),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_207),
.B(n_4),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_263),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_212),
.B(n_4),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_263),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_280),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_270),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_270),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_285),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_290),
.B(n_6),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_256),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_280),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_281),
.Y(n_353)
);

CKINVDCx8_ASAP7_75t_R g354 ( 
.A(n_231),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_281),
.Y(n_355)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_256),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_191),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_192),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_195),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_256),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_308),
.B(n_6),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_212),
.B(n_7),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_193),
.B(n_7),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_198),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_308),
.B(n_9),
.Y(n_365)
);

CKINVDCx11_ASAP7_75t_R g366 ( 
.A(n_188),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g367 ( 
.A(n_199),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_203),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_200),
.B(n_9),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_204),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_206),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_202),
.B(n_10),
.Y(n_372)
);

OAI21x1_ASAP7_75t_L g373 ( 
.A1(n_208),
.A2(n_103),
.B(n_170),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_210),
.Y(n_374)
);

INVx6_ASAP7_75t_L g375 ( 
.A(n_283),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_217),
.B(n_12),
.Y(n_376)
);

AOI22x1_ASAP7_75t_SL g377 ( 
.A1(n_188),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_211),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_220),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_225),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_233),
.B(n_16),
.Y(n_381)
);

CKINVDCx11_ASAP7_75t_R g382 ( 
.A(n_214),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_235),
.Y(n_383)
);

AND2x6_ASAP7_75t_L g384 ( 
.A(n_236),
.B(n_238),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_241),
.Y(n_385)
);

NOR2x1p5_ASAP7_75t_L g386 ( 
.A(n_340),
.B(n_356),
.Y(n_386)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_316),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_363),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_314),
.A2(n_309),
.B1(n_189),
.B2(n_201),
.Y(n_389)
);

BUFx10_ASAP7_75t_L g390 ( 
.A(n_375),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_356),
.B(n_222),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_358),
.B(n_244),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_314),
.A2(n_309),
.B1(n_187),
.B2(n_189),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_369),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_369),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_317),
.B(n_196),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_375),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_327),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_316),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_375),
.Y(n_403)
);

OR2x6_ASAP7_75t_L g404 ( 
.A(n_340),
.B(n_228),
.Y(n_404)
);

BUFx10_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_372),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_317),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_358),
.B(n_245),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_316),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_334),
.Y(n_411)
);

AO21x2_ASAP7_75t_L g412 ( 
.A1(n_373),
.A2(n_253),
.B(n_248),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_317),
.B(n_197),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_331),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_317),
.B(n_299),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_323),
.B(n_265),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_323),
.B(n_265),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_331),
.Y(n_418)
);

INVx6_ASAP7_75t_L g419 ( 
.A(n_357),
.Y(n_419)
);

OR2x6_ASAP7_75t_L g420 ( 
.A(n_337),
.B(n_242),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_347),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_323),
.B(n_254),
.Y(n_422)
);

OR2x6_ASAP7_75t_L g423 ( 
.A(n_312),
.B(n_243),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_376),
.A2(n_344),
.B1(n_362),
.B2(n_364),
.Y(n_424)
);

AO22x2_ASAP7_75t_L g425 ( 
.A1(n_377),
.A2(n_287),
.B1(n_252),
.B2(n_214),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_364),
.B(n_260),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_376),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_315),
.Y(n_428)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_351),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_351),
.B(n_360),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_344),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_351),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_362),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_342),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_324),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_L g436 ( 
.A1(n_374),
.A2(n_269),
.B1(n_279),
.B2(n_268),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_348),
.Y(n_437)
);

INVx8_ASAP7_75t_L g438 ( 
.A(n_360),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_360),
.B(n_299),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_312),
.B(n_304),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_315),
.A2(n_201),
.B1(n_246),
.B2(n_187),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_325),
.Y(n_442)
);

INVxp33_ASAP7_75t_L g443 ( 
.A(n_366),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_315),
.A2(n_301),
.B1(n_288),
.B2(n_262),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_325),
.Y(n_445)
);

OAI22xp33_ASAP7_75t_L g446 ( 
.A1(n_354),
.A2(n_276),
.B1(n_288),
.B2(n_246),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_326),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_379),
.B(n_277),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_384),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_313),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_367),
.B(n_378),
.Y(n_451)
);

OR2x6_ASAP7_75t_L g452 ( 
.A(n_361),
.B(n_266),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_315),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_379),
.B(n_289),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_328),
.Y(n_455)
);

INVx8_ASAP7_75t_L g456 ( 
.A(n_384),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_383),
.B(n_291),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_354),
.B(n_304),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_365),
.A2(n_262),
.B1(n_301),
.B2(n_215),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_383),
.A2(n_194),
.B1(n_292),
.B2(n_221),
.Y(n_460)
);

AND2x6_ASAP7_75t_L g461 ( 
.A(n_368),
.B(n_294),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_368),
.B(n_295),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_380),
.B(n_190),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_327),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_380),
.B(n_296),
.Y(n_465)
);

BUFx24_ASAP7_75t_SL g466 ( 
.A(n_441),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_390),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_450),
.B(n_384),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_390),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_416),
.B(n_339),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_389),
.A2(n_276),
.B1(n_382),
.B2(n_377),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_417),
.B(n_391),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_391),
.B(n_359),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_435),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_430),
.A2(n_384),
.B(n_373),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_L g476 ( 
.A(n_456),
.B(n_384),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_359),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_429),
.B(n_384),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_442),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_411),
.Y(n_480)
);

OAI22xp33_ASAP7_75t_L g481 ( 
.A1(n_433),
.A2(n_350),
.B1(n_385),
.B2(n_380),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_393),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_449),
.B(n_357),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_456),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_449),
.B(n_357),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_414),
.A2(n_385),
.B1(n_328),
.B2(n_371),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_398),
.B(n_381),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_413),
.B(n_311),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_438),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_456),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_L g491 ( 
.A(n_441),
.B(n_329),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_405),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_405),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_422),
.B(n_332),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_423),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_433),
.B(n_335),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_434),
.B(n_335),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_438),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_434),
.B(n_319),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_438),
.B(n_319),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_419),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_415),
.B(n_320),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_410),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_387),
.B(n_370),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_387),
.B(n_370),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_451),
.B(n_320),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_388),
.A2(n_330),
.B(n_305),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_431),
.B(n_407),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_432),
.B(n_321),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_418),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_439),
.B(n_321),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_445),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_387),
.B(n_370),
.Y(n_513)
);

O2A1O1Ixp33_ASAP7_75t_L g514 ( 
.A1(n_427),
.A2(n_408),
.B(n_426),
.C(n_394),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_420),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_447),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_420),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_461),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_423),
.B(n_333),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_420),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_455),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_394),
.B(n_336),
.Y(n_522)
);

OAI22xp33_ASAP7_75t_L g523 ( 
.A1(n_389),
.A2(n_355),
.B1(n_353),
.B2(n_352),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_392),
.A2(n_353),
.B1(n_352),
.B2(n_336),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_408),
.B(n_346),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_426),
.B(n_346),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_421),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_428),
.B(n_370),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_448),
.B(n_205),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_396),
.B(n_370),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_448),
.B(n_209),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_386),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_440),
.B(n_300),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_404),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_437),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_458),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_459),
.B(n_371),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_454),
.B(n_224),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_397),
.B(n_399),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_457),
.B(n_226),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_463),
.B(n_302),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_402),
.Y(n_542)
);

NOR2x1_ASAP7_75t_R g543 ( 
.A(n_443),
.B(n_227),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_402),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_457),
.B(n_232),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_462),
.B(n_237),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_462),
.B(n_240),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_409),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_400),
.B(n_303),
.Y(n_549)
);

BUFx6f_ASAP7_75t_SL g550 ( 
.A(n_404),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_470),
.B(n_499),
.Y(n_551)
);

OA22x2_ASAP7_75t_L g552 ( 
.A1(n_466),
.A2(n_444),
.B1(n_395),
.B2(n_459),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_503),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_480),
.B(n_395),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_503),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_489),
.B(n_406),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_509),
.Y(n_557)
);

AO22x1_ASAP7_75t_L g558 ( 
.A1(n_517),
.A2(n_446),
.B1(n_444),
.B2(n_461),
.Y(n_558)
);

OAI21xp33_ASAP7_75t_L g559 ( 
.A1(n_472),
.A2(n_460),
.B(n_436),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_539),
.A2(n_409),
.B(n_412),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_542),
.Y(n_561)
);

BUFx12f_ASAP7_75t_L g562 ( 
.A(n_532),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_536),
.A2(n_452),
.B1(n_403),
.B2(n_461),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_468),
.A2(n_412),
.B(n_465),
.Y(n_564)
);

AOI21x1_ASAP7_75t_L g565 ( 
.A1(n_507),
.A2(n_465),
.B(n_330),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_515),
.B(n_520),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_544),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_514),
.A2(n_330),
.B(n_452),
.Y(n_568)
);

CKINVDCx10_ASAP7_75t_R g569 ( 
.A(n_550),
.Y(n_569)
);

NOR2x1_ASAP7_75t_L g570 ( 
.A(n_537),
.B(n_271),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_481),
.B(n_371),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_481),
.B(n_371),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_L g573 ( 
.A(n_490),
.B(n_251),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_497),
.B(n_519),
.Y(n_574)
);

O2A1O1Ixp5_ASAP7_75t_SL g575 ( 
.A1(n_504),
.A2(n_306),
.B(n_307),
.C(n_219),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_473),
.B(n_371),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_478),
.A2(n_218),
.B(n_223),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_548),
.Y(n_578)
);

O2A1O1Ixp33_ASAP7_75t_L g579 ( 
.A1(n_523),
.A2(n_267),
.B(n_310),
.C(n_318),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_473),
.B(n_371),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_475),
.A2(n_349),
.B(n_464),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_489),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_491),
.A2(n_425),
.B1(n_259),
.B2(n_261),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_498),
.B(n_264),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_498),
.A2(n_425),
.B1(n_272),
.B2(n_274),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_529),
.B(n_531),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_508),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_495),
.B(n_17),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_534),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_538),
.B(n_275),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_540),
.B(n_282),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_545),
.B(n_284),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_518),
.B(n_293),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_474),
.Y(n_594)
);

AO22x1_ASAP7_75t_L g595 ( 
.A1(n_467),
.A2(n_297),
.B1(n_19),
.B2(n_24),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_522),
.B(n_18),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_479),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_525),
.B(n_19),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_477),
.B(n_24),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_510),
.A2(n_310),
.B1(n_338),
.B2(n_343),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_523),
.B(n_469),
.Y(n_601)
);

BUFx6f_ASAP7_75t_SL g602 ( 
.A(n_492),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_490),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_526),
.B(n_25),
.Y(n_604)
);

CKINVDCx8_ASAP7_75t_R g605 ( 
.A(n_550),
.Y(n_605)
);

O2A1O1Ixp33_ASAP7_75t_L g606 ( 
.A1(n_496),
.A2(n_524),
.B(n_506),
.C(n_494),
.Y(n_606)
);

OR2x2_ASAP7_75t_SL g607 ( 
.A(n_471),
.B(n_26),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_493),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_546),
.B(n_26),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_500),
.A2(n_345),
.B1(n_341),
.B2(n_30),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_512),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_547),
.B(n_27),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_483),
.A2(n_401),
.B(n_345),
.Y(n_613)
);

AND3x2_ASAP7_75t_L g614 ( 
.A(n_543),
.B(n_27),
.C(n_28),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_L g615 ( 
.A1(n_488),
.A2(n_341),
.B(n_109),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_487),
.B(n_30),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_516),
.A2(n_341),
.B1(n_33),
.B2(n_34),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_490),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_485),
.A2(n_110),
.B(n_165),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_484),
.B(n_32),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_484),
.B(n_32),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_487),
.B(n_35),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_533),
.B(n_36),
.Y(n_623)
);

AO21x2_ASAP7_75t_L g624 ( 
.A1(n_504),
.A2(n_112),
.B(n_163),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_528),
.Y(n_625)
);

A2O1A1Ixp33_ASAP7_75t_L g626 ( 
.A1(n_488),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_502),
.A2(n_113),
.B(n_162),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_533),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_502),
.B(n_511),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_521),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_485),
.A2(n_118),
.B(n_44),
.Y(n_631)
);

A2O1A1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_511),
.A2(n_39),
.B(n_46),
.C(n_47),
.Y(n_632)
);

CKINVDCx14_ASAP7_75t_R g633 ( 
.A(n_541),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_549),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_535),
.Y(n_635)
);

AOI22x1_ASAP7_75t_L g636 ( 
.A1(n_535),
.A2(n_58),
.B1(n_60),
.B2(n_63),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_549),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_560),
.A2(n_476),
.B(n_530),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_551),
.B(n_486),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_587),
.Y(n_640)
);

AO32x2_ASAP7_75t_L g641 ( 
.A1(n_617),
.A2(n_513),
.A3(n_505),
.B1(n_530),
.B2(n_482),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_582),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_630),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_557),
.B(n_527),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_552),
.A2(n_501),
.B1(n_80),
.B2(n_81),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_594),
.Y(n_646)
);

AOI221x1_ASAP7_75t_L g647 ( 
.A1(n_615),
.A2(n_79),
.B1(n_83),
.B2(n_84),
.C(n_85),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_597),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_586),
.A2(n_95),
.B(n_96),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_589),
.B(n_182),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_554),
.B(n_108),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_611),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_601),
.B(n_559),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_629),
.A2(n_128),
.B(n_129),
.Y(n_654)
);

OA21x2_ASAP7_75t_L g655 ( 
.A1(n_565),
.A2(n_572),
.B(n_571),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_582),
.Y(n_656)
);

AND2x2_ASAP7_75t_SL g657 ( 
.A(n_588),
.B(n_582),
.Y(n_657)
);

CKINVDCx11_ASAP7_75t_R g658 ( 
.A(n_605),
.Y(n_658)
);

AO32x2_ASAP7_75t_L g659 ( 
.A1(n_610),
.A2(n_585),
.A3(n_600),
.B1(n_625),
.B2(n_575),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_588),
.B(n_136),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_603),
.Y(n_661)
);

AO31x2_ASAP7_75t_L g662 ( 
.A1(n_632),
.A2(n_137),
.A3(n_138),
.B(n_140),
.Y(n_662)
);

NOR2xp67_ASAP7_75t_L g663 ( 
.A(n_583),
.B(n_141),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_566),
.B(n_158),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_552),
.B(n_142),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_596),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_608),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_598),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_SL g669 ( 
.A1(n_603),
.A2(n_149),
.B(n_150),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_633),
.B(n_152),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_604),
.Y(n_671)
);

A2O1A1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_623),
.A2(n_157),
.B(n_622),
.C(n_616),
.Y(n_672)
);

NOR2x1_ASAP7_75t_SL g673 ( 
.A(n_603),
.B(n_618),
.Y(n_673)
);

AO31x2_ASAP7_75t_L g674 ( 
.A1(n_626),
.A2(n_577),
.A3(n_576),
.B(n_580),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_561),
.Y(n_675)
);

OAI21x1_ASAP7_75t_SL g676 ( 
.A1(n_563),
.A2(n_637),
.B(n_579),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_558),
.B(n_612),
.Y(n_677)
);

AO31x2_ASAP7_75t_L g678 ( 
.A1(n_619),
.A2(n_631),
.A3(n_613),
.B(n_567),
.Y(n_678)
);

INVx8_ASAP7_75t_L g679 ( 
.A(n_602),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_602),
.B(n_562),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_609),
.B(n_570),
.Y(n_681)
);

AO31x2_ASAP7_75t_L g682 ( 
.A1(n_578),
.A2(n_553),
.A3(n_555),
.B(n_591),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_628),
.Y(n_683)
);

OAI21x1_ASAP7_75t_SL g684 ( 
.A1(n_634),
.A2(n_636),
.B(n_592),
.Y(n_684)
);

INVx5_ASAP7_75t_L g685 ( 
.A(n_635),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_595),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_590),
.B(n_556),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_620),
.B(n_621),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_584),
.A2(n_573),
.B1(n_593),
.B2(n_614),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_624),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_SL g691 ( 
.A1(n_569),
.A2(n_498),
.B(n_489),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_607),
.Y(n_692)
);

NOR2xp67_ASAP7_75t_L g693 ( 
.A(n_583),
.B(n_515),
.Y(n_693)
);

BUFx2_ASAP7_75t_R g694 ( 
.A(n_605),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_551),
.B(n_587),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_551),
.B(n_587),
.Y(n_696)
);

O2A1O1Ixp33_ASAP7_75t_SL g697 ( 
.A1(n_632),
.A2(n_622),
.B(n_616),
.C(n_627),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_551),
.B(n_587),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_551),
.B(n_587),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_551),
.B(n_587),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_551),
.B(n_587),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_587),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_560),
.A2(n_551),
.B(n_564),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_568),
.A2(n_564),
.B(n_560),
.Y(n_704)
);

CKINVDCx11_ASAP7_75t_R g705 ( 
.A(n_605),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_551),
.B(n_587),
.Y(n_706)
);

A2O1A1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_606),
.A2(n_514),
.B(n_586),
.C(n_568),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_587),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_587),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_551),
.B(n_587),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g711 ( 
.A1(n_568),
.A2(n_564),
.B(n_560),
.Y(n_711)
);

O2A1O1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_551),
.A2(n_559),
.B(n_622),
.C(n_616),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_582),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_582),
.B(n_480),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_551),
.B(n_587),
.Y(n_715)
);

INVx5_ASAP7_75t_L g716 ( 
.A(n_582),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_605),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_551),
.A2(n_433),
.B1(n_574),
.B2(n_424),
.Y(n_718)
);

OAI22x1_ASAP7_75t_L g719 ( 
.A1(n_583),
.A2(n_395),
.B1(n_389),
.B2(n_441),
.Y(n_719)
);

AO22x2_ASAP7_75t_L g720 ( 
.A1(n_588),
.A2(n_585),
.B1(n_377),
.B2(n_599),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_SL g721 ( 
.A1(n_607),
.A2(n_471),
.B1(n_444),
.B2(n_441),
.Y(n_721)
);

AO31x2_ASAP7_75t_L g722 ( 
.A1(n_568),
.A2(n_581),
.A3(n_572),
.B(n_571),
.Y(n_722)
);

AO22x2_ASAP7_75t_L g723 ( 
.A1(n_588),
.A2(n_585),
.B1(n_377),
.B2(n_599),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_582),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_SL g725 ( 
.A1(n_650),
.A2(n_707),
.B(n_649),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_640),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_661),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_655),
.Y(n_728)
);

BUFx2_ASAP7_75t_SL g729 ( 
.A(n_717),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_702),
.Y(n_730)
);

AO21x2_ASAP7_75t_L g731 ( 
.A1(n_684),
.A2(n_653),
.B(n_676),
.Y(n_731)
);

AOI21xp33_ASAP7_75t_L g732 ( 
.A1(n_712),
.A2(n_677),
.B(n_718),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_697),
.A2(n_672),
.B(n_638),
.Y(n_733)
);

NOR2x1_ASAP7_75t_SL g734 ( 
.A(n_716),
.B(n_661),
.Y(n_734)
);

INVxp67_ASAP7_75t_SL g735 ( 
.A(n_695),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_708),
.Y(n_736)
);

OA21x2_ASAP7_75t_L g737 ( 
.A1(n_647),
.A2(n_645),
.B(n_654),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_667),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_696),
.B(n_698),
.Y(n_739)
);

AOI21xp33_ASAP7_75t_L g740 ( 
.A1(n_681),
.A2(n_683),
.B(n_686),
.Y(n_740)
);

OAI21xp5_ASAP7_75t_L g741 ( 
.A1(n_699),
.A2(n_715),
.B(n_706),
.Y(n_741)
);

OAI21x1_ASAP7_75t_L g742 ( 
.A1(n_669),
.A2(n_660),
.B(n_690),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_700),
.B(n_701),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_709),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_710),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_716),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_643),
.B(n_644),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_646),
.B(n_716),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_648),
.B(n_652),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_661),
.Y(n_750)
);

BUFx2_ASAP7_75t_SL g751 ( 
.A(n_650),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_642),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_720),
.B(n_723),
.Y(n_753)
);

AO21x2_ASAP7_75t_L g754 ( 
.A1(n_666),
.A2(n_671),
.B(n_668),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_639),
.A2(n_687),
.B(n_688),
.Y(n_755)
);

OAI21xp5_ASAP7_75t_L g756 ( 
.A1(n_651),
.A2(n_665),
.B(n_663),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_719),
.B(n_714),
.Y(n_757)
);

CKINVDCx6p67_ASAP7_75t_R g758 ( 
.A(n_679),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_675),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_720),
.B(n_723),
.Y(n_760)
);

OA21x2_ASAP7_75t_L g761 ( 
.A1(n_722),
.A2(n_690),
.B(n_641),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_692),
.Y(n_762)
);

AOI21x1_ASAP7_75t_L g763 ( 
.A1(n_664),
.A2(n_693),
.B(n_656),
.Y(n_763)
);

OAI21x1_ASAP7_75t_SL g764 ( 
.A1(n_673),
.A2(n_689),
.B(n_657),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_664),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_682),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_721),
.B(n_691),
.Y(n_767)
);

INVx4_ASAP7_75t_L g768 ( 
.A(n_679),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_670),
.B(n_680),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_682),
.B(n_724),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_673),
.A2(n_685),
.B(n_642),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_685),
.A2(n_713),
.B1(n_694),
.B2(n_641),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_713),
.B(n_674),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_713),
.B(n_674),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_674),
.B(n_678),
.Y(n_775)
);

AO31x2_ASAP7_75t_L g776 ( 
.A1(n_662),
.A2(n_659),
.A3(n_658),
.B(n_705),
.Y(n_776)
);

AO21x2_ASAP7_75t_L g777 ( 
.A1(n_659),
.A2(n_711),
.B(n_704),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_662),
.B(n_695),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_640),
.Y(n_779)
);

AO21x1_ASAP7_75t_L g780 ( 
.A1(n_712),
.A2(n_653),
.B(n_703),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_695),
.B(n_696),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_695),
.B(n_696),
.Y(n_782)
);

AND2x2_ASAP7_75t_SL g783 ( 
.A(n_657),
.B(n_650),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_661),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_721),
.A2(n_683),
.B1(n_692),
.B2(n_552),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_695),
.B(n_696),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_695),
.B(n_696),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_695),
.B(n_696),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_667),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_695),
.B(n_696),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_758),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_790),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_728),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_739),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_735),
.B(n_782),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_782),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_735),
.B(n_743),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_766),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_786),
.B(n_781),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_745),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_746),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_746),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_759),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_748),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_786),
.B(n_741),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_787),
.B(n_788),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_751),
.B(n_785),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_785),
.B(n_757),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_749),
.B(n_754),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_749),
.B(n_753),
.Y(n_810)
);

AO21x2_ASAP7_75t_L g811 ( 
.A1(n_733),
.A2(n_780),
.B(n_732),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_773),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_726),
.Y(n_813)
);

NOR2x1_ASAP7_75t_L g814 ( 
.A(n_772),
.B(n_771),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_749),
.B(n_760),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_730),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_789),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_736),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_748),
.B(n_783),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_747),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_744),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_779),
.Y(n_822)
);

OR2x6_ASAP7_75t_L g823 ( 
.A(n_725),
.B(n_764),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_770),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_774),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_774),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_783),
.Y(n_827)
);

OR2x6_ASAP7_75t_L g828 ( 
.A(n_771),
.B(n_763),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_740),
.B(n_765),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_768),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_755),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_778),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_778),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_775),
.B(n_727),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_752),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_775),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_738),
.Y(n_837)
);

CKINVDCx10_ASAP7_75t_R g838 ( 
.A(n_729),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_752),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_762),
.B(n_767),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_798),
.Y(n_841)
);

AOI221xp5_ASAP7_75t_L g842 ( 
.A1(n_796),
.A2(n_756),
.B1(n_769),
.B2(n_768),
.C(n_777),
.Y(n_842)
);

OAI21xp33_ASAP7_75t_L g843 ( 
.A1(n_799),
.A2(n_727),
.B(n_750),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_827),
.A2(n_731),
.B1(n_784),
.B2(n_750),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_793),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_802),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_834),
.B(n_777),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_797),
.B(n_761),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_834),
.B(n_761),
.Y(n_849)
);

NOR2xp67_ASAP7_75t_L g850 ( 
.A(n_797),
.B(n_784),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_831),
.B(n_805),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_824),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_812),
.B(n_776),
.Y(n_853)
);

CKINVDCx14_ASAP7_75t_R g854 ( 
.A(n_791),
.Y(n_854)
);

OR2x2_ASAP7_75t_SL g855 ( 
.A(n_808),
.B(n_737),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_809),
.B(n_795),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_802),
.Y(n_857)
);

OR2x6_ASAP7_75t_L g858 ( 
.A(n_823),
.B(n_742),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_856),
.B(n_847),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_856),
.B(n_836),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_848),
.B(n_847),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_848),
.B(n_808),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_846),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_851),
.B(n_795),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_841),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_849),
.B(n_836),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_858),
.B(n_832),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_850),
.Y(n_868)
);

OR2x6_ASAP7_75t_L g869 ( 
.A(n_858),
.B(n_823),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_851),
.B(n_805),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_849),
.B(n_825),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_845),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_853),
.B(n_826),
.Y(n_873)
);

AOI21xp33_ASAP7_75t_L g874 ( 
.A1(n_843),
.A2(n_807),
.B(n_811),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_854),
.B(n_830),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_853),
.B(n_832),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_846),
.B(n_830),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_858),
.B(n_833),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_869),
.B(n_867),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_870),
.B(n_852),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_859),
.B(n_810),
.Y(n_881)
);

NOR2x1_ASAP7_75t_L g882 ( 
.A(n_875),
.B(n_846),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_865),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_868),
.B(n_843),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_861),
.B(n_852),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_872),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_859),
.B(n_810),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_861),
.B(n_807),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_865),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_860),
.B(n_815),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_862),
.B(n_817),
.Y(n_891)
);

OR2x6_ASAP7_75t_L g892 ( 
.A(n_869),
.B(n_858),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_862),
.B(n_837),
.Y(n_893)
);

NAND4xp25_ASAP7_75t_L g894 ( 
.A(n_874),
.B(n_842),
.C(n_840),
.D(n_850),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_860),
.B(n_815),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_881),
.B(n_866),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_888),
.B(n_876),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_885),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_887),
.B(n_866),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_883),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_886),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_879),
.B(n_871),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_889),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_880),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_893),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_893),
.B(n_876),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_884),
.A2(n_842),
.B(n_806),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_900),
.Y(n_908)
);

OAI21xp33_ASAP7_75t_L g909 ( 
.A1(n_904),
.A2(n_894),
.B(n_884),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_900),
.Y(n_910)
);

INVxp33_ASAP7_75t_L g911 ( 
.A(n_906),
.Y(n_911)
);

OAI32xp33_ASAP7_75t_L g912 ( 
.A1(n_906),
.A2(n_877),
.A3(n_891),
.B1(n_857),
.B2(n_888),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_907),
.A2(n_882),
.B(n_891),
.C(n_879),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_896),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_898),
.B(n_890),
.Y(n_915)
);

OAI22xp33_ASAP7_75t_SL g916 ( 
.A1(n_905),
.A2(n_892),
.B1(n_879),
.B2(n_869),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_SL g917 ( 
.A1(n_896),
.A2(n_863),
.B(n_819),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_897),
.A2(n_892),
.B(n_869),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_901),
.A2(n_892),
.B(n_869),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_917),
.A2(n_892),
.B1(n_902),
.B2(n_899),
.Y(n_920)
);

AOI222xp33_ASAP7_75t_L g921 ( 
.A1(n_909),
.A2(n_895),
.B1(n_903),
.B2(n_899),
.C1(n_792),
.C2(n_902),
.Y(n_921)
);

AOI21xp33_ASAP7_75t_SL g922 ( 
.A1(n_913),
.A2(n_874),
.B(n_838),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_918),
.A2(n_867),
.B1(n_878),
.B2(n_873),
.Y(n_923)
);

AOI332xp33_ASAP7_75t_L g924 ( 
.A1(n_908),
.A2(n_821),
.A3(n_822),
.B1(n_818),
.B2(n_816),
.B3(n_813),
.C1(n_864),
.C2(n_806),
.Y(n_924)
);

AOI211xp5_ASAP7_75t_L g925 ( 
.A1(n_922),
.A2(n_916),
.B(n_912),
.C(n_913),
.Y(n_925)
);

NAND3xp33_ASAP7_75t_L g926 ( 
.A(n_921),
.B(n_919),
.C(n_910),
.Y(n_926)
);

NAND3xp33_ASAP7_75t_L g927 ( 
.A(n_923),
.B(n_911),
.C(n_844),
.Y(n_927)
);

OAI21xp33_ASAP7_75t_L g928 ( 
.A1(n_925),
.A2(n_920),
.B(n_914),
.Y(n_928)
);

OAI21xp33_ASAP7_75t_L g929 ( 
.A1(n_926),
.A2(n_915),
.B(n_823),
.Y(n_929)
);

NAND3xp33_ASAP7_75t_SL g930 ( 
.A(n_928),
.B(n_927),
.C(n_924),
.Y(n_930)
);

NOR2x1p5_ASAP7_75t_L g931 ( 
.A(n_929),
.B(n_838),
.Y(n_931)
);

OAI211xp5_ASAP7_75t_L g932 ( 
.A1(n_930),
.A2(n_794),
.B(n_800),
.C(n_820),
.Y(n_932)
);

AOI221xp5_ASAP7_75t_L g933 ( 
.A1(n_931),
.A2(n_821),
.B1(n_816),
.B2(n_818),
.C(n_813),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_932),
.B(n_901),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_933),
.A2(n_801),
.B(n_814),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_934),
.Y(n_936)
);

OA22x2_ASAP7_75t_L g937 ( 
.A1(n_935),
.A2(n_801),
.B1(n_822),
.B2(n_823),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_934),
.A2(n_863),
.B1(n_858),
.B2(n_829),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_936),
.A2(n_937),
.B1(n_938),
.B2(n_829),
.Y(n_939)
);

NAND3xp33_ASAP7_75t_L g940 ( 
.A(n_936),
.B(n_802),
.C(n_803),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_936),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_936),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_936),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_942),
.Y(n_944)
);

OAI22xp33_ASAP7_75t_L g945 ( 
.A1(n_941),
.A2(n_857),
.B1(n_828),
.B2(n_858),
.Y(n_945)
);

OAI211xp5_ASAP7_75t_L g946 ( 
.A1(n_943),
.A2(n_839),
.B(n_814),
.C(n_857),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_SL g947 ( 
.A1(n_940),
.A2(n_855),
.B1(n_828),
.B2(n_839),
.Y(n_947)
);

OAI21xp33_ASAP7_75t_SL g948 ( 
.A1(n_939),
.A2(n_819),
.B(n_803),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_942),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_942),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_950),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_944),
.A2(n_734),
.B(n_828),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_949),
.B(n_804),
.Y(n_953)
);

AOI21xp33_ASAP7_75t_L g954 ( 
.A1(n_948),
.A2(n_839),
.B(n_835),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_951),
.Y(n_955)
);

OA21x2_ASAP7_75t_L g956 ( 
.A1(n_953),
.A2(n_946),
.B(n_947),
.Y(n_956)
);

OR2x6_ASAP7_75t_L g957 ( 
.A(n_955),
.B(n_952),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_957),
.A2(n_954),
.B1(n_956),
.B2(n_945),
.Y(n_958)
);


endmodule