module fake_jpeg_13045_n_44 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_44);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_44;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

AO22x1_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_9),
.B1(n_15),
.B2(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_18),
.B(n_0),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_20),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_26),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_29),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_1),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_34),
.C(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_1),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_4),
.C(n_5),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_21),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_37),
.Y(n_39)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_12),
.C(n_13),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_14),
.C(n_16),
.Y(n_41)
);

NAND2xp33_ASAP7_75t_SL g42 ( 
.A(n_41),
.B(n_39),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);


endmodule