module fake_jpeg_18347_n_121 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_22),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_0),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_1),
.Y(n_76)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_58),
.Y(n_64)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_55),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_74),
.B1(n_75),
.B2(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_3),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_59),
.A2(n_43),
.B1(n_48),
.B2(n_52),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_51),
.B1(n_50),
.B2(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_1),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_72),
.B(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_83),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_2),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_67),
.Y(n_91)
);

NOR2xp67_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_2),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_54),
.B(n_21),
.C(n_23),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_86),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_39),
.B1(n_19),
.B2(n_20),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_17),
.C(n_37),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_24),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_5),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_3),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_4),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_100),
.Y(n_104)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_85),
.B1(n_7),
.B2(n_9),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_102),
.A2(n_107),
.B(n_95),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_98),
.A2(n_85),
.B1(n_10),
.B2(n_12),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_92),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

OAI322xp33_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_109),
.A3(n_110),
.B1(n_104),
.B2(n_106),
.C1(n_105),
.C2(n_102),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_28),
.C(n_13),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_112),
.A2(n_113),
.B(n_30),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_111),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_27),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_31),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_14),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_16),
.B(n_26),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_32),
.C(n_35),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_38),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_6),
.Y(n_121)
);


endmodule