module fake_jpeg_11499_n_644 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_644);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_644;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVxp33_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_12),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_14),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_33),
.A2(n_8),
.B1(n_17),
.B2(n_15),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_62),
.A2(n_56),
.B1(n_55),
.B2(n_29),
.Y(n_193)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_64),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_66),
.Y(n_149)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_68),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_69),
.Y(n_186)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_71),
.Y(n_174)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_74),
.Y(n_167)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_77),
.Y(n_189)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_80),
.Y(n_194)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_81),
.Y(n_161)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_82),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_25),
.B(n_7),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_115),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_84),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_85),
.Y(n_203)
);

BUFx24_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

CKINVDCx6p67_ASAP7_75t_R g214 ( 
.A(n_86),
.Y(n_214)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_87),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_40),
.B(n_7),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_89),
.B(n_120),
.Y(n_140)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g144 ( 
.A(n_90),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_91),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_93),
.Y(n_184)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_94),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_95),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_97),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_98),
.Y(n_195)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_99),
.Y(n_179)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_101),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_102),
.Y(n_211)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

INVx4_ASAP7_75t_SL g105 ( 
.A(n_20),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_122),
.Y(n_143)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_22),
.Y(n_109)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_53),
.B(n_7),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_130),
.B(n_28),
.C(n_50),
.Y(n_147)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_22),
.Y(n_112)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_113),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_41),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_32),
.B(n_8),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_26),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_41),
.Y(n_118)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_118),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_25),
.B(n_8),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_18),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_40),
.B(n_8),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_29),
.B(n_6),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_44),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_41),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_47),
.Y(n_124)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_22),
.Y(n_125)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_21),
.Y(n_126)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_126),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_21),
.Y(n_129)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

HAxp5_ASAP7_75t_SL g130 ( 
.A(n_19),
.B(n_0),
.CON(n_130),
.SN(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_21),
.B1(n_33),
.B2(n_45),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_131),
.A2(n_132),
.B1(n_152),
.B2(n_175),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_86),
.A2(n_45),
.B1(n_33),
.B2(n_52),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_110),
.A2(n_28),
.B1(n_19),
.B2(n_45),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_136),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_142),
.B(n_164),
.Y(n_228)
);

AO22x1_ASAP7_75t_L g278 ( 
.A1(n_147),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_148),
.B(n_157),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_99),
.A2(n_96),
.B1(n_95),
.B2(n_127),
.Y(n_152)
);

NAND3xp33_ASAP7_75t_L g286 ( 
.A(n_156),
.B(n_188),
.C(n_190),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_46),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_92),
.B(n_46),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_158),
.B(n_160),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_92),
.B(n_56),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_100),
.B(n_44),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_86),
.B(n_61),
.C(n_60),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_165),
.B(n_187),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_102),
.B(n_48),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_170),
.B(n_173),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_48),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_130),
.A2(n_52),
.B1(n_60),
.B2(n_32),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_72),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_106),
.B(n_59),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_111),
.B(n_59),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_105),
.B(n_38),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_192),
.B(n_51),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_193),
.A2(n_212),
.B1(n_213),
.B2(n_35),
.Y(n_246)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_128),
.Y(n_196)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_73),
.B(n_37),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_202),
.B(n_31),
.Y(n_258)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_112),
.Y(n_204)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_93),
.A2(n_35),
.B1(n_38),
.B2(n_61),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_124),
.A2(n_55),
.B1(n_37),
.B2(n_26),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_143),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_218),
.Y(n_349)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_219),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_131),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_220)
);

AOI22x1_ASAP7_75t_L g307 ( 
.A1(n_220),
.A2(n_133),
.B1(n_199),
.B2(n_171),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_162),
.Y(n_221)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_221),
.Y(n_302)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_223),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_140),
.B(n_58),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_225),
.B(n_231),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_151),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_227),
.B(n_255),
.Y(n_315)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_229),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_134),
.B(n_58),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_232),
.Y(n_313)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_175),
.A2(n_69),
.B1(n_113),
.B2(n_101),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_234),
.A2(n_252),
.B1(n_210),
.B2(n_217),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_162),
.Y(n_235)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_235),
.Y(n_323)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_159),
.Y(n_236)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_236),
.Y(n_306)
);

INVx11_ASAP7_75t_L g237 ( 
.A(n_144),
.Y(n_237)
);

INVx11_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_166),
.Y(n_238)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_238),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_143),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_239),
.Y(n_309)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_240),
.Y(n_299)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_144),
.Y(n_241)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_241),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_192),
.A2(n_114),
.B1(n_77),
.B2(n_98),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_242),
.A2(n_248),
.B1(n_271),
.B2(n_281),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_162),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_243),
.B(n_246),
.Y(n_320)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_135),
.Y(n_244)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_244),
.Y(n_329)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_178),
.Y(n_245)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_245),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_138),
.B(n_23),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_247),
.B(n_273),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_141),
.A2(n_84),
.B1(n_91),
.B2(n_85),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_146),
.A2(n_104),
.B1(n_51),
.B2(n_31),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_250),
.Y(n_297)
);

INVx13_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_251),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_132),
.A2(n_88),
.B1(n_74),
.B2(n_90),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_181),
.Y(n_253)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_253),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_189),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_254),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_151),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_155),
.Y(n_256)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_256),
.Y(n_331)
);

OAI21xp33_ASAP7_75t_L g295 ( 
.A1(n_257),
.A2(n_269),
.B(n_272),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_258),
.B(n_249),
.Y(n_304)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_154),
.Y(n_259)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_259),
.Y(n_348)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_197),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_260),
.Y(n_352)
);

OA22x2_ASAP7_75t_L g261 ( 
.A1(n_207),
.A2(n_30),
.B1(n_23),
.B2(n_2),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_SL g305 ( 
.A1(n_261),
.A2(n_217),
.B(n_210),
.C(n_167),
.Y(n_305)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_139),
.Y(n_263)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_263),
.Y(n_335)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_183),
.Y(n_264)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_264),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_197),
.Y(n_266)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_266),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_184),
.Y(n_267)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_267),
.Y(n_338)
);

INVx8_ASAP7_75t_L g268 ( 
.A(n_145),
.Y(n_268)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_268),
.Y(n_350)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_182),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_169),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_270),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_L g271 ( 
.A1(n_212),
.A2(n_30),
.B1(n_9),
.B2(n_11),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_161),
.B(n_0),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_185),
.B(n_0),
.Y(n_273)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_214),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_274),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_169),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_275),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_191),
.B(n_1),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_276),
.B(n_288),
.Y(n_312)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_183),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_277),
.B(n_4),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_292),
.Y(n_294)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_211),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_279),
.B(n_282),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_176),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_280),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_150),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_155),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_180),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_283),
.B(n_285),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_194),
.A2(n_5),
.B1(n_6),
.B2(n_11),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_284),
.A2(n_287),
.B1(n_293),
.B2(n_153),
.Y(n_345)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_145),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_201),
.A2(n_5),
.B1(n_6),
.B2(n_17),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_174),
.B(n_1),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_180),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_289),
.B(n_290),
.Y(n_346)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_176),
.Y(n_290)
);

INVx11_ASAP7_75t_L g292 ( 
.A(n_214),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_133),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_293)
);

OAI22x1_ASAP7_75t_SL g301 ( 
.A1(n_226),
.A2(n_177),
.B1(n_163),
.B2(n_168),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_301),
.A2(n_307),
.B1(n_308),
.B2(n_314),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_304),
.B(n_310),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_345),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_265),
.A2(n_199),
.B1(n_171),
.B2(n_172),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_225),
.B(n_198),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_218),
.A2(n_209),
.B1(n_205),
.B2(n_172),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_319),
.A2(n_333),
.B1(n_292),
.B2(n_237),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_273),
.B(n_209),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_321),
.B(n_328),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_L g327 ( 
.A1(n_220),
.A2(n_208),
.B1(n_195),
.B2(n_205),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_327),
.A2(n_334),
.B1(n_267),
.B2(n_268),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_247),
.B(n_150),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_230),
.A2(n_149),
.B1(n_186),
.B2(n_203),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_L g334 ( 
.A1(n_271),
.A2(n_149),
.B1(n_186),
.B2(n_203),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_239),
.A2(n_137),
.B(n_153),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_336),
.A2(n_351),
.B(n_267),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_291),
.B(n_1),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_347),
.B(n_241),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_288),
.A2(n_1),
.B(n_4),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_353),
.Y(n_358)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_299),
.Y(n_355)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_355),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_328),
.A2(n_262),
.B1(n_276),
.B2(n_228),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_356),
.A2(n_357),
.B1(n_371),
.B2(n_382),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_311),
.A2(n_231),
.B1(n_278),
.B2(n_261),
.Y(n_357)
);

A2O1A1Ixp33_ASAP7_75t_L g360 ( 
.A1(n_294),
.A2(n_257),
.B(n_286),
.C(n_272),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_360),
.B(n_362),
.Y(n_404)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_338),
.Y(n_361)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_361),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_311),
.B(n_272),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_300),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_366),
.Y(n_403)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_299),
.Y(n_365)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_365),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_300),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_367),
.B(n_380),
.Y(n_401)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_315),
.Y(n_368)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_368),
.Y(n_417)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_369),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_321),
.B(n_288),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_370),
.B(n_377),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_294),
.A2(n_261),
.B1(n_263),
.B2(n_244),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_348),
.Y(n_372)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_372),
.Y(n_420)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_348),
.Y(n_373)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_373),
.Y(n_422)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_303),
.Y(n_375)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_375),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_349),
.B(n_312),
.C(n_309),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_376),
.B(n_379),
.C(n_398),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_312),
.B(n_257),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_378),
.A2(n_297),
.B1(n_301),
.B2(n_334),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_295),
.B(n_233),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_269),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_346),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_381),
.B(n_385),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_320),
.A2(n_261),
.B1(n_223),
.B2(n_229),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g383 ( 
.A(n_318),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_383),
.Y(n_405)
);

AO21x2_ASAP7_75t_SL g384 ( 
.A1(n_305),
.A2(n_274),
.B(n_251),
.Y(n_384)
);

OA22x2_ASAP7_75t_L g431 ( 
.A1(n_384),
.A2(n_331),
.B1(n_316),
.B2(n_343),
.Y(n_431)
);

A2O1A1Ixp33_ASAP7_75t_L g385 ( 
.A1(n_310),
.A2(n_296),
.B(n_320),
.C(n_349),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_386),
.A2(n_393),
.B1(n_298),
.B2(n_313),
.Y(n_424)
);

O2A1O1Ixp33_ASAP7_75t_L g387 ( 
.A1(n_297),
.A2(n_275),
.B(n_224),
.C(n_222),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_387),
.A2(n_392),
.B(n_396),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_325),
.B(n_240),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_388),
.B(n_391),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_322),
.Y(n_389)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_389),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_390),
.A2(n_340),
.B(n_335),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_317),
.B(n_264),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_296),
.B(n_277),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_320),
.A2(n_232),
.B1(n_260),
.B2(n_219),
.Y(n_393)
);

INVx3_ASAP7_75t_SL g394 ( 
.A(n_322),
.Y(n_394)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_394),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_308),
.A2(n_282),
.B1(n_285),
.B2(n_283),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_395),
.A2(n_393),
.B1(n_364),
.B2(n_366),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_306),
.B(n_256),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_397),
.Y(n_418)
);

MAJx2_ASAP7_75t_L g398 ( 
.A(n_333),
.B(n_243),
.C(n_289),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_298),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_399),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_336),
.B(n_279),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_390),
.C(n_379),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_409),
.A2(n_410),
.B1(n_415),
.B2(n_382),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_374),
.A2(n_307),
.B1(n_330),
.B2(n_327),
.Y(n_410)
);

INVxp33_ASAP7_75t_L g460 ( 
.A(n_411),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_357),
.B(n_351),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_412),
.B(n_359),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_406),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_374),
.A2(n_307),
.B1(n_341),
.B2(n_337),
.Y(n_415)
);

OA21x2_ASAP7_75t_SL g416 ( 
.A1(n_362),
.A2(n_332),
.B(n_342),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_416),
.B(n_355),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_363),
.A2(n_324),
.B(n_316),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_419),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_400),
.A2(n_302),
.B(n_323),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_421),
.A2(n_426),
.B(n_385),
.Y(n_453)
);

OAI22xp33_ASAP7_75t_SL g444 ( 
.A1(n_424),
.A2(n_378),
.B1(n_373),
.B2(n_372),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_376),
.B(n_329),
.C(n_335),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_427),
.B(n_438),
.C(n_391),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_363),
.A2(n_350),
.B1(n_302),
.B2(n_323),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_430),
.A2(n_384),
.B(n_380),
.Y(n_449)
);

AO22x2_ASAP7_75t_L g456 ( 
.A1(n_431),
.A2(n_437),
.B1(n_384),
.B2(n_386),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_363),
.A2(n_326),
.B1(n_344),
.B2(n_352),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_436),
.A2(n_384),
.B1(n_394),
.B2(n_397),
.Y(n_454)
);

OA22x2_ASAP7_75t_L g437 ( 
.A1(n_384),
.A2(n_331),
.B1(n_329),
.B2(n_303),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_354),
.B(n_343),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_403),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_440),
.B(n_446),
.Y(n_480)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_403),
.Y(n_441)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_441),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_442),
.A2(n_451),
.B1(n_437),
.B2(n_431),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_444),
.A2(n_454),
.B1(n_463),
.B2(n_408),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_445),
.B(n_455),
.C(n_457),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_425),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_402),
.Y(n_447)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_447),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_367),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_448),
.B(n_450),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_449),
.A2(n_453),
.B(n_458),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_381),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_415),
.A2(n_410),
.B1(n_409),
.B2(n_419),
.Y(n_451)
);

INVxp33_ASAP7_75t_SL g452 ( 
.A(n_425),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_452),
.B(n_466),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_456),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_406),
.B(n_392),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_413),
.A2(n_358),
.B(n_368),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_354),
.Y(n_459)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_459),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_426),
.A2(n_387),
.B(n_360),
.Y(n_461)
);

AO21x1_ASAP7_75t_L g502 ( 
.A1(n_461),
.A2(n_468),
.B(n_405),
.Y(n_502)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_402),
.Y(n_462)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_462),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_423),
.A2(n_359),
.B1(n_370),
.B2(n_371),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_414),
.Y(n_464)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_464),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_408),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_465),
.B(n_474),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_433),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_404),
.B(n_377),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_467),
.B(n_473),
.C(n_416),
.Y(n_499)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_414),
.Y(n_469)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_469),
.Y(n_486)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_420),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_471),
.Y(n_488)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_420),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_417),
.B(n_356),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_472),
.B(n_428),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_404),
.B(n_396),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_422),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_475),
.B(n_438),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_451),
.A2(n_423),
.B1(n_412),
.B2(n_430),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_476),
.A2(n_479),
.B1(n_495),
.B2(n_500),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_477),
.B(n_499),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_427),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_478),
.B(n_481),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_442),
.A2(n_412),
.B1(n_436),
.B2(n_411),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_457),
.B(n_432),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_432),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_483),
.B(n_505),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_440),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_487),
.B(n_497),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_492),
.A2(n_496),
.B1(n_498),
.B2(n_461),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_465),
.A2(n_424),
.B1(n_421),
.B2(n_417),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_463),
.A2(n_401),
.B1(n_437),
.B2(n_431),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_466),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_454),
.A2(n_401),
.B1(n_437),
.B2(n_431),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_502),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_453),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_503),
.B(n_509),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_446),
.A2(n_422),
.B1(n_431),
.B2(n_437),
.Y(n_504)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_504),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_473),
.B(n_365),
.Y(n_505)
);

A2O1A1Ixp33_ASAP7_75t_L g506 ( 
.A1(n_449),
.A2(n_428),
.B(n_398),
.C(n_439),
.Y(n_506)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_506),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_476),
.A2(n_443),
.B1(n_441),
.B2(n_460),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_510),
.A2(n_514),
.B1(n_492),
.B2(n_496),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_SL g511 ( 
.A(n_491),
.B(n_443),
.Y(n_511)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_511),
.Y(n_550)
);

XOR2x2_ASAP7_75t_L g513 ( 
.A(n_491),
.B(n_468),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_513),
.B(n_535),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_479),
.A2(n_445),
.B1(n_472),
.B2(n_475),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_515),
.A2(n_516),
.B1(n_495),
.B2(n_488),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_490),
.A2(n_474),
.B1(n_471),
.B2(n_470),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_478),
.B(n_458),
.C(n_459),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_520),
.B(n_524),
.C(n_527),
.Y(n_555)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_480),
.Y(n_523)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_523),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_484),
.B(n_469),
.C(n_464),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_SL g525 ( 
.A(n_482),
.B(n_456),
.Y(n_525)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_525),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_484),
.B(n_462),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_526),
.B(n_531),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_481),
.B(n_447),
.C(n_439),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_499),
.B(n_407),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_477),
.B(n_407),
.C(n_433),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_532),
.B(n_536),
.C(n_538),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_483),
.B(n_398),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_533),
.B(n_534),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_505),
.B(n_375),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_480),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_489),
.B(n_418),
.C(n_361),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_502),
.B(n_456),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_537),
.B(n_507),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_489),
.B(n_418),
.C(n_369),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_482),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_539),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_SL g575 ( 
.A(n_540),
.B(n_537),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_528),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_542),
.B(n_547),
.Y(n_579)
);

AOI21xp33_ASAP7_75t_SL g543 ( 
.A1(n_513),
.A2(n_508),
.B(n_506),
.Y(n_543)
);

BUFx24_ASAP7_75t_SL g568 ( 
.A(n_543),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_536),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_544),
.B(n_546),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_538),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_512),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_551),
.B(n_558),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_529),
.A2(n_501),
.B1(n_498),
.B2(n_507),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_552),
.Y(n_584)
);

NOR3xp33_ASAP7_75t_SL g553 ( 
.A(n_522),
.B(n_488),
.C(n_494),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_553),
.A2(n_554),
.B1(n_530),
.B2(n_514),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_526),
.B(n_494),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_524),
.B(n_486),
.C(n_493),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_559),
.B(n_561),
.C(n_563),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_518),
.B(n_486),
.C(n_493),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_529),
.A2(n_485),
.B1(n_456),
.B2(n_434),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_SL g576 ( 
.A1(n_562),
.A2(n_434),
.B1(n_429),
.B2(n_394),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_518),
.B(n_485),
.C(n_418),
.Y(n_563)
);

NOR2x1p5_ASAP7_75t_L g564 ( 
.A(n_533),
.B(n_456),
.Y(n_564)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_564),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_541),
.B(n_531),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_569),
.B(n_575),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_548),
.A2(n_530),
.B(n_510),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_570),
.A2(n_580),
.B(n_582),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_553),
.B(n_517),
.Y(n_571)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_571),
.Y(n_592)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_572),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_555),
.B(n_527),
.C(n_520),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_573),
.B(n_577),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_545),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_574),
.B(n_581),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_576),
.A2(n_389),
.B1(n_344),
.B2(n_326),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_555),
.B(n_532),
.C(n_519),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_SL g578 ( 
.A1(n_560),
.A2(n_534),
.B(n_521),
.Y(n_578)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_578),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_550),
.A2(n_519),
.B(n_521),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_559),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_551),
.A2(n_429),
.B(n_399),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_557),
.Y(n_583)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_583),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_571),
.A2(n_546),
.B1(n_544),
.B2(n_564),
.Y(n_587)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_587),
.Y(n_604)
);

CKINVDCx14_ASAP7_75t_R g589 ( 
.A(n_579),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_589),
.B(n_566),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_567),
.B(n_561),
.C(n_556),
.Y(n_590)
);

NOR2xp67_ASAP7_75t_SL g614 ( 
.A(n_590),
.B(n_591),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_567),
.B(n_573),
.C(n_577),
.Y(n_591)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_574),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_598),
.A2(n_603),
.B1(n_584),
.B2(n_389),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_565),
.B(n_558),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_599),
.B(n_600),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_569),
.B(n_541),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_565),
.B(n_556),
.C(n_563),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_601),
.B(n_549),
.C(n_578),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_570),
.A2(n_564),
.B(n_549),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_602),
.A2(n_582),
.B(n_585),
.Y(n_605)
);

AOI21x1_ASAP7_75t_L g625 ( 
.A1(n_605),
.A2(n_606),
.B(n_593),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_592),
.A2(n_585),
.B(n_575),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_SL g607 ( 
.A(n_586),
.B(n_568),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_607),
.B(n_616),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_609),
.B(n_610),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_601),
.B(n_566),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_611),
.B(n_612),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_590),
.B(n_580),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_613),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_591),
.B(n_352),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_615),
.B(n_617),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_594),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_595),
.B(n_254),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_608),
.B(n_595),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_618),
.B(n_623),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_610),
.B(n_594),
.C(n_592),
.Y(n_623)
);

NOR2x1_ASAP7_75t_L g624 ( 
.A(n_616),
.B(n_596),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_624),
.A2(n_606),
.B(n_605),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_L g630 ( 
.A1(n_625),
.A2(n_593),
.B(n_602),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_612),
.B(n_600),
.Y(n_627)
);

XOR2xp5_ASAP7_75t_L g629 ( 
.A(n_627),
.B(n_613),
.Y(n_629)
);

OAI321xp33_ASAP7_75t_L g628 ( 
.A1(n_619),
.A2(n_604),
.A3(n_598),
.B1(n_597),
.B2(n_596),
.C(n_587),
.Y(n_628)
);

AOI31xp33_ASAP7_75t_L g635 ( 
.A1(n_628),
.A2(n_634),
.A3(n_620),
.B(n_621),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_629),
.B(n_620),
.C(n_608),
.Y(n_636)
);

AOI21xp33_ASAP7_75t_L g637 ( 
.A1(n_630),
.A2(n_588),
.B(n_597),
.Y(n_637)
);

AO21x1_ASAP7_75t_L g631 ( 
.A1(n_622),
.A2(n_614),
.B(n_599),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_631),
.A2(n_633),
.B(n_588),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_624),
.B(n_618),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g640 ( 
.A1(n_635),
.A2(n_638),
.B(n_221),
.Y(n_640)
);

A2O1A1O1Ixp25_ASAP7_75t_L g639 ( 
.A1(n_636),
.A2(n_637),
.B(n_632),
.C(n_626),
.D(n_603),
.Y(n_639)
);

BUFx24_ASAP7_75t_SL g641 ( 
.A(n_639),
.Y(n_641)
);

NAND3xp33_ASAP7_75t_L g642 ( 
.A(n_641),
.B(n_640),
.C(n_235),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_642),
.B(n_313),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_643),
.B(n_266),
.Y(n_644)
);


endmodule