module fake_jpeg_13970_n_407 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_407);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_407;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_15),
.B(n_3),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_48),
.Y(n_96)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_49),
.Y(n_79)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_60),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_22),
.Y(n_52)
);

INVx5_ASAP7_75t_SL g110 ( 
.A(n_52),
.Y(n_110)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_14),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_73),
.Y(n_100)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_56),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_1),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_18),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_62),
.Y(n_111)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_63),
.Y(n_82)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_36),
.Y(n_104)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_30),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_78),
.B(n_98),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_40),
.A2(n_31),
.B1(n_36),
.B2(n_26),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_87),
.A2(n_108),
.B1(n_26),
.B2(n_68),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_40),
.B(n_29),
.C(n_20),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_21),
.C(n_23),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_52),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_31),
.B1(n_35),
.B2(n_33),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_101),
.A2(n_28),
.B1(n_19),
.B2(n_70),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_104),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_35),
.B(n_21),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_19),
.B(n_24),
.C(n_27),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_36),
.B1(n_26),
.B2(n_27),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_41),
.B(n_33),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_32),
.Y(n_125)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_115),
.Y(n_170)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_116),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_24),
.B(n_27),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_108),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_110),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_125),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_119),
.B(n_138),
.Y(n_193)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_110),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_122),
.Y(n_167)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_123),
.Y(n_191)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_23),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_129),
.Y(n_158)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_134),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_32),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_99),
.A2(n_47),
.B1(n_58),
.B2(n_26),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_130),
.A2(n_139),
.B(n_79),
.Y(n_172)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_132),
.A2(n_150),
.B1(n_151),
.B2(n_153),
.Y(n_166)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_133),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_81),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_137),
.Y(n_175)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_136),
.Y(n_187)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_105),
.A2(n_19),
.B1(n_24),
.B2(n_26),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_142),
.Y(n_192)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_149),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_148),
.A2(n_96),
.B1(n_87),
.B2(n_112),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_82),
.B(n_28),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_96),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_90),
.A2(n_65),
.B1(n_61),
.B2(n_59),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_46),
.B1(n_57),
.B2(n_45),
.Y(n_162)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_155),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_159),
.B(n_5),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_117),
.B(n_86),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_169),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_162),
.A2(n_171),
.B1(n_144),
.B2(n_124),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_141),
.B1(n_120),
.B2(n_150),
.Y(n_200)
);

NAND2xp33_ASAP7_75t_SL g165 ( 
.A(n_122),
.B(n_82),
.Y(n_165)
);

NAND2xp33_ASAP7_75t_SL g231 ( 
.A(n_165),
.B(n_181),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_125),
.B(n_103),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_112),
.B1(n_103),
.B2(n_92),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_2),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_79),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_138),
.C(n_137),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_129),
.B(n_107),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_185),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_147),
.A2(n_114),
.B1(n_109),
.B2(n_92),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_109),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_1),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_4),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_119),
.B(n_58),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_188),
.B(n_48),
.Y(n_215)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_194),
.Y(n_233)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_195),
.Y(n_240)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_197),
.Y(n_261)
);

OA21x2_ASAP7_75t_L g198 ( 
.A1(n_185),
.A2(n_130),
.B(n_133),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_121),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_199),
.B(n_221),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_208),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g254 ( 
.A(n_201),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_146),
.B(n_145),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_202),
.A2(n_212),
.B(n_216),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_158),
.A2(n_131),
.B1(n_127),
.B2(n_143),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_203),
.A2(n_223),
.B1(n_225),
.B2(n_227),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_183),
.A2(n_152),
.B1(n_155),
.B2(n_136),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_158),
.A2(n_153),
.B1(n_151),
.B2(n_142),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_219),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_159),
.A2(n_34),
.B(n_85),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_165),
.B(n_175),
.Y(n_234)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_213),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_224),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_172),
.B(n_2),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_170),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_34),
.C(n_5),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_220)
);

INVxp33_ASAP7_75t_SL g266 ( 
.A(n_220),
.Y(n_266)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_229),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_174),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_223)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_173),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_170),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_160),
.B(n_7),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_226),
.B(n_179),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_174),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_188),
.B1(n_186),
.B2(n_178),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_230),
.B1(n_167),
.B2(n_166),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_8),
.C(n_9),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_169),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_234),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_203),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_245),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_247),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_204),
.A2(n_175),
.B(n_173),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_239),
.A2(n_253),
.B(n_259),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_242),
.A2(n_209),
.B1(n_197),
.B2(n_195),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_214),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_167),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_230),
.Y(n_272)
);

AO22x1_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_170),
.B1(n_176),
.B2(n_156),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_248),
.B(n_256),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_204),
.A2(n_192),
.B(n_191),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_196),
.B(n_218),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_265),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_196),
.B(n_192),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_191),
.B(n_190),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_202),
.B(n_179),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_177),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_212),
.A2(n_191),
.B(n_187),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_216),
.B(n_212),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_210),
.B(n_157),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_246),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_267),
.B(n_272),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_200),
.B1(n_228),
.B2(n_211),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_268),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_269),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_222),
.C(n_219),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_290),
.C(n_260),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_213),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_275),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_246),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_281),
.Y(n_314)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_233),
.Y(n_277)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_278),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_254),
.B1(n_236),
.B2(n_265),
.Y(n_280)
);

INVxp33_ASAP7_75t_SL g281 ( 
.A(n_232),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_249),
.A2(n_198),
.B1(n_227),
.B2(n_223),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_259),
.A2(n_198),
.B1(n_229),
.B2(n_216),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_285),
.A2(n_292),
.B1(n_264),
.B2(n_250),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_243),
.B(n_157),
.Y(n_286)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_286),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_247),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_288),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_247),
.Y(n_288)
);

INVxp33_ASAP7_75t_L g289 ( 
.A(n_239),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_235),
.B(n_179),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_255),
.A2(n_234),
.B1(n_242),
.B2(n_251),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_291),
.A2(n_258),
.B1(n_241),
.B2(n_250),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_243),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_293),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_253),
.Y(n_294)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_294),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_260),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_296),
.B(n_313),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_287),
.A2(n_251),
.B1(n_252),
.B2(n_266),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_300),
.A2(n_268),
.B1(n_282),
.B2(n_258),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_318),
.C(n_274),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_303),
.Y(n_326)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_285),
.A2(n_238),
.B1(n_252),
.B2(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_308),
.Y(n_334)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_309),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_270),
.B(n_264),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_315),
.A2(n_288),
.B1(n_294),
.B2(n_271),
.Y(n_323)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_293),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_279),
.B(n_257),
.C(n_261),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_279),
.B(n_241),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_319),
.B(n_291),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_280),
.A2(n_258),
.B1(n_261),
.B2(n_240),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_320),
.A2(n_284),
.B1(n_276),
.B2(n_272),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_322),
.B(n_335),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_323),
.A2(n_327),
.B1(n_333),
.B2(n_341),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_271),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_324),
.B(n_330),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_301),
.A2(n_295),
.B1(n_272),
.B2(n_267),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_314),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_311),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_302),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_331),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_275),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_295),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_338),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_284),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_301),
.B(n_283),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_298),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_337),
.A2(n_334),
.B1(n_326),
.B2(n_320),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_314),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_339),
.B(n_316),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_315),
.A2(n_278),
.B1(n_277),
.B2(n_269),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_299),
.C(n_304),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_344),
.B(n_348),
.Y(n_365)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_345),
.Y(n_358)
);

AOI21x1_ASAP7_75t_L g347 ( 
.A1(n_340),
.A2(n_304),
.B(n_312),
.Y(n_347)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_347),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_330),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_331),
.B(n_319),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_297),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_299),
.C(n_307),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_350),
.B(n_354),
.C(n_344),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_351),
.B(n_321),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_353),
.A2(n_341),
.B1(n_333),
.B2(n_336),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_300),
.C(n_306),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_355),
.B(n_357),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_305),
.Y(n_357)
);

NAND2x1p5_ASAP7_75t_L g359 ( 
.A(n_354),
.B(n_324),
.Y(n_359)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_359),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_362),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_337),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_363),
.B(n_350),
.Y(n_373)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_342),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_364),
.B(n_370),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_369),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_355),
.A2(n_305),
.B1(n_322),
.B2(n_310),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_368),
.B(n_357),
.Y(n_371)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_356),
.Y(n_370)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_371),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_373),
.A2(n_367),
.B1(n_368),
.B2(n_244),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_366),
.B(n_346),
.C(n_349),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_375),
.B(n_378),
.Y(n_386)
);

A2O1A1Ixp33_ASAP7_75t_SL g377 ( 
.A1(n_361),
.A2(n_352),
.B(n_346),
.C(n_257),
.Y(n_377)
);

AO21x1_ASAP7_75t_L g389 ( 
.A1(n_377),
.A2(n_10),
.B(n_12),
.Y(n_389)
);

BUFx24_ASAP7_75t_SL g378 ( 
.A(n_358),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_369),
.B(n_352),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_379),
.B(n_9),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_359),
.A2(n_240),
.B1(n_244),
.B2(n_168),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_381),
.A2(n_244),
.B1(n_168),
.B2(n_367),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_374),
.A2(n_365),
.B(n_360),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_382),
.A2(n_373),
.B(n_372),
.Y(n_391)
);

AND2x2_ASAP7_75t_SL g392 ( 
.A(n_384),
.B(n_387),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_389),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_380),
.A2(n_177),
.B1(n_176),
.B2(n_156),
.Y(n_387)
);

OR2x6_ASAP7_75t_SL g393 ( 
.A(n_388),
.B(n_390),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_376),
.A2(n_10),
.B(n_12),
.Y(n_390)
);

AO21x2_ASAP7_75t_L g400 ( 
.A1(n_391),
.A2(n_13),
.B(n_14),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_386),
.B(n_377),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_395),
.B(n_396),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_383),
.B(n_10),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_391),
.A2(n_382),
.B1(n_389),
.B2(n_390),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_397),
.B(n_398),
.C(n_400),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_394),
.B(n_388),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_399),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_402),
.Y(n_403)
);

AOI21x1_ASAP7_75t_L g404 ( 
.A1(n_403),
.A2(n_401),
.B(n_393),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_404),
.A2(n_392),
.B(n_13),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_405),
.B(n_13),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_406),
.A2(n_13),
.B(n_14),
.Y(n_407)
);


endmodule