module fake_netlist_6_4740_n_1825 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1825);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1825;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g174 ( 
.A(n_0),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_20),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_76),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_99),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_161),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_35),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_43),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_43),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_55),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_38),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_108),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_84),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_171),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_104),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_8),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_29),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_28),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_83),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_117),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_51),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_48),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_128),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_131),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_60),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_8),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_127),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_88),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_39),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_38),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_63),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_72),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_46),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_152),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_41),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_63),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_28),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_162),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_67),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_4),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_100),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_95),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_122),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_69),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_86),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_39),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_64),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_155),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_52),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_167),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_56),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_133),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_23),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_59),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_7),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_21),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_124),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_123),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_37),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_154),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_129),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_52),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_12),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_5),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_98),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_64),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_138),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_48),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_106),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_27),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_30),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_60),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_147),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_26),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_148),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_10),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_25),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_21),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_24),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_102),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_130),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_170),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_3),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_6),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_56),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_25),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_80),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_49),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_134),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_58),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_149),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_135),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_101),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_44),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_0),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_150),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_34),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_73),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_94),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_13),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_16),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_109),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_136),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_59),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_23),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_1),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_3),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_137),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_165),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_55),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_26),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_156),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_1),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_31),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_114),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_87),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_81),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_31),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_85),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_91),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_139),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_118),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_45),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_160),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_35),
.Y(n_303)
);

INVxp33_ASAP7_75t_L g304 ( 
.A(n_70),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_29),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_53),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_6),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_15),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_145),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_33),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_5),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_75),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_19),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_46),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_166),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_32),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_22),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_41),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_153),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_27),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_18),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_36),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_142),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_163),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_18),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_47),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_82),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_19),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_34),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_44),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_140),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_132),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_169),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_93),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_47),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_74),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_96),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_16),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_10),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_115),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_9),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_178),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_189),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_190),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_246),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_191),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_182),
.B(n_2),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_246),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_233),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_197),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_246),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_200),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_202),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_205),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_206),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_233),
.B(n_7),
.Y(n_356)
);

NOR2xp67_ASAP7_75t_L g357 ( 
.A(n_175),
.B(n_9),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_182),
.B(n_11),
.Y(n_358)
);

BUFx6f_ASAP7_75t_SL g359 ( 
.A(n_315),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_243),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_246),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_246),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_341),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_246),
.Y(n_364)
);

BUFx10_ASAP7_75t_L g365 ( 
.A(n_188),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_217),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_301),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_216),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_222),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_301),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_220),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_301),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_223),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_225),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_213),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_303),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_226),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_176),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_176),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_228),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_243),
.B(n_11),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_301),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_337),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_301),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_195),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_235),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_236),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_195),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_211),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_211),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_258),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_333),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_325),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_325),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_174),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_239),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_181),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_174),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_180),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_245),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_341),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_180),
.Y(n_402)
);

BUFx2_ASAP7_75t_SL g403 ( 
.A(n_188),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_337),
.B(n_12),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_183),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_186),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_247),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_181),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_299),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_186),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_192),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_251),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_224),
.B(n_13),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_253),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_177),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_260),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_192),
.Y(n_417)
);

BUFx2_ASAP7_75t_SL g418 ( 
.A(n_212),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_194),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_265),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_303),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_194),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_207),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_207),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_209),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_267),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_269),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_209),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_409),
.B(n_212),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_370),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_403),
.B(n_304),
.Y(n_431)
);

AND2x6_ASAP7_75t_L g432 ( 
.A(n_356),
.B(n_297),
.Y(n_432)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_370),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_345),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_345),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_378),
.B(n_299),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_348),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_348),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_351),
.Y(n_439)
);

INVx5_ASAP7_75t_L g440 ( 
.A(n_365),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_351),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_361),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_361),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_362),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_362),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_364),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_364),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_367),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_403),
.B(n_238),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_367),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_372),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_372),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_382),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_347),
.B(n_315),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_382),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_358),
.B(n_315),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_384),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_384),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_379),
.B(n_328),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_418),
.B(n_340),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_385),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_415),
.B(n_328),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_356),
.B(n_177),
.Y(n_464)
);

OA21x2_ASAP7_75t_L g465 ( 
.A1(n_388),
.A2(n_231),
.B(n_214),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_418),
.B(n_395),
.Y(n_466)
);

OA21x2_ASAP7_75t_L g467 ( 
.A1(n_388),
.A2(n_231),
.B(n_214),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_381),
.A2(n_244),
.B1(n_266),
.B2(n_273),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_389),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_376),
.B(n_184),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_376),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_389),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_390),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_390),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_421),
.B(n_184),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_393),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_375),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_393),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_421),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_394),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_395),
.B(n_193),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_405),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_394),
.Y(n_483)
);

NAND2xp33_ASAP7_75t_R g484 ( 
.A(n_404),
.B(n_185),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_398),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_398),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_349),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_399),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_399),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_406),
.B(n_193),
.Y(n_490)
);

NAND2x1_ASAP7_75t_L g491 ( 
.A(n_406),
.B(n_297),
.Y(n_491)
);

NAND3xp33_ASAP7_75t_L g492 ( 
.A(n_402),
.B(n_240),
.C(n_234),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_410),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_410),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_411),
.B(n_196),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_411),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_417),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_360),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_428),
.Y(n_499)
);

INVx6_ASAP7_75t_L g500 ( 
.A(n_365),
.Y(n_500)
);

AND2x6_ASAP7_75t_L g501 ( 
.A(n_417),
.B(n_297),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_414),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_419),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_383),
.B(n_196),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_419),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_432),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_465),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_431),
.B(n_342),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_433),
.Y(n_509)
);

AND2x6_ASAP7_75t_L g510 ( 
.A(n_464),
.B(n_201),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_454),
.B(n_456),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_465),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_435),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_433),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_435),
.Y(n_515)
);

NAND3xp33_ASAP7_75t_L g516 ( 
.A(n_431),
.B(n_374),
.C(n_344),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_435),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_465),
.Y(n_518)
);

OR2x6_ASAP7_75t_L g519 ( 
.A(n_498),
.B(n_357),
.Y(n_519)
);

INVxp33_ASAP7_75t_L g520 ( 
.A(n_471),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_435),
.Y(n_521)
);

INVx5_ASAP7_75t_L g522 ( 
.A(n_432),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_439),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_449),
.B(n_343),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_477),
.Y(n_525)
);

AO21x2_ASAP7_75t_L g526 ( 
.A1(n_454),
.A2(n_210),
.B(n_201),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_449),
.B(n_346),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_502),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_439),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_439),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_439),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_456),
.B(n_350),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_464),
.A2(n_229),
.B1(n_339),
.B2(n_313),
.Y(n_533)
);

BUFx4f_ASAP7_75t_L g534 ( 
.A(n_465),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_L g535 ( 
.A(n_432),
.B(n_297),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_461),
.B(n_352),
.Y(n_536)
);

AND2x2_ASAP7_75t_SL g537 ( 
.A(n_464),
.B(n_210),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_441),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_464),
.A2(n_229),
.B1(n_313),
.B2(n_339),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_465),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_502),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_464),
.A2(n_504),
.B1(n_432),
.B2(n_475),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_441),
.Y(n_543)
);

INVx8_ASAP7_75t_L g544 ( 
.A(n_432),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_477),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_465),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_464),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_461),
.B(n_353),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_498),
.B(n_354),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_467),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_467),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_471),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_467),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_441),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_440),
.B(n_355),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_467),
.Y(n_556)
);

AND2x6_ASAP7_75t_L g557 ( 
.A(n_481),
.B(n_219),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_SL g558 ( 
.A(n_484),
.B(n_504),
.Y(n_558)
);

BUFx10_ASAP7_75t_L g559 ( 
.A(n_500),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_479),
.B(n_368),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_479),
.B(n_371),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_429),
.B(n_373),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_441),
.Y(n_563)
);

AND2x6_ASAP7_75t_L g564 ( 
.A(n_481),
.B(n_219),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_442),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_442),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_489),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_429),
.B(n_377),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_467),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_466),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_442),
.Y(n_571)
);

AO22x2_ASAP7_75t_L g572 ( 
.A1(n_504),
.A2(n_413),
.B1(n_252),
.B2(n_311),
.Y(n_572)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_466),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_489),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_433),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_436),
.B(n_422),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_433),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_467),
.Y(n_578)
);

INVxp33_ASAP7_75t_L g579 ( 
.A(n_487),
.Y(n_579)
);

AND2x2_ASAP7_75t_SL g580 ( 
.A(n_468),
.B(n_230),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_489),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_442),
.Y(n_582)
);

AO22x2_ASAP7_75t_L g583 ( 
.A1(n_470),
.A2(n_413),
.B1(n_252),
.B2(n_311),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_493),
.Y(n_584)
);

AND2x6_ASAP7_75t_L g585 ( 
.A(n_481),
.B(n_230),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_440),
.B(n_500),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_482),
.B(n_380),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_482),
.B(n_386),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_440),
.B(n_387),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_433),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_444),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_444),
.Y(n_592)
);

INVxp33_ASAP7_75t_SL g593 ( 
.A(n_487),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_437),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_432),
.A2(n_306),
.B1(n_240),
.B2(n_330),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_470),
.B(n_396),
.Y(n_596)
);

AND2x6_ASAP7_75t_L g597 ( 
.A(n_481),
.B(n_270),
.Y(n_597)
);

INVx8_ASAP7_75t_L g598 ( 
.A(n_432),
.Y(n_598)
);

NAND3xp33_ASAP7_75t_L g599 ( 
.A(n_484),
.B(n_407),
.C(n_400),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_493),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_481),
.B(n_270),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_475),
.B(n_412),
.Y(n_602)
);

AND2x6_ASAP7_75t_L g603 ( 
.A(n_481),
.B(n_281),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_475),
.B(n_420),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_493),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_490),
.B(n_281),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_444),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_494),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_432),
.A2(n_307),
.B1(n_234),
.B2(n_242),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_500),
.B(n_416),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_440),
.B(n_365),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_460),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_468),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_433),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_460),
.Y(n_615)
);

AO22x2_ASAP7_75t_L g616 ( 
.A1(n_492),
.A2(n_306),
.B1(n_284),
.B2(n_242),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_440),
.B(n_363),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_492),
.B(n_255),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_432),
.A2(n_326),
.B1(n_289),
.B2(n_307),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_440),
.B(n_365),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_437),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_440),
.B(n_401),
.Y(n_622)
);

NAND3xp33_ASAP7_75t_L g623 ( 
.A(n_468),
.B(n_203),
.C(n_187),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_444),
.Y(n_624)
);

NAND3xp33_ASAP7_75t_L g625 ( 
.A(n_436),
.B(n_208),
.C(n_204),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_432),
.A2(n_490),
.B1(n_495),
.B2(n_436),
.Y(n_626)
);

AND2x6_ASAP7_75t_L g627 ( 
.A(n_490),
.B(n_286),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_460),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_440),
.B(n_426),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_446),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_463),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_440),
.B(n_427),
.Y(n_632)
);

INVxp33_ASAP7_75t_L g633 ( 
.A(n_463),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_432),
.A2(n_326),
.B1(n_288),
.B2(n_289),
.Y(n_634)
);

BUFx6f_ASAP7_75t_SL g635 ( 
.A(n_490),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_432),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_446),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_463),
.B(n_255),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_490),
.Y(n_639)
);

BUFx4f_ASAP7_75t_L g640 ( 
.A(n_500),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_494),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_440),
.B(n_179),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_490),
.B(n_397),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_494),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_496),
.Y(n_645)
);

OR2x6_ASAP7_75t_L g646 ( 
.A(n_495),
.B(n_257),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_495),
.A2(n_284),
.B1(n_288),
.B2(n_308),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_446),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_495),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_496),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_437),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_500),
.B(n_221),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_500),
.B(n_259),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_500),
.B(n_312),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_496),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_495),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_495),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_656),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_511),
.A2(n_408),
.B1(n_369),
.B2(n_391),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_570),
.B(n_499),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_513),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_542),
.B(n_297),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_573),
.B(n_499),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_536),
.B(n_499),
.Y(n_664)
);

NAND3xp33_ASAP7_75t_L g665 ( 
.A(n_558),
.B(n_218),
.C(n_215),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_633),
.B(n_359),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_656),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_639),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_525),
.B(n_366),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_553),
.A2(n_283),
.B1(n_257),
.B2(n_308),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_553),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_537),
.B(n_499),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_581),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_537),
.B(n_499),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_526),
.B(n_499),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_558),
.B(n_271),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_615),
.B(n_359),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_532),
.A2(n_392),
.B1(n_290),
.B2(n_319),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_639),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_581),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_649),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_649),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_631),
.B(n_422),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_545),
.Y(n_684)
);

BUFx6f_ASAP7_75t_SL g685 ( 
.A(n_580),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_L g686 ( 
.A(n_510),
.B(n_274),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_605),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_524),
.B(n_359),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_527),
.B(n_604),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_526),
.B(n_483),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_534),
.B(n_276),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_L g692 ( 
.A1(n_618),
.A2(n_264),
.B1(n_254),
.B2(n_314),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_512),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_526),
.B(n_483),
.Y(n_694)
);

OR2x6_ASAP7_75t_L g695 ( 
.A(n_552),
.B(n_283),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_605),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_552),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_548),
.B(n_483),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_631),
.B(n_483),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_512),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_608),
.Y(n_701)
);

NAND3xp33_ASAP7_75t_L g702 ( 
.A(n_516),
.B(n_232),
.C(n_227),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_560),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_608),
.Y(n_704)
);

BUFx8_ASAP7_75t_L g705 ( 
.A(n_612),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_641),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_547),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_509),
.B(n_514),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_641),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_644),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_509),
.B(n_514),
.Y(n_711)
);

NAND3xp33_ASAP7_75t_L g712 ( 
.A(n_561),
.B(n_241),
.C(n_237),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_509),
.B(n_483),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_514),
.B(n_483),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_575),
.B(n_445),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_579),
.B(n_520),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_547),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_644),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_575),
.B(n_445),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_612),
.Y(n_720)
);

NOR3xp33_ASAP7_75t_L g721 ( 
.A(n_623),
.B(n_249),
.C(n_248),
.Y(n_721)
);

NAND2xp33_ASAP7_75t_L g722 ( 
.A(n_510),
.B(n_557),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_562),
.B(n_250),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_568),
.B(n_256),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_534),
.B(n_512),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_576),
.B(n_646),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_513),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_645),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_507),
.A2(n_330),
.B1(n_329),
.B2(n_322),
.Y(n_729)
);

NAND3xp33_ASAP7_75t_L g730 ( 
.A(n_625),
.B(n_262),
.C(n_261),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_610),
.A2(n_293),
.B1(n_277),
.B2(n_280),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_645),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_515),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_534),
.B(n_512),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_515),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_L g736 ( 
.A(n_510),
.B(n_287),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_507),
.A2(n_329),
.B1(n_322),
.B2(n_314),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_596),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_650),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_575),
.B(n_445),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_576),
.B(n_198),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_512),
.B(n_294),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_628),
.B(n_198),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_546),
.B(n_295),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_R g745 ( 
.A(n_528),
.B(n_298),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_580),
.A2(n_519),
.B1(n_657),
.B2(n_602),
.Y(n_746)
);

OR2x6_ASAP7_75t_L g747 ( 
.A(n_638),
.B(n_618),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_577),
.B(n_447),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_638),
.B(n_423),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_546),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_577),
.B(n_590),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_517),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_577),
.B(n_447),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_646),
.B(n_423),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_590),
.B(n_447),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_590),
.B(n_485),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_614),
.B(n_485),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_518),
.A2(n_316),
.B1(n_324),
.B2(n_327),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_614),
.B(n_485),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_587),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_614),
.B(n_485),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_628),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_521),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_650),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_588),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_657),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_546),
.B(n_486),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_546),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_546),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_567),
.Y(n_770)
);

NAND2xp33_ASAP7_75t_L g771 ( 
.A(n_510),
.B(n_300),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_519),
.A2(n_309),
.B1(n_334),
.B2(n_332),
.Y(n_772)
);

NAND3xp33_ASAP7_75t_SL g773 ( 
.A(n_613),
.B(n_272),
.C(n_318),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_574),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_584),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_600),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_655),
.Y(n_777)
);

NAND2x1_ASAP7_75t_L g778 ( 
.A(n_506),
.B(n_453),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_518),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_540),
.A2(n_316),
.B1(n_324),
.B2(n_327),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_519),
.B(n_198),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_540),
.A2(n_286),
.B1(n_503),
.B2(n_497),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_550),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_508),
.B(n_263),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_550),
.B(n_486),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_626),
.B(n_302),
.Y(n_786)
);

OR2x6_ASAP7_75t_L g787 ( 
.A(n_638),
.B(n_424),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_551),
.B(n_486),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_551),
.B(n_486),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_599),
.B(n_549),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_556),
.B(n_488),
.Y(n_791)
);

INVx8_ASAP7_75t_L g792 ( 
.A(n_510),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_556),
.Y(n_793)
);

INVx4_ASAP7_75t_L g794 ( 
.A(n_544),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_569),
.A2(n_503),
.B1(n_497),
.B2(n_505),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_569),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_519),
.B(n_643),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_578),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_578),
.B(n_488),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_601),
.B(n_488),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_601),
.B(n_488),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_601),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_646),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_638),
.B(n_198),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_652),
.B(n_505),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_616),
.A2(n_503),
.B1(n_497),
.B2(n_505),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_654),
.B(n_653),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_510),
.B(n_505),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_618),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_642),
.B(n_448),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_522),
.B(n_323),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_646),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_521),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_636),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_523),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_522),
.B(n_331),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_522),
.B(n_336),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_593),
.B(n_268),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_593),
.B(n_275),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_583),
.B(n_199),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_SL g821 ( 
.A(n_528),
.B(n_199),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_523),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_547),
.B(n_448),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_529),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_557),
.B(n_448),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_583),
.B(n_199),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_659),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_693),
.B(n_506),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_689),
.A2(n_635),
.B1(n_603),
.B2(n_564),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_689),
.B(n_629),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_673),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_703),
.B(n_632),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_746),
.B(n_640),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_814),
.Y(n_834)
);

AOI21x1_ASAP7_75t_L g835 ( 
.A1(n_691),
.A2(n_589),
.B(n_555),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_680),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_672),
.A2(n_640),
.B1(n_635),
.B2(n_636),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_769),
.B(n_557),
.Y(n_838)
);

BUFx4f_ASAP7_75t_L g839 ( 
.A(n_747),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_708),
.A2(n_640),
.B(n_711),
.Y(n_840)
);

NAND2x1p5_ASAP7_75t_L g841 ( 
.A(n_814),
.B(n_506),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_751),
.A2(n_598),
.B(n_544),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_662),
.A2(n_676),
.B(n_786),
.C(n_674),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_696),
.Y(n_844)
);

AO21x2_ASAP7_75t_L g845 ( 
.A1(n_742),
.A2(n_622),
.B(n_617),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_794),
.A2(n_598),
.B(n_544),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_794),
.A2(n_598),
.B(n_544),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_807),
.B(n_671),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_767),
.A2(n_598),
.B(n_522),
.Y(n_849)
);

O2A1O1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_662),
.A2(n_618),
.B(n_535),
.C(n_647),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_671),
.B(n_557),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_696),
.Y(n_852)
);

O2A1O1Ixp5_ASAP7_75t_L g853 ( 
.A1(n_742),
.A2(n_611),
.B(n_620),
.C(n_586),
.Y(n_853)
);

AO21x1_ASAP7_75t_L g854 ( 
.A1(n_744),
.A2(n_691),
.B(n_674),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_782),
.B(n_557),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_684),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_693),
.A2(n_522),
.B(n_559),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_693),
.A2(n_559),
.B(n_535),
.Y(n_858)
);

BUFx12f_ASAP7_75t_L g859 ( 
.A(n_705),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_693),
.B(n_559),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_790),
.A2(n_539),
.B(n_533),
.C(n_609),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_814),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_684),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_782),
.B(n_557),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_683),
.B(n_564),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_683),
.B(n_564),
.Y(n_866)
);

NOR3xp33_ASAP7_75t_L g867 ( 
.A(n_773),
.B(n_797),
.C(n_818),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_758),
.A2(n_635),
.B1(n_619),
.B2(n_634),
.Y(n_868)
);

BUFx8_ASAP7_75t_SL g869 ( 
.A(n_669),
.Y(n_869)
);

OAI21xp33_ASAP7_75t_L g870 ( 
.A1(n_818),
.A2(n_572),
.B(n_583),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_813),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_758),
.A2(n_595),
.B1(n_616),
.B2(n_541),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_700),
.B(n_594),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_676),
.A2(n_491),
.B(n_648),
.C(n_637),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_779),
.B(n_564),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_720),
.B(n_278),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_779),
.B(n_564),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_700),
.B(n_594),
.Y(n_878)
);

OAI321xp33_ASAP7_75t_L g879 ( 
.A1(n_692),
.A2(n_425),
.A3(n_428),
.B1(n_616),
.B2(n_572),
.C(n_583),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_700),
.A2(n_651),
.B(n_621),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_750),
.A2(n_651),
.B(n_621),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_796),
.B(n_564),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_750),
.B(n_594),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_750),
.A2(n_594),
.B(n_637),
.Y(n_884)
);

O2A1O1Ixp5_ASAP7_75t_L g885 ( 
.A1(n_744),
.A2(n_491),
.B(n_630),
.C(n_531),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_720),
.B(n_572),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_SL g887 ( 
.A1(n_664),
.A2(n_491),
.B(n_630),
.C(n_531),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_780),
.A2(n_616),
.B1(n_572),
.B2(n_624),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_726),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_675),
.A2(n_585),
.B(n_627),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_796),
.B(n_585),
.Y(n_891)
);

AOI21xp33_ASAP7_75t_L g892 ( 
.A1(n_784),
.A2(n_296),
.B(n_279),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_716),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_813),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_690),
.A2(n_585),
.B(n_627),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_750),
.B(n_594),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_798),
.B(n_585),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_768),
.A2(n_538),
.B(n_529),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_809),
.B(n_282),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_741),
.B(n_425),
.Y(n_900)
);

OAI21xp33_ASAP7_75t_L g901 ( 
.A1(n_819),
.A2(n_292),
.B(n_285),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_768),
.A2(n_648),
.B(n_563),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_790),
.A2(n_554),
.B(n_624),
.C(n_607),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_768),
.A2(n_543),
.B(n_607),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_768),
.A2(n_563),
.B(n_554),
.Y(n_905)
);

OAI321xp33_ASAP7_75t_L g906 ( 
.A1(n_692),
.A2(n_476),
.A3(n_459),
.B1(n_451),
.B2(n_452),
.C(n_480),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_786),
.A2(n_543),
.B(n_530),
.C(n_538),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_687),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_660),
.A2(n_530),
.B(n_571),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_822),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_663),
.A2(n_565),
.B(n_582),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_694),
.A2(n_627),
.B(n_606),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_762),
.B(n_459),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_785),
.A2(n_627),
.B(n_606),
.Y(n_914)
);

OAI321xp33_ASAP7_75t_L g915 ( 
.A1(n_784),
.A2(n_723),
.A3(n_724),
.B1(n_819),
.B2(n_826),
.C(n_820),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_798),
.B(n_585),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_814),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_726),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_738),
.B(n_291),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_701),
.B(n_585),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_780),
.A2(n_566),
.B1(n_571),
.B2(n_591),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_698),
.B(n_566),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_725),
.A2(n_592),
.B(n_591),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_704),
.B(n_706),
.Y(n_924)
);

OAI22xp33_ASAP7_75t_L g925 ( 
.A1(n_747),
.A2(n_317),
.B1(n_310),
.B2(n_305),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_734),
.A2(n_592),
.B(n_446),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_734),
.A2(n_430),
.B(n_450),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_709),
.B(n_597),
.Y(n_928)
);

OAI321xp33_ASAP7_75t_L g929 ( 
.A1(n_723),
.A2(n_476),
.A3(n_459),
.B1(n_451),
.B2(n_452),
.C(n_462),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_760),
.B(n_320),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_756),
.A2(n_430),
.B(n_450),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_765),
.B(n_321),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_757),
.A2(n_430),
.B(n_450),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_792),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_766),
.B(n_472),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_658),
.B(n_335),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_788),
.A2(n_791),
.B(n_789),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_724),
.A2(n_476),
.B(n_451),
.C(n_452),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_759),
.A2(n_430),
.B(n_450),
.Y(n_939)
);

OAI21xp33_ASAP7_75t_L g940 ( 
.A1(n_821),
.A2(n_338),
.B(n_462),
.Y(n_940)
);

OAI22x1_ASAP7_75t_L g941 ( 
.A1(n_697),
.A2(n_743),
.B1(n_781),
.B2(n_678),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_710),
.B(n_597),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_667),
.B(n_14),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_718),
.B(n_597),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_783),
.B(n_472),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_688),
.A2(n_469),
.B(n_462),
.C(n_473),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_728),
.B(n_597),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_732),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_793),
.A2(n_453),
.B(n_434),
.C(n_458),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_677),
.B(n_462),
.Y(n_950)
);

AOI21x1_ASAP7_75t_L g951 ( 
.A1(n_799),
.A2(n_458),
.B(n_473),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_761),
.A2(n_458),
.B(n_434),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_805),
.A2(n_458),
.B(n_434),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_739),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_764),
.B(n_597),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_713),
.A2(n_627),
.B(n_606),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_770),
.Y(n_957)
);

OR2x6_ASAP7_75t_L g958 ( 
.A(n_747),
.B(n_469),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_774),
.B(n_597),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_714),
.A2(n_434),
.B(n_453),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_775),
.B(n_603),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_776),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_777),
.B(n_603),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_715),
.A2(n_434),
.B(n_453),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_688),
.B(n_603),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_802),
.A2(n_469),
.B(n_473),
.C(n_480),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_754),
.B(n_603),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_665),
.A2(n_469),
.B(n_473),
.C(n_480),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_749),
.B(n_14),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_670),
.B(n_603),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_668),
.B(n_15),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_804),
.B(n_480),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_707),
.B(n_478),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_719),
.A2(n_434),
.B(n_453),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_740),
.A2(n_453),
.B(n_438),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_679),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_800),
.A2(n_627),
.B(n_606),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_745),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_707),
.B(n_478),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_717),
.B(n_478),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_822),
.Y(n_981)
);

OR2x6_ASAP7_75t_L g982 ( 
.A(n_787),
.B(n_478),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_681),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_801),
.A2(n_606),
.B(n_501),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_699),
.A2(n_606),
.B(n_22),
.C(n_24),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_682),
.A2(n_803),
.B1(n_812),
.B2(n_754),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_670),
.A2(n_478),
.B1(n_474),
.B2(n_472),
.Y(n_987)
);

NOR2x1p5_ASAP7_75t_SL g988 ( 
.A(n_661),
.B(n_501),
.Y(n_988)
);

AND2x6_ASAP7_75t_SL g989 ( 
.A(n_695),
.B(n_787),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_787),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_727),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_695),
.B(n_17),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_729),
.A2(n_478),
.B1(n_474),
.B2(n_472),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_824),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_729),
.B(n_478),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_666),
.A2(n_478),
.B(n_474),
.C(n_472),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_685),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_748),
.A2(n_437),
.B(n_438),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_733),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_792),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_730),
.Y(n_1001)
);

AO21x2_ASAP7_75t_L g1002 ( 
.A1(n_811),
.A2(n_501),
.B(n_107),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_737),
.B(n_478),
.Y(n_1003)
);

NOR2xp67_ASAP7_75t_L g1004 ( 
.A(n_712),
.B(n_103),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_666),
.A2(n_472),
.B(n_474),
.C(n_443),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_737),
.B(n_717),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_795),
.B(n_474),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_753),
.A2(n_437),
.B(n_438),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_755),
.A2(n_437),
.B(n_438),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_722),
.A2(n_437),
.B(n_438),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_R g1011 ( 
.A(n_792),
.B(n_97),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_848),
.B(n_795),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_893),
.B(n_685),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_915),
.A2(n_721),
.B(n_702),
.C(n_823),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_863),
.B(n_772),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_844),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_832),
.B(n_731),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_867),
.B(n_808),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_867),
.A2(n_771),
.B1(n_736),
.B2(n_686),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_SL g1020 ( 
.A1(n_971),
.A2(n_806),
.B(n_810),
.C(n_825),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_917),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_830),
.B(n_806),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_918),
.B(n_735),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_892),
.A2(n_817),
.B(n_816),
.C(n_811),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_SL g1025 ( 
.A1(n_971),
.A2(n_763),
.B(n_752),
.C(n_815),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_900),
.B(n_924),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_852),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_872),
.A2(n_817),
.B1(n_816),
.B2(n_778),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_917),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_841),
.A2(n_437),
.B(n_443),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_908),
.B(n_472),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_SL g1032 ( 
.A1(n_965),
.A2(n_501),
.B(n_110),
.C(n_111),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_948),
.B(n_472),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_843),
.A2(n_472),
.B(n_474),
.C(n_443),
.Y(n_1034)
);

NAND2x1p5_ASAP7_75t_L g1035 ( 
.A(n_934),
.B(n_474),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_934),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_954),
.B(n_474),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_901),
.A2(n_17),
.B(n_30),
.C(n_32),
.Y(n_1038)
);

OAI22x1_ASAP7_75t_L g1039 ( 
.A1(n_886),
.A2(n_33),
.B1(n_36),
.B2(n_40),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_841),
.A2(n_437),
.B(n_443),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_913),
.B(n_474),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_871),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_SL g1043 ( 
.A(n_868),
.B(n_501),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_972),
.B(n_438),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_838),
.A2(n_438),
.B(n_443),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_831),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_R g1047 ( 
.A(n_978),
.B(n_112),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_SL g1048 ( 
.A(n_839),
.B(n_501),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_957),
.B(n_438),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_967),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_833),
.A2(n_438),
.B(n_443),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_934),
.Y(n_1052)
);

INVxp67_ASAP7_75t_L g1053 ( 
.A(n_876),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_834),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_967),
.B(n_443),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_R g1056 ( 
.A(n_827),
.B(n_92),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_836),
.B(n_443),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_850),
.A2(n_443),
.B(n_455),
.C(n_457),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_958),
.Y(n_1059)
);

INVx4_ASAP7_75t_L g1060 ( 
.A(n_934),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_857),
.A2(n_455),
.B(n_457),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_889),
.B(n_455),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_969),
.A2(n_919),
.B(n_925),
.C(n_899),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_856),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_894),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_858),
.A2(n_455),
.B(n_457),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_930),
.B(n_40),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_840),
.A2(n_828),
.B(n_860),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_828),
.A2(n_455),
.B(n_457),
.Y(n_1069)
);

O2A1O1Ixp5_ASAP7_75t_L g1070 ( 
.A1(n_854),
.A2(n_90),
.B(n_173),
.C(n_168),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_937),
.B(n_457),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_950),
.B(n_457),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_888),
.B(n_457),
.Y(n_1073)
);

AO32x2_ASAP7_75t_L g1074 ( 
.A1(n_921),
.A2(n_42),
.A3(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_969),
.A2(n_455),
.B(n_457),
.C(n_54),
.Y(n_1075)
);

AO21x1_ASAP7_75t_L g1076 ( 
.A1(n_1006),
.A2(n_42),
.B(n_50),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_1001),
.B(n_455),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_932),
.B(n_54),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_962),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_834),
.B(n_455),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_919),
.B(n_57),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_910),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_870),
.B(n_57),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_925),
.A2(n_58),
.B(n_61),
.C(n_62),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_932),
.B(n_61),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_876),
.B(n_65),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_981),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_879),
.B(n_119),
.Y(n_1088)
);

INVx1_ASAP7_75t_SL g1089 ( 
.A(n_992),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_899),
.A2(n_65),
.B(n_66),
.C(n_501),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_936),
.B(n_66),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_990),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_861),
.A2(n_68),
.B(n_71),
.C(n_77),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_994),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_976),
.B(n_501),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_859),
.Y(n_1096)
);

OAI22x1_ASAP7_75t_L g1097 ( 
.A1(n_986),
.A2(n_78),
.B1(n_79),
.B2(n_89),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_990),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_842),
.A2(n_847),
.B(n_846),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_983),
.A2(n_501),
.B1(n_116),
.B2(n_120),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_849),
.A2(n_113),
.B(n_125),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_R g1102 ( 
.A(n_997),
.B(n_862),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_941),
.B(n_839),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_991),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_999),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_936),
.B(n_126),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_970),
.A2(n_501),
.B1(n_144),
.B2(n_146),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_890),
.A2(n_141),
.B(n_157),
.Y(n_1108)
);

HB1xp67_ASAP7_75t_L g1109 ( 
.A(n_958),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_855),
.A2(n_159),
.B(n_164),
.C(n_501),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_966),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_865),
.B(n_501),
.Y(n_1112)
);

INVx4_ASAP7_75t_L g1113 ( 
.A(n_1000),
.Y(n_1113)
);

INVx3_ASAP7_75t_SL g1114 ( 
.A(n_958),
.Y(n_1114)
);

BUFx12f_ASAP7_75t_L g1115 ( 
.A(n_989),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_895),
.A2(n_912),
.B(n_977),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_943),
.A2(n_985),
.B(n_940),
.C(n_938),
.Y(n_1117)
);

OAI21xp33_ASAP7_75t_L g1118 ( 
.A1(n_866),
.A2(n_864),
.B(n_961),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_829),
.A2(n_914),
.B(n_963),
.C(n_959),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_982),
.A2(n_1007),
.B1(n_1003),
.B2(n_995),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_851),
.A2(n_956),
.B(n_896),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_920),
.A2(n_928),
.B(n_955),
.C(n_942),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_982),
.A2(n_862),
.B1(n_875),
.B2(n_882),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_1000),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1000),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_869),
.B(n_906),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_922),
.B(n_845),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1011),
.B(n_944),
.Y(n_1128)
);

CKINVDCx6p67_ASAP7_75t_R g1129 ( 
.A(n_982),
.Y(n_1129)
);

BUFx4f_ASAP7_75t_L g1130 ( 
.A(n_1000),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_946),
.A2(n_1005),
.B(n_996),
.C(n_903),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_947),
.A2(n_874),
.B(n_885),
.C(n_929),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_951),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_877),
.B(n_916),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_845),
.A2(n_1004),
.B1(n_891),
.B2(n_897),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_945),
.Y(n_1136)
);

INVxp67_ASAP7_75t_SL g1137 ( 
.A(n_873),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1011),
.Y(n_1138)
);

INVx4_ASAP7_75t_L g1139 ( 
.A(n_1002),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_873),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_907),
.A2(n_984),
.B(n_949),
.C(n_923),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_837),
.B(n_973),
.Y(n_1142)
);

BUFx12f_ASAP7_75t_L g1143 ( 
.A(n_988),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_973),
.B(n_980),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_878),
.A2(n_883),
.B(n_896),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_968),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_926),
.A2(n_960),
.B(n_853),
.C(n_974),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_945),
.B(n_935),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_935),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_922),
.B(n_883),
.Y(n_1150)
);

AOI22x1_ASAP7_75t_L g1151 ( 
.A1(n_909),
.A2(n_911),
.B1(n_953),
.B2(n_964),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_878),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_SL g1153 ( 
.A1(n_1010),
.A2(n_884),
.B(n_905),
.C(n_904),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_927),
.A2(n_952),
.B(n_975),
.C(n_902),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_979),
.B(n_980),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_987),
.A2(n_993),
.B1(n_880),
.B2(n_881),
.Y(n_1156)
);

CKINVDCx8_ASAP7_75t_R g1157 ( 
.A(n_1002),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_887),
.A2(n_898),
.B(n_1009),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_931),
.A2(n_933),
.B1(n_939),
.B2(n_998),
.Y(n_1159)
);

INVxp67_ASAP7_75t_L g1160 ( 
.A(n_1008),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_835),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_841),
.A2(n_640),
.B(n_794),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_841),
.A2(n_640),
.B(n_794),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_918),
.B(n_889),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_967),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1116),
.A2(n_1058),
.B(n_1119),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1162),
.A2(n_1163),
.B(n_1132),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1063),
.A2(n_1106),
.B(n_1078),
.C(n_1085),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1068),
.A2(n_1099),
.B(n_1158),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_SL g1170 ( 
.A1(n_1076),
.A2(n_1108),
.B(n_1038),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1034),
.A2(n_1120),
.B(n_1160),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_SL g1172 ( 
.A1(n_1093),
.A2(n_1020),
.B(n_1088),
.C(n_1081),
.Y(n_1172)
);

AOI221x1_ASAP7_75t_L g1173 ( 
.A1(n_1091),
.A2(n_1086),
.B1(n_1075),
.B2(n_1028),
.C(n_1147),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1151),
.A2(n_1051),
.B(n_1121),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1161),
.A2(n_1139),
.A3(n_1141),
.B(n_1123),
.Y(n_1175)
);

OR2x6_ASAP7_75t_L g1176 ( 
.A(n_1138),
.B(n_1059),
.Y(n_1176)
);

OA21x2_ASAP7_75t_L g1177 ( 
.A1(n_1127),
.A2(n_1142),
.B(n_1071),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1022),
.B(n_1026),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_1139),
.A2(n_1123),
.A3(n_1156),
.B(n_1127),
.Y(n_1179)
);

NAND2xp33_ASAP7_75t_R g1180 ( 
.A(n_1102),
.B(n_1047),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1094),
.Y(n_1181)
);

NAND2xp33_ASAP7_75t_L g1182 ( 
.A(n_1026),
.B(n_1050),
.Y(n_1182)
);

AO31x2_ASAP7_75t_L g1183 ( 
.A1(n_1156),
.A2(n_1120),
.A3(n_1028),
.B(n_1154),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_1064),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1145),
.A2(n_1045),
.B(n_1066),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1019),
.A2(n_1024),
.B(n_1128),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1072),
.A2(n_1017),
.B(n_1012),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1072),
.A2(n_1012),
.B(n_1153),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1042),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1053),
.A2(n_1084),
.B(n_1067),
.C(n_1103),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1015),
.B(n_1164),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1131),
.A2(n_1018),
.B(n_1122),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1089),
.B(n_1126),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1134),
.A2(n_1071),
.B(n_1044),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_SL g1195 ( 
.A(n_1130),
.B(n_1021),
.Y(n_1195)
);

NAND2xp33_ASAP7_75t_L g1196 ( 
.A(n_1050),
.B(n_1165),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1056),
.B(n_1164),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1118),
.A2(n_1117),
.B(n_1144),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1014),
.A2(n_1146),
.B(n_1135),
.Y(n_1199)
);

AOI221xp5_ASAP7_75t_SL g1200 ( 
.A1(n_1039),
.A2(n_1090),
.B1(n_1022),
.B2(n_1083),
.C(n_1073),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1150),
.A2(n_1155),
.B(n_1073),
.Y(n_1201)
);

NOR2x1_ASAP7_75t_R g1202 ( 
.A(n_1096),
.B(n_1115),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_SL g1203 ( 
.A1(n_1097),
.A2(n_1052),
.B(n_1113),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1098),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1105),
.B(n_1046),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1065),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1104),
.B(n_1016),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1027),
.B(n_1082),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1070),
.A2(n_1111),
.B(n_1150),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1092),
.B(n_1109),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1159),
.A2(n_1025),
.B(n_1101),
.Y(n_1211)
);

AO21x2_ASAP7_75t_L g1212 ( 
.A1(n_1133),
.A2(n_1032),
.B(n_1061),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1165),
.B(n_1023),
.Y(n_1213)
);

OR2x2_ASAP7_75t_L g1214 ( 
.A(n_1114),
.B(n_1087),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_1130),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1137),
.A2(n_1043),
.B(n_1080),
.Y(n_1216)
);

BUFx4f_ASAP7_75t_L g1217 ( 
.A(n_1125),
.Y(n_1217)
);

AO32x2_ASAP7_75t_L g1218 ( 
.A1(n_1074),
.A2(n_1157),
.A3(n_1021),
.B1(n_1036),
.B2(n_1113),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1043),
.A2(n_1110),
.B(n_1149),
.C(n_1107),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1049),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1023),
.B(n_1041),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1069),
.A2(n_1057),
.B(n_1030),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1148),
.A2(n_1057),
.B(n_1112),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1059),
.B(n_1129),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1140),
.B(n_1152),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1040),
.A2(n_1080),
.B(n_1031),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1140),
.B(n_1152),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1055),
.A2(n_1077),
.B(n_1033),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1037),
.A2(n_1062),
.B(n_1029),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1136),
.A2(n_1095),
.B(n_1100),
.C(n_1054),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1048),
.A2(n_1035),
.B(n_1054),
.Y(n_1231)
);

OAI22x1_ASAP7_75t_L g1232 ( 
.A1(n_1074),
.A2(n_1060),
.B1(n_1036),
.B2(n_1124),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1035),
.A2(n_1143),
.B(n_1052),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1048),
.A2(n_1060),
.B(n_1124),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1059),
.Y(n_1235)
);

BUFx8_ASAP7_75t_L g1236 ( 
.A(n_1125),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1074),
.Y(n_1237)
);

NOR2xp67_ASAP7_75t_L g1238 ( 
.A(n_1053),
.B(n_684),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1099),
.A2(n_1158),
.B(n_1068),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1026),
.B(n_689),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1022),
.B(n_689),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_SL g1242 ( 
.A1(n_1093),
.A2(n_1106),
.B(n_1063),
.C(n_1020),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1125),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1053),
.B(n_703),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1102),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1099),
.A2(n_1158),
.B(n_1068),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1034),
.A2(n_1058),
.A3(n_854),
.B(n_1161),
.Y(n_1247)
);

AOI221xp5_ASAP7_75t_L g1248 ( 
.A1(n_1091),
.A2(n_692),
.B1(n_1063),
.B2(n_1086),
.C(n_1085),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1106),
.A2(n_689),
.B1(n_669),
.B2(n_827),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1091),
.A2(n_1086),
.B1(n_511),
.B2(n_1085),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1162),
.A2(n_640),
.B(n_693),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1099),
.A2(n_1158),
.B(n_1068),
.Y(n_1252)
);

BUFx12f_ASAP7_75t_L g1253 ( 
.A(n_1096),
.Y(n_1253)
);

CKINVDCx6p67_ASAP7_75t_R g1254 ( 
.A(n_1096),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1036),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1079),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1162),
.A2(n_640),
.B(n_693),
.Y(n_1257)
);

CKINVDCx6p67_ASAP7_75t_R g1258 ( 
.A(n_1096),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1064),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1026),
.A2(n_780),
.B1(n_758),
.B2(n_511),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1099),
.A2(n_1158),
.B(n_1068),
.Y(n_1261)
);

AO21x1_ASAP7_75t_L g1262 ( 
.A1(n_1063),
.A2(n_1106),
.B(n_830),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1116),
.A2(n_1058),
.B(n_1119),
.Y(n_1263)
);

NAND2xp33_ASAP7_75t_L g1264 ( 
.A(n_1081),
.B(n_1011),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1022),
.B(n_689),
.Y(n_1265)
);

AOI221xp5_ASAP7_75t_SL g1266 ( 
.A1(n_1063),
.A2(n_1091),
.B1(n_1078),
.B2(n_1085),
.C(n_1084),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1162),
.A2(n_640),
.B(n_693),
.Y(n_1267)
);

INVxp67_ASAP7_75t_SL g1268 ( 
.A(n_1026),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1053),
.B(n_525),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_SL g1270 ( 
.A1(n_1093),
.A2(n_1106),
.B(n_1063),
.C(n_1020),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1079),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1089),
.B(n_525),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1064),
.Y(n_1273)
);

AOI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1142),
.A2(n_835),
.B(n_1018),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1026),
.B(n_689),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1053),
.B(n_525),
.Y(n_1276)
);

AOI31xp67_ASAP7_75t_L g1277 ( 
.A1(n_1133),
.A2(n_1142),
.A3(n_1019),
.B(n_1135),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1099),
.A2(n_1158),
.B(n_1068),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1026),
.B(n_689),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1162),
.A2(n_640),
.B(n_693),
.Y(n_1280)
);

O2A1O1Ixp33_ASAP7_75t_SL g1281 ( 
.A1(n_1093),
.A2(n_1106),
.B(n_1063),
.C(n_1020),
.Y(n_1281)
);

AO21x2_ASAP7_75t_L g1282 ( 
.A1(n_1034),
.A2(n_1058),
.B(n_1116),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1026),
.A2(n_780),
.B1(n_758),
.B2(n_511),
.Y(n_1283)
);

BUFx10_ASAP7_75t_L g1284 ( 
.A(n_1013),
.Y(n_1284)
);

BUFx2_ASAP7_75t_R g1285 ( 
.A(n_1096),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1099),
.A2(n_1158),
.B(n_1068),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1162),
.A2(n_640),
.B(n_693),
.Y(n_1287)
);

AO21x2_ASAP7_75t_L g1288 ( 
.A1(n_1034),
.A2(n_1058),
.B(n_1116),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1034),
.A2(n_1058),
.A3(n_854),
.B(n_1161),
.Y(n_1289)
);

AOI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1142),
.A2(n_835),
.B(n_1018),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1026),
.B(n_689),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1162),
.A2(n_640),
.B(n_693),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1162),
.A2(n_640),
.B(n_693),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1089),
.B(n_545),
.Y(n_1294)
);

A2O1A1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1063),
.A2(n_511),
.B(n_689),
.C(n_1106),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1099),
.A2(n_1158),
.B(n_1068),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1099),
.A2(n_1158),
.B(n_1068),
.Y(n_1297)
);

O2A1O1Ixp5_ASAP7_75t_L g1298 ( 
.A1(n_1078),
.A2(n_689),
.B(n_1085),
.C(n_1091),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1053),
.B(n_703),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_SL g1300 ( 
.A1(n_1076),
.A2(n_843),
.B(n_1108),
.Y(n_1300)
);

BUFx12f_ASAP7_75t_L g1301 ( 
.A(n_1096),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1079),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1125),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1053),
.B(n_703),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1022),
.B(n_689),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1102),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1162),
.A2(n_640),
.B(n_693),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1022),
.B(n_689),
.Y(n_1308)
);

BUFx4f_ASAP7_75t_SL g1309 ( 
.A(n_1096),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1034),
.A2(n_1058),
.A3(n_854),
.B(n_1161),
.Y(n_1310)
);

NAND2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1130),
.B(n_917),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1236),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1248),
.A2(n_1250),
.B1(n_1262),
.B2(n_1249),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1240),
.A2(n_1275),
.B1(n_1291),
.B2(n_1279),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1217),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1168),
.B(n_1295),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1260),
.A2(n_1283),
.B1(n_1305),
.B2(n_1241),
.Y(n_1317)
);

BUFx12f_ASAP7_75t_L g1318 ( 
.A(n_1253),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1260),
.A2(n_1283),
.B1(n_1308),
.B2(n_1241),
.Y(n_1319)
);

CKINVDCx11_ASAP7_75t_R g1320 ( 
.A(n_1301),
.Y(n_1320)
);

INVx4_ASAP7_75t_L g1321 ( 
.A(n_1217),
.Y(n_1321)
);

INVx6_ASAP7_75t_L g1322 ( 
.A(n_1236),
.Y(n_1322)
);

BUFx4f_ASAP7_75t_L g1323 ( 
.A(n_1254),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1256),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1265),
.A2(n_1305),
.B1(n_1308),
.B2(n_1199),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1193),
.A2(n_1268),
.B1(n_1170),
.B2(n_1264),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1265),
.A2(n_1199),
.B1(n_1192),
.B2(n_1178),
.Y(n_1327)
);

BUFx8_ASAP7_75t_L g1328 ( 
.A(n_1259),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1215),
.B(n_1224),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1272),
.Y(n_1330)
);

INVx6_ASAP7_75t_L g1331 ( 
.A(n_1215),
.Y(n_1331)
);

BUFx10_ASAP7_75t_L g1332 ( 
.A(n_1245),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1192),
.A2(n_1178),
.B1(n_1198),
.B2(n_1191),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1197),
.A2(n_1182),
.B1(n_1284),
.B2(n_1300),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1271),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1184),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1273),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1166),
.A2(n_1263),
.B1(n_1186),
.B2(n_1171),
.Y(n_1338)
);

BUFx2_ASAP7_75t_SL g1339 ( 
.A(n_1306),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1189),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1302),
.Y(n_1341)
);

AOI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1266),
.A2(n_1244),
.B1(n_1304),
.B2(n_1299),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1205),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1166),
.A2(n_1263),
.B1(n_1171),
.B2(n_1201),
.Y(n_1344)
);

INVx6_ASAP7_75t_L g1345 ( 
.A(n_1243),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1180),
.Y(n_1346)
);

INVx4_ASAP7_75t_SL g1347 ( 
.A(n_1243),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1298),
.A2(n_1187),
.B1(n_1266),
.B2(n_1294),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1206),
.A2(n_1209),
.B1(n_1282),
.B2(n_1288),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1303),
.Y(n_1350)
);

BUFx10_ASAP7_75t_L g1351 ( 
.A(n_1210),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1176),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1285),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1177),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1269),
.B(n_1276),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1177),
.Y(n_1356)
);

OAI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1173),
.A2(n_1238),
.B1(n_1195),
.B2(n_1176),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1209),
.A2(n_1288),
.B1(n_1282),
.B2(n_1204),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1169),
.A2(n_1280),
.B(n_1251),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_SL g1360 ( 
.A1(n_1284),
.A2(n_1195),
.B1(n_1237),
.B2(n_1309),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1190),
.A2(n_1214),
.B1(n_1219),
.B2(n_1213),
.Y(n_1361)
);

OAI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1221),
.A2(n_1232),
.B1(n_1220),
.B2(n_1227),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1208),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1223),
.A2(n_1188),
.B1(n_1194),
.B2(n_1207),
.Y(n_1364)
);

BUFx2_ASAP7_75t_SL g1365 ( 
.A(n_1303),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1311),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1200),
.A2(n_1242),
.B1(n_1281),
.B2(n_1270),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1235),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1223),
.A2(n_1216),
.B1(n_1167),
.B2(n_1225),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1225),
.B(n_1227),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1211),
.A2(n_1228),
.B1(n_1196),
.B2(n_1229),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1212),
.A2(n_1234),
.B1(n_1255),
.B2(n_1258),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1218),
.Y(n_1373)
);

BUFx8_ASAP7_75t_L g1374 ( 
.A(n_1303),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1212),
.A2(n_1255),
.B1(n_1231),
.B2(n_1174),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1233),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1230),
.A2(n_1203),
.B1(n_1307),
.B2(n_1293),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1218),
.B(n_1183),
.Y(n_1378)
);

CKINVDCx11_ASAP7_75t_R g1379 ( 
.A(n_1202),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1175),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_SL g1381 ( 
.A1(n_1172),
.A2(n_1252),
.B1(n_1286),
.B2(n_1246),
.Y(n_1381)
);

CKINVDCx10_ASAP7_75t_R g1382 ( 
.A(n_1277),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1257),
.Y(n_1383)
);

OAI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1274),
.A2(n_1290),
.B1(n_1292),
.B2(n_1267),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1287),
.A2(n_1183),
.B1(n_1179),
.B2(n_1247),
.Y(n_1385)
);

NAND2x1p5_ASAP7_75t_L g1386 ( 
.A(n_1226),
.B(n_1222),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_SL g1387 ( 
.A1(n_1239),
.A2(n_1278),
.B1(n_1297),
.B2(n_1261),
.Y(n_1387)
);

BUFx8_ASAP7_75t_L g1388 ( 
.A(n_1289),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1289),
.B(n_1310),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1185),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1296),
.A2(n_1248),
.B1(n_1250),
.B2(n_1091),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1193),
.A2(n_1086),
.B1(n_1091),
.B2(n_821),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1193),
.A2(n_1086),
.B1(n_1091),
.B2(n_821),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1184),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1193),
.A2(n_1086),
.B1(n_1091),
.B2(n_821),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1240),
.B(n_1275),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1217),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1181),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1181),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1181),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_SL g1401 ( 
.A(n_1236),
.Y(n_1401)
);

CKINVDCx11_ASAP7_75t_R g1402 ( 
.A(n_1253),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1245),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1240),
.B(n_1275),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1240),
.B(n_1275),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1248),
.A2(n_1250),
.B1(n_1091),
.B2(n_1078),
.Y(n_1406)
);

BUFx8_ASAP7_75t_L g1407 ( 
.A(n_1253),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1181),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1240),
.B(n_1275),
.Y(n_1409)
);

CKINVDCx11_ASAP7_75t_R g1410 ( 
.A(n_1253),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1309),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1181),
.Y(n_1412)
);

BUFx4f_ASAP7_75t_SL g1413 ( 
.A(n_1253),
.Y(n_1413)
);

INVx6_ASAP7_75t_L g1414 ( 
.A(n_1236),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1193),
.A2(n_1086),
.B1(n_1091),
.B2(n_821),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1236),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1248),
.A2(n_1250),
.B1(n_1091),
.B2(n_1078),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_SL g1418 ( 
.A1(n_1249),
.A2(n_1250),
.B(n_1248),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1248),
.A2(n_1250),
.B1(n_1091),
.B2(n_1078),
.Y(n_1419)
);

BUFx10_ASAP7_75t_L g1420 ( 
.A(n_1245),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1184),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1248),
.A2(n_1250),
.B1(n_1091),
.B2(n_1078),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_SL g1423 ( 
.A(n_1250),
.B(n_1248),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1181),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1236),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1184),
.Y(n_1426)
);

AO21x2_ASAP7_75t_L g1427 ( 
.A1(n_1359),
.A2(n_1384),
.B(n_1390),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_1330),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1378),
.B(n_1316),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1354),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1386),
.A2(n_1377),
.B(n_1385),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1325),
.B(n_1314),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1388),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1388),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1325),
.B(n_1314),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1356),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1376),
.B(n_1380),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1316),
.B(n_1373),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1389),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1375),
.A2(n_1371),
.B(n_1376),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1380),
.Y(n_1441)
);

AOI211x1_ASAP7_75t_L g1442 ( 
.A1(n_1423),
.A2(n_1361),
.B(n_1409),
.C(n_1405),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1375),
.A2(n_1371),
.B(n_1349),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1324),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1344),
.A2(n_1349),
.B(n_1338),
.Y(n_1445)
);

INVx4_ASAP7_75t_L g1446 ( 
.A(n_1383),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1346),
.B(n_1342),
.Y(n_1447)
);

INVx4_ASAP7_75t_L g1448 ( 
.A(n_1366),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1317),
.B(n_1319),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1370),
.Y(n_1450)
);

INVxp33_ASAP7_75t_L g1451 ( 
.A(n_1337),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1352),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1327),
.B(n_1317),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1319),
.B(n_1338),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1358),
.B(n_1327),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1335),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1341),
.Y(n_1457)
);

CKINVDCx11_ASAP7_75t_R g1458 ( 
.A(n_1411),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1406),
.A2(n_1422),
.B1(n_1419),
.B2(n_1417),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1343),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1328),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1367),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1344),
.A2(n_1358),
.B(n_1364),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1363),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1331),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1333),
.B(n_1348),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1368),
.Y(n_1467)
);

AOI221xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1406),
.A2(n_1417),
.B1(n_1419),
.B2(n_1422),
.C(n_1313),
.Y(n_1468)
);

NAND3xp33_ASAP7_75t_L g1469 ( 
.A(n_1392),
.B(n_1393),
.C(n_1395),
.Y(n_1469)
);

NOR2x1_ASAP7_75t_SL g1470 ( 
.A(n_1418),
.B(n_1398),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1399),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1348),
.B(n_1333),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1400),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1369),
.B(n_1366),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1362),
.B(n_1313),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1391),
.B(n_1369),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1391),
.B(n_1412),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_SL g1478 ( 
.A(n_1401),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1362),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1424),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1364),
.A2(n_1372),
.B(n_1408),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1340),
.B(n_1396),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1384),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1382),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1404),
.B(n_1326),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1387),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1381),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1372),
.B(n_1360),
.Y(n_1488)
);

INVx2_ASAP7_75t_SL g1489 ( 
.A(n_1331),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1351),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1334),
.B(n_1355),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1357),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1357),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1415),
.B(n_1329),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1329),
.A2(n_1339),
.B1(n_1414),
.B2(n_1322),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1347),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1321),
.A2(n_1315),
.B(n_1397),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1347),
.Y(n_1498)
);

CKINVDCx11_ASAP7_75t_R g1499 ( 
.A(n_1320),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1421),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1331),
.Y(n_1501)
);

BUFx2_ASAP7_75t_SL g1502 ( 
.A(n_1351),
.Y(n_1502)
);

OAI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1321),
.A2(n_1426),
.B(n_1394),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1315),
.B(n_1397),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1328),
.A2(n_1336),
.B1(n_1414),
.B2(n_1322),
.Y(n_1505)
);

OA21x2_ASAP7_75t_L g1506 ( 
.A1(n_1443),
.A2(n_1353),
.B(n_1347),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1450),
.B(n_1350),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1429),
.B(n_1312),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1443),
.A2(n_1365),
.B(n_1403),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1460),
.Y(n_1510)
);

AOI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1432),
.A2(n_1414),
.B(n_1322),
.Y(n_1511)
);

O2A1O1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1459),
.A2(n_1312),
.B(n_1416),
.C(n_1425),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1459),
.A2(n_1425),
.B1(n_1416),
.B2(n_1323),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1468),
.A2(n_1323),
.B(n_1420),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1438),
.B(n_1374),
.Y(n_1515)
);

A2O1A1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1469),
.A2(n_1468),
.B(n_1447),
.C(n_1484),
.Y(n_1516)
);

O2A1O1Ixp33_ASAP7_75t_SL g1517 ( 
.A1(n_1484),
.A2(n_1379),
.B(n_1407),
.C(n_1413),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1452),
.B(n_1491),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1491),
.B(n_1345),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1469),
.A2(n_1475),
.B1(n_1442),
.B2(n_1453),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1446),
.B(n_1420),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1475),
.A2(n_1413),
.B(n_1332),
.C(n_1407),
.Y(n_1522)
);

A2O1A1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1479),
.A2(n_1410),
.B(n_1402),
.C(n_1318),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1482),
.B(n_1467),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1479),
.A2(n_1449),
.B(n_1485),
.C(n_1476),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_1500),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1461),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1477),
.B(n_1494),
.Y(n_1528)
);

INVx5_ASAP7_75t_L g1529 ( 
.A(n_1446),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1477),
.B(n_1494),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1442),
.A2(n_1453),
.B1(n_1492),
.B2(n_1493),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1446),
.B(n_1451),
.Y(n_1532)
);

AO21x1_ASAP7_75t_L g1533 ( 
.A1(n_1485),
.A2(n_1435),
.B(n_1432),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1503),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1492),
.A2(n_1493),
.B1(n_1435),
.B2(n_1449),
.Y(n_1535)
);

NAND4xp25_ASAP7_75t_L g1536 ( 
.A(n_1428),
.B(n_1490),
.C(n_1503),
.D(n_1462),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1428),
.B(n_1458),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1490),
.B(n_1478),
.Y(n_1538)
);

A2O1A1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1454),
.A2(n_1472),
.B(n_1466),
.C(n_1488),
.Y(n_1539)
);

OAI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1454),
.A2(n_1481),
.B(n_1455),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1462),
.A2(n_1445),
.B1(n_1488),
.B2(n_1495),
.Y(n_1541)
);

A2O1A1Ixp33_ASAP7_75t_L g1542 ( 
.A1(n_1455),
.A2(n_1431),
.B(n_1495),
.C(n_1433),
.Y(n_1542)
);

AO32x2_ASAP7_75t_L g1543 ( 
.A1(n_1448),
.A2(n_1489),
.A3(n_1465),
.B1(n_1501),
.B2(n_1439),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1437),
.B(n_1456),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1502),
.B(n_1499),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1481),
.A2(n_1463),
.B(n_1483),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1474),
.A2(n_1434),
.B1(n_1433),
.B2(n_1445),
.Y(n_1547)
);

INVxp33_ASAP7_75t_SL g1548 ( 
.A(n_1502),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1445),
.A2(n_1505),
.B1(n_1434),
.B2(n_1463),
.Y(n_1549)
);

OAI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1463),
.A2(n_1483),
.B(n_1440),
.Y(n_1550)
);

OA21x2_ASAP7_75t_L g1551 ( 
.A1(n_1440),
.A2(n_1431),
.B(n_1487),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1497),
.B(n_1465),
.Y(n_1552)
);

O2A1O1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1487),
.A2(n_1486),
.B(n_1497),
.C(n_1504),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1461),
.B(n_1489),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1444),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1445),
.A2(n_1431),
.B(n_1474),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1457),
.B(n_1464),
.Y(n_1557)
);

OAI211xp5_ASAP7_75t_L g1558 ( 
.A1(n_1486),
.A2(n_1471),
.B(n_1480),
.C(n_1473),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1556),
.B(n_1430),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1544),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1550),
.B(n_1430),
.Y(n_1561)
);

NOR2x1p5_ASAP7_75t_L g1562 ( 
.A(n_1536),
.B(n_1461),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1556),
.B(n_1436),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1534),
.B(n_1470),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1510),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1546),
.B(n_1540),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1558),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1548),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1555),
.Y(n_1569)
);

OAI222xp33_ASAP7_75t_L g1570 ( 
.A1(n_1520),
.A2(n_1513),
.B1(n_1535),
.B2(n_1541),
.C1(n_1531),
.C2(n_1512),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1507),
.Y(n_1571)
);

INVxp67_ASAP7_75t_SL g1572 ( 
.A(n_1557),
.Y(n_1572)
);

BUFx2_ASAP7_75t_L g1573 ( 
.A(n_1543),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1543),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1551),
.B(n_1436),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1543),
.Y(n_1576)
);

INVx4_ASAP7_75t_L g1577 ( 
.A(n_1529),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1533),
.B(n_1474),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1551),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1540),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1520),
.A2(n_1474),
.B1(n_1471),
.B2(n_1473),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1545),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1509),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1566),
.B(n_1506),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1560),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1566),
.B(n_1509),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1574),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1569),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1560),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1567),
.B(n_1529),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1575),
.Y(n_1591)
);

AOI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1570),
.A2(n_1516),
.B1(n_1539),
.B2(n_1525),
.C(n_1535),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1573),
.B(n_1549),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1575),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1572),
.B(n_1528),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1569),
.Y(n_1596)
);

AND2x4_ASAP7_75t_SL g1597 ( 
.A(n_1577),
.B(n_1565),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1566),
.B(n_1547),
.Y(n_1598)
);

OR2x6_ASAP7_75t_SL g1599 ( 
.A(n_1568),
.B(n_1549),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1573),
.B(n_1427),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1573),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1565),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1569),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1567),
.A2(n_1541),
.B1(n_1513),
.B2(n_1531),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1580),
.B(n_1427),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1580),
.B(n_1427),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1574),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1559),
.B(n_1542),
.Y(n_1608)
);

OAI221xp5_ASAP7_75t_L g1609 ( 
.A1(n_1581),
.A2(n_1514),
.B1(n_1523),
.B2(n_1522),
.C(n_1553),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1578),
.B(n_1532),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1578),
.B(n_1511),
.Y(n_1611)
);

AOI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1570),
.A2(n_1514),
.B1(n_1530),
.B2(n_1517),
.C(n_1526),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1559),
.B(n_1441),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1581),
.A2(n_1524),
.B1(n_1538),
.B2(n_1537),
.C(n_1480),
.Y(n_1614)
);

OAI222xp33_ASAP7_75t_L g1615 ( 
.A1(n_1568),
.A2(n_1515),
.B1(n_1508),
.B2(n_1518),
.C1(n_1552),
.C2(n_1519),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1591),
.Y(n_1616)
);

INVxp67_ASAP7_75t_SL g1617 ( 
.A(n_1587),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1601),
.B(n_1576),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1601),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1601),
.B(n_1583),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1595),
.B(n_1571),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1586),
.B(n_1584),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1586),
.B(n_1583),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1591),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1586),
.B(n_1583),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1610),
.B(n_1582),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1584),
.B(n_1583),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1593),
.B(n_1572),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1588),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1584),
.B(n_1579),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1588),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1600),
.B(n_1579),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1600),
.B(n_1579),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1589),
.B(n_1591),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1608),
.B(n_1559),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1594),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1593),
.B(n_1561),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1608),
.B(n_1563),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1608),
.B(n_1563),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1585),
.B(n_1563),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1596),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1610),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1602),
.Y(n_1643)
);

AND2x4_ASAP7_75t_SL g1644 ( 
.A(n_1604),
.B(n_1577),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1603),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1595),
.B(n_1571),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1600),
.B(n_1579),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1619),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1626),
.A2(n_1592),
.B1(n_1612),
.B2(n_1604),
.Y(n_1649)
);

A2O1A1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1626),
.A2(n_1612),
.B(n_1592),
.C(n_1642),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1642),
.B(n_1621),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1619),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1619),
.Y(n_1653)
);

OAI211xp5_ASAP7_75t_SL g1654 ( 
.A1(n_1621),
.A2(n_1614),
.B(n_1609),
.C(n_1611),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1635),
.B(n_1599),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1617),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1634),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1617),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1634),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1635),
.B(n_1638),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1646),
.B(n_1598),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1646),
.B(n_1598),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1643),
.Y(n_1663)
);

INVxp67_ASAP7_75t_SL g1664 ( 
.A(n_1628),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1628),
.B(n_1593),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1635),
.B(n_1597),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1638),
.B(n_1598),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1643),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1629),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1629),
.Y(n_1670)
);

INVxp33_ASAP7_75t_L g1671 ( 
.A(n_1638),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1639),
.B(n_1602),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1639),
.B(n_1614),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1634),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1629),
.Y(n_1675)
);

AND2x2_ASAP7_75t_SL g1676 ( 
.A(n_1644),
.B(n_1564),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1631),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1628),
.B(n_1587),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1639),
.B(n_1622),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1644),
.B(n_1613),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1637),
.B(n_1607),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1631),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1644),
.A2(n_1609),
.B(n_1611),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1631),
.Y(n_1684)
);

INVx2_ASAP7_75t_SL g1685 ( 
.A(n_1634),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1634),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1634),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1641),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1622),
.B(n_1599),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1641),
.Y(n_1690)
);

OAI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1649),
.A2(n_1599),
.B1(n_1590),
.B2(n_1637),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1667),
.B(n_1637),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1660),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1660),
.B(n_1622),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1649),
.B(n_1644),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1650),
.B(n_1640),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1669),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1663),
.B(n_1640),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1669),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1689),
.B(n_1618),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1670),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1666),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1663),
.B(n_1640),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1689),
.B(n_1618),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1652),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1665),
.B(n_1616),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1652),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1666),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1681),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1683),
.B(n_1623),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1670),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1675),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1681),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1668),
.B(n_1623),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1651),
.B(n_1623),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1673),
.B(n_1625),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1655),
.B(n_1625),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1654),
.A2(n_1562),
.B1(n_1590),
.B2(n_1564),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1665),
.B(n_1616),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1655),
.B(n_1618),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1676),
.B(n_1625),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1676),
.B(n_1627),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1661),
.B(n_1582),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1675),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1662),
.B(n_1616),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1679),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1677),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1697),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1702),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1697),
.Y(n_1730)
);

OAI21xp33_ASAP7_75t_L g1731 ( 
.A1(n_1696),
.A2(n_1671),
.B(n_1676),
.Y(n_1731)
);

NOR2x1_ASAP7_75t_L g1732 ( 
.A(n_1691),
.B(n_1648),
.Y(n_1732)
);

AOI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1718),
.A2(n_1666),
.B1(n_1672),
.B2(n_1562),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1695),
.B(n_1664),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1723),
.B(n_1710),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1718),
.A2(n_1666),
.B1(n_1680),
.B2(n_1679),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1699),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1699),
.Y(n_1738)
);

AOI322xp5_ASAP7_75t_L g1739 ( 
.A1(n_1716),
.A2(n_1656),
.A3(n_1658),
.B1(n_1632),
.B2(n_1633),
.C1(n_1647),
.C2(n_1605),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1701),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1701),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1692),
.B(n_1521),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1711),
.Y(n_1743)
);

INVx1_ASAP7_75t_SL g1744 ( 
.A(n_1702),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_SL g1745 ( 
.A1(n_1708),
.A2(n_1698),
.B1(n_1703),
.B2(n_1656),
.Y(n_1745)
);

INVx2_ASAP7_75t_SL g1746 ( 
.A(n_1708),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1711),
.Y(n_1747)
);

NAND3xp33_ASAP7_75t_L g1748 ( 
.A(n_1709),
.B(n_1653),
.C(n_1648),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1712),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1712),
.Y(n_1750)
);

OAI322xp33_ASAP7_75t_L g1751 ( 
.A1(n_1726),
.A2(n_1658),
.A3(n_1653),
.B1(n_1678),
.B2(n_1685),
.C1(n_1677),
.C2(n_1684),
.Y(n_1751)
);

AOI21xp33_ASAP7_75t_L g1752 ( 
.A1(n_1705),
.A2(n_1678),
.B(n_1682),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1709),
.B(n_1682),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1724),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_SL g1755 ( 
.A(n_1732),
.B(n_1721),
.Y(n_1755)
);

AOI322xp5_ASAP7_75t_L g1756 ( 
.A1(n_1731),
.A2(n_1704),
.A3(n_1700),
.B1(n_1720),
.B2(n_1722),
.C1(n_1721),
.C2(n_1715),
.Y(n_1756)
);

OAI221xp5_ASAP7_75t_L g1757 ( 
.A1(n_1733),
.A2(n_1714),
.B1(n_1717),
.B2(n_1692),
.C(n_1726),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1736),
.A2(n_1704),
.B1(n_1700),
.B2(n_1720),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1728),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1746),
.B(n_1726),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1730),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1735),
.B(n_1709),
.Y(n_1762)
);

INVx1_ASAP7_75t_SL g1763 ( 
.A(n_1744),
.Y(n_1763)
);

A2O1A1Ixp33_ASAP7_75t_L g1764 ( 
.A1(n_1748),
.A2(n_1722),
.B(n_1713),
.C(n_1606),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1737),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1745),
.A2(n_1713),
.B(n_1707),
.Y(n_1766)
);

OAI222xp33_ASAP7_75t_L g1767 ( 
.A1(n_1744),
.A2(n_1693),
.B1(n_1713),
.B2(n_1725),
.C1(n_1685),
.C2(n_1694),
.Y(n_1767)
);

AOI21xp33_ASAP7_75t_SL g1768 ( 
.A1(n_1734),
.A2(n_1707),
.B(n_1705),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1738),
.Y(n_1769)
);

NAND4xp25_ASAP7_75t_SL g1770 ( 
.A(n_1739),
.B(n_1693),
.C(n_1725),
.D(n_1705),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1729),
.B(n_1742),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1753),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1740),
.B(n_1693),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1763),
.B(n_1741),
.Y(n_1774)
);

OAI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1755),
.A2(n_1752),
.B1(n_1753),
.B2(n_1707),
.C(n_1747),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1773),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1773),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_SL g1778 ( 
.A(n_1762),
.B(n_1751),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1760),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1758),
.A2(n_1694),
.B1(n_1754),
.B2(n_1750),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1762),
.B(n_1743),
.Y(n_1781)
);

OAI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1764),
.A2(n_1752),
.B(n_1749),
.Y(n_1782)
);

OAI221xp5_ASAP7_75t_L g1783 ( 
.A1(n_1764),
.A2(n_1719),
.B1(n_1706),
.B2(n_1727),
.C(n_1724),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1760),
.Y(n_1784)
);

NAND4xp25_ASAP7_75t_L g1785 ( 
.A(n_1778),
.B(n_1771),
.C(n_1780),
.D(n_1774),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_L g1786 ( 
.A(n_1782),
.B(n_1766),
.C(n_1768),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1779),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1784),
.B(n_1759),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1779),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1776),
.B(n_1772),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1777),
.B(n_1756),
.Y(n_1791)
);

NOR2xp67_ASAP7_75t_L g1792 ( 
.A(n_1775),
.B(n_1770),
.Y(n_1792)
);

OAI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1781),
.A2(n_1767),
.B(n_1757),
.Y(n_1793)
);

AOI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1786),
.A2(n_1793),
.B1(n_1785),
.B2(n_1791),
.C(n_1783),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1787),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1792),
.B(n_1761),
.Y(n_1796)
);

AOI211x1_ASAP7_75t_L g1797 ( 
.A1(n_1790),
.A2(n_1769),
.B(n_1765),
.C(n_1727),
.Y(n_1797)
);

AOI221xp5_ASAP7_75t_L g1798 ( 
.A1(n_1789),
.A2(n_1694),
.B1(n_1719),
.B2(n_1706),
.C(n_1687),
.Y(n_1798)
);

AOI221xp5_ASAP7_75t_L g1799 ( 
.A1(n_1794),
.A2(n_1788),
.B1(n_1694),
.B2(n_1686),
.C(n_1674),
.Y(n_1799)
);

AOI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1796),
.A2(n_1674),
.B1(n_1687),
.B2(n_1686),
.C(n_1657),
.Y(n_1800)
);

INVxp33_ASAP7_75t_SL g1801 ( 
.A(n_1795),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1797),
.Y(n_1802)
);

AOI222xp33_ASAP7_75t_L g1803 ( 
.A1(n_1798),
.A2(n_1620),
.B1(n_1615),
.B2(n_1605),
.C1(n_1606),
.C2(n_1627),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1795),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1799),
.A2(n_1659),
.B1(n_1657),
.B2(n_1684),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1804),
.Y(n_1806)
);

NAND3x1_ASAP7_75t_L g1807 ( 
.A(n_1802),
.B(n_1620),
.C(n_1688),
.Y(n_1807)
);

NOR3xp33_ASAP7_75t_SL g1808 ( 
.A(n_1801),
.B(n_1615),
.C(n_1554),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1803),
.B(n_1659),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1806),
.B(n_1800),
.Y(n_1810)
);

NAND3xp33_ASAP7_75t_L g1811 ( 
.A(n_1809),
.B(n_1527),
.C(n_1688),
.Y(n_1811)
);

NAND3xp33_ASAP7_75t_L g1812 ( 
.A(n_1808),
.B(n_1690),
.C(n_1620),
.Y(n_1812)
);

OAI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1812),
.A2(n_1807),
.B1(n_1805),
.B2(n_1690),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1813),
.A2(n_1810),
.B1(n_1811),
.B2(n_1606),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_SL g1815 ( 
.A1(n_1814),
.A2(n_1504),
.B1(n_1501),
.B2(n_1515),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1814),
.A2(n_1616),
.B1(n_1624),
.B2(n_1636),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_SL g1817 ( 
.A1(n_1815),
.A2(n_1504),
.B1(n_1498),
.B2(n_1496),
.Y(n_1817)
);

INVxp67_ASAP7_75t_L g1818 ( 
.A(n_1816),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1817),
.A2(n_1636),
.B1(n_1624),
.B2(n_1627),
.Y(n_1819)
);

AOI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1818),
.A2(n_1630),
.B1(n_1633),
.B2(n_1632),
.Y(n_1820)
);

AOI32xp33_ASAP7_75t_L g1821 ( 
.A1(n_1819),
.A2(n_1597),
.A3(n_1630),
.B1(n_1633),
.B2(n_1632),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1821),
.A2(n_1820),
.B1(n_1630),
.B2(n_1647),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1822),
.Y(n_1823)
);

AOI221xp5_ASAP7_75t_L g1824 ( 
.A1(n_1823),
.A2(n_1624),
.B1(n_1636),
.B2(n_1645),
.C(n_1641),
.Y(n_1824)
);

AOI211xp5_ASAP7_75t_L g1825 ( 
.A1(n_1824),
.A2(n_1496),
.B(n_1498),
.C(n_1636),
.Y(n_1825)
);


endmodule