module fake_ariane_472_n_790 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_790);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_790;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_166;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_56),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_46),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_42),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_8),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_69),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_5),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_16),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_117),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_20),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_49),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_148),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_86),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_79),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_3),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_5),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_12),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_13),
.Y(n_178)
);

BUFx2_ASAP7_75t_SL g179 ( 
.A(n_109),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_9),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_54),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_4),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_62),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_64),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_17),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_137),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_4),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_126),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_11),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_93),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_85),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_67),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_87),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_133),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_59),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_38),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_68),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_2),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_15),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_60),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_36),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_139),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_74),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_70),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_116),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_103),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_201),
.B(n_0),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_0),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g212 ( 
.A1(n_157),
.A2(n_1),
.B(n_2),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_159),
.B(n_1),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_178),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_216)
);

OA21x2_ASAP7_75t_L g217 ( 
.A1(n_160),
.A2(n_9),
.B(n_10),
.Y(n_217)
);

BUFx8_ASAP7_75t_SL g218 ( 
.A(n_183),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

AND2x4_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_10),
.Y(n_220)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_161),
.B(n_11),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_165),
.B(n_12),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_186),
.Y(n_229)
);

OA21x2_ASAP7_75t_L g230 ( 
.A1(n_168),
.A2(n_13),
.B(n_14),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

BUFx8_ASAP7_75t_SL g232 ( 
.A(n_163),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_164),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_170),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_174),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_176),
.A2(n_14),
.B1(n_18),
.B2(n_19),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_181),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_180),
.B(n_153),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

OAI21x1_ASAP7_75t_L g245 ( 
.A1(n_194),
.A2(n_21),
.B(n_22),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_196),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

AND2x6_ASAP7_75t_L g249 ( 
.A(n_203),
.B(n_23),
.Y(n_249)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_24),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_208),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_188),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_215),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_215),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_232),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_155),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_232),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_218),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_218),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_252),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_215),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_252),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_235),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_235),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_224),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_236),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_215),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_236),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_179),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_236),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_219),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_236),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_219),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_244),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_R g280 ( 
.A(n_247),
.B(n_156),
.Y(n_280)
);

NAND2xp33_ASAP7_75t_R g281 ( 
.A(n_212),
.B(n_158),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_240),
.B(n_162),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_244),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_251),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_247),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_247),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_248),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_248),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_211),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_211),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_210),
.Y(n_292)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_221),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_219),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_210),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_223),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_223),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_225),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_225),
.Y(n_299)
);

NAND2x1_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_249),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_243),
.Y(n_301)
);

NAND2xp33_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_249),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_227),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_269),
.Y(n_304)
);

AO221x1_ASAP7_75t_L g305 ( 
.A1(n_253),
.A2(n_214),
.B1(n_216),
.B2(n_238),
.C(n_209),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_276),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_227),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_285),
.B(n_243),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_263),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_266),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_256),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_257),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_276),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_291),
.B(n_280),
.Y(n_315)
);

NAND2xp33_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_249),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_231),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_265),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_284),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_231),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g322 ( 
.A(n_274),
.Y(n_322)
);

NOR3xp33_ASAP7_75t_L g323 ( 
.A(n_258),
.B(n_209),
.C(n_228),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_233),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_288),
.B(n_250),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_254),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_254),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_255),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_233),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_259),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_255),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_264),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_270),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_283),
.B(n_250),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_273),
.B(n_213),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_L g336 ( 
.A(n_279),
.B(n_221),
.C(n_220),
.Y(n_336)
);

NAND3xp33_ASAP7_75t_L g337 ( 
.A(n_275),
.B(n_221),
.C(n_220),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_277),
.B(n_234),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_271),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_264),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_272),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_272),
.B(n_234),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_278),
.B(n_242),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_267),
.B(n_220),
.Y(n_344)
);

NOR3xp33_ASAP7_75t_L g345 ( 
.A(n_260),
.B(n_239),
.C(n_238),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_278),
.B(n_242),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_268),
.B(n_238),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_294),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_261),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_294),
.B(n_249),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_271),
.B(n_241),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_271),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_262),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_271),
.B(n_249),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_281),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_292),
.B(n_249),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_290),
.B(n_212),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_285),
.B(n_166),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_290),
.B(n_212),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_253),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_285),
.B(n_167),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_269),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_322),
.A2(n_191),
.B1(n_171),
.B2(n_172),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_301),
.B(n_169),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_322),
.B(n_182),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_311),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_349),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_312),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_307),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_330),
.B(n_184),
.Y(n_371)
);

O2A1O1Ixp33_ASAP7_75t_L g372 ( 
.A1(n_361),
.A2(n_217),
.B(n_230),
.C(n_245),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_241),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_322),
.B(n_185),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_333),
.B(n_245),
.Y(n_375)
);

CKINVDCx11_ASAP7_75t_R g376 ( 
.A(n_304),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

AND2x6_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_229),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_322),
.B(n_187),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_306),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_358),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_322),
.B(n_189),
.Y(n_383)
);

AND2x6_ASAP7_75t_L g384 ( 
.A(n_360),
.B(n_229),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_342),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_322),
.B(n_192),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_335),
.B(n_202),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_327),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_342),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_303),
.B(n_206),
.Y(n_390)
);

NAND2x1p5_ASAP7_75t_L g391 ( 
.A(n_363),
.B(n_217),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_310),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_328),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_329),
.B(n_207),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_343),
.Y(n_395)
);

INVx5_ASAP7_75t_L g396 ( 
.A(n_339),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_314),
.Y(n_397)
);

BUFx8_ASAP7_75t_L g398 ( 
.A(n_347),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_331),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_309),
.B(n_217),
.Y(n_400)
);

OR2x6_ASAP7_75t_L g401 ( 
.A(n_315),
.B(n_230),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_L g402 ( 
.A1(n_336),
.A2(n_230),
.B1(n_241),
.B2(n_246),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_303),
.B(n_241),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_332),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_359),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_308),
.B(n_241),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_313),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_344),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_318),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_334),
.A2(n_229),
.B1(n_246),
.B2(n_27),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_308),
.B(n_246),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_340),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_339),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_323),
.B(n_305),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_341),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_317),
.B(n_246),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_329),
.A2(n_229),
.B1(n_246),
.B2(n_28),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_317),
.B(n_25),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_325),
.A2(n_337),
.B1(n_324),
.B2(n_321),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_321),
.Y(n_420)
);

NOR2x2_ASAP7_75t_L g421 ( 
.A(n_355),
.B(n_26),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_348),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_320),
.Y(n_423)
);

OR2x6_ASAP7_75t_L g424 ( 
.A(n_362),
.B(n_324),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_338),
.B(n_29),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_338),
.B(n_151),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_345),
.B(n_30),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_343),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_339),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_302),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_346),
.Y(n_431)
);

AND3x1_ASAP7_75t_SL g432 ( 
.A(n_346),
.B(n_34),
.C(n_35),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_376),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_356),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_387),
.A2(n_300),
.B1(n_354),
.B2(n_350),
.Y(n_435)
);

OAI21xp33_ASAP7_75t_L g436 ( 
.A1(n_371),
.A2(n_316),
.B(n_350),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_414),
.A2(n_352),
.B1(n_351),
.B2(n_40),
.Y(n_437)
);

O2A1O1Ixp33_ASAP7_75t_L g438 ( 
.A1(n_369),
.A2(n_352),
.B(n_39),
.C(n_41),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_419),
.B(n_392),
.Y(n_439)
);

AOI221xp5_ASAP7_75t_L g440 ( 
.A1(n_370),
.A2(n_381),
.B1(n_405),
.B2(n_408),
.C(n_427),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_374),
.A2(n_37),
.B(n_43),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_407),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_390),
.B(n_44),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_367),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_377),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_423),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_379),
.A2(n_45),
.B(n_47),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_429),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_368),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_396),
.Y(n_450)
);

INVx3_ASAP7_75t_SL g451 ( 
.A(n_421),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_366),
.A2(n_48),
.B(n_50),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_431),
.B(n_51),
.Y(n_453)
);

OAI21xp33_ASAP7_75t_L g454 ( 
.A1(n_365),
.A2(n_364),
.B(n_394),
.Y(n_454)
);

AO21x1_ASAP7_75t_L g455 ( 
.A1(n_418),
.A2(n_150),
.B(n_53),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_52),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_373),
.B(n_55),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_424),
.B(n_380),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_398),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_424),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_460)
);

INVx5_ASAP7_75t_L g461 ( 
.A(n_378),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_398),
.B(n_63),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_385),
.B(n_65),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_385),
.A2(n_66),
.B(n_71),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_380),
.B(n_72),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_409),
.B(n_73),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

AO32x2_ASAP7_75t_L g468 ( 
.A1(n_432),
.A2(n_75),
.A3(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_389),
.A2(n_80),
.B(n_81),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_382),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_396),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_383),
.A2(n_82),
.B(n_83),
.Y(n_472)
);

O2A1O1Ixp33_ASAP7_75t_L g473 ( 
.A1(n_389),
.A2(n_84),
.B(n_88),
.C(n_89),
.Y(n_473)
);

A2O1A1Ixp33_ASAP7_75t_L g474 ( 
.A1(n_395),
.A2(n_90),
.B(n_91),
.C(n_92),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_397),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_425),
.B(n_94),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_395),
.B(n_95),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_386),
.A2(n_96),
.B(n_97),
.Y(n_478)
);

OAI22x1_ASAP7_75t_L g479 ( 
.A1(n_375),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_397),
.Y(n_480)
);

OAI22x1_ASAP7_75t_L g481 ( 
.A1(n_375),
.A2(n_101),
.B1(n_102),
.B2(n_104),
.Y(n_481)
);

INVx3_ASAP7_75t_SL g482 ( 
.A(n_401),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_388),
.Y(n_483)
);

AND2x6_ASAP7_75t_L g484 ( 
.A(n_400),
.B(n_105),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_412),
.B(n_106),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_413),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_415),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_422),
.B(n_107),
.Y(n_488)
);

INVx5_ASAP7_75t_L g489 ( 
.A(n_378),
.Y(n_489)
);

NAND2x1p5_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_413),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_461),
.B(n_378),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_449),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_436),
.A2(n_426),
.B(n_372),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_448),
.Y(n_494)
);

AO21x2_ASAP7_75t_L g495 ( 
.A1(n_463),
.A2(n_402),
.B(n_416),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_461),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_451),
.Y(n_497)
);

AOI22x1_ASAP7_75t_L g498 ( 
.A1(n_441),
.A2(n_391),
.B1(n_393),
.B2(n_399),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_446),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_450),
.B(n_401),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_489),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_448),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_442),
.Y(n_503)
);

AOI22x1_ASAP7_75t_L g504 ( 
.A1(n_447),
.A2(n_404),
.B1(n_410),
.B2(n_411),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_489),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_489),
.Y(n_506)
);

NAND2x1p5_ASAP7_75t_L g507 ( 
.A(n_450),
.B(n_430),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_487),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_445),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_434),
.B(n_384),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_464),
.A2(n_406),
.B(n_403),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_439),
.B(n_384),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_444),
.Y(n_513)
);

AOI22x1_ASAP7_75t_L g514 ( 
.A1(n_479),
.A2(n_417),
.B1(n_384),
.B2(n_378),
.Y(n_514)
);

BUFx2_ASAP7_75t_SL g515 ( 
.A(n_433),
.Y(n_515)
);

AO21x2_ASAP7_75t_L g516 ( 
.A1(n_469),
.A2(n_384),
.B(n_110),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_470),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_467),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_483),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_467),
.B(n_111),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_485),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_471),
.Y(n_522)
);

AO21x2_ASAP7_75t_L g523 ( 
.A1(n_477),
.A2(n_112),
.B(n_113),
.Y(n_523)
);

AO21x2_ASAP7_75t_L g524 ( 
.A1(n_437),
.A2(n_114),
.B(n_115),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_440),
.B(n_118),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_458),
.B(n_119),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_488),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_444),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_466),
.B(n_121),
.Y(n_529)
);

BUFx10_ASAP7_75t_L g530 ( 
.A(n_471),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g531 ( 
.A1(n_455),
.A2(n_122),
.B(n_124),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_454),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_475),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_480),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_453),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_459),
.Y(n_536)
);

AO21x2_ASAP7_75t_L g537 ( 
.A1(n_456),
.A2(n_130),
.B(n_132),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_482),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_529),
.A2(n_460),
.B1(n_443),
.B2(n_465),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_529),
.A2(n_486),
.B1(n_462),
.B2(n_476),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_503),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_508),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_499),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_491),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_494),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_499),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_509),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_519),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_517),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_517),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_492),
.Y(n_551)
);

AOI21x1_ASAP7_75t_L g552 ( 
.A1(n_493),
.A2(n_457),
.B(n_435),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_501),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_533),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_494),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_534),
.Y(n_556)
);

BUFx10_ASAP7_75t_L g557 ( 
.A(n_497),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_500),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_521),
.B(n_484),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_491),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_502),
.B(n_513),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_491),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_500),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_530),
.Y(n_564)
);

NAND2x1p5_ASAP7_75t_L g565 ( 
.A(n_501),
.B(n_478),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_510),
.A2(n_481),
.B1(n_484),
.B2(n_474),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_502),
.B(n_468),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_530),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_501),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_500),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_521),
.A2(n_484),
.B1(n_472),
.B2(n_452),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_510),
.A2(n_468),
.B1(n_438),
.B2(n_473),
.Y(n_572)
);

CKINVDCx14_ASAP7_75t_R g573 ( 
.A(n_497),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_500),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_SL g575 ( 
.A1(n_514),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_527),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_513),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_522),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_522),
.Y(n_579)
);

BUFx2_ASAP7_75t_R g580 ( 
.A(n_515),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_527),
.A2(n_524),
.B1(n_535),
.B2(n_525),
.Y(n_581)
);

OR2x6_ASAP7_75t_L g582 ( 
.A(n_538),
.B(n_143),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_520),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_541),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_544),
.B(n_560),
.Y(n_585)
);

NOR3xp33_ASAP7_75t_SL g586 ( 
.A(n_540),
.B(n_526),
.C(n_512),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_567),
.B(n_507),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_551),
.B(n_528),
.Y(n_588)
);

NOR3xp33_ASAP7_75t_SL g589 ( 
.A(n_540),
.B(n_536),
.C(n_538),
.Y(n_589)
);

NOR3xp33_ASAP7_75t_SL g590 ( 
.A(n_539),
.B(n_538),
.C(n_530),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_545),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_551),
.B(n_554),
.Y(n_592)
);

NAND3xp33_ASAP7_75t_SL g593 ( 
.A(n_566),
.B(n_532),
.C(n_507),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_549),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_R g595 ( 
.A(n_573),
.B(n_538),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_557),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_539),
.A2(n_532),
.B(n_511),
.Y(n_597)
);

CKINVDCx16_ASAP7_75t_R g598 ( 
.A(n_557),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_555),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_561),
.B(n_518),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_577),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_580),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_544),
.B(n_560),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_550),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_562),
.B(n_518),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_562),
.B(n_518),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_558),
.B(n_506),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_542),
.B(n_506),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_563),
.B(n_506),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_547),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_583),
.B(n_501),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_564),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_570),
.B(n_505),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_548),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_553),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_556),
.B(n_579),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_578),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_553),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_553),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_568),
.B(n_505),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_574),
.B(n_520),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_569),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_543),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_546),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_581),
.A2(n_524),
.B1(n_559),
.B2(n_516),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_569),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_SL g627 ( 
.A1(n_582),
.A2(n_516),
.B1(n_531),
.B2(n_537),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_572),
.A2(n_511),
.B(n_531),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_582),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_580),
.B(n_496),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_559),
.Y(n_631)
);

NOR2x1_ASAP7_75t_L g632 ( 
.A(n_582),
.B(n_523),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_565),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_584),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_614),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_592),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_587),
.B(n_575),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_623),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_591),
.B(n_575),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_633),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_601),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_587),
.B(n_631),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_610),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_624),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_594),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_616),
.B(n_531),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_617),
.B(n_523),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_608),
.B(n_495),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_626),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_604),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_608),
.B(n_523),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_589),
.B(n_496),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_628),
.B(n_537),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_628),
.B(n_537),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_599),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_588),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_593),
.B(n_565),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_621),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_600),
.B(n_490),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_597),
.B(n_552),
.Y(n_660)
);

AO22x1_ASAP7_75t_L g661 ( 
.A1(n_632),
.A2(n_571),
.B1(n_576),
.B2(n_490),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_607),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_597),
.B(n_144),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_632),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_586),
.B(n_145),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_613),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_627),
.A2(n_504),
.B1(n_498),
.B2(n_149),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_622),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_590),
.B(n_585),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_585),
.B(n_146),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_613),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_603),
.B(n_618),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_634),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_SL g674 ( 
.A1(n_665),
.A2(n_630),
.B(n_625),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_649),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_645),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_634),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_656),
.B(n_636),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_642),
.B(n_598),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_635),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_645),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_640),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_663),
.B(n_639),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_641),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_647),
.B(n_618),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_642),
.B(n_612),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_647),
.B(n_603),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_642),
.B(n_622),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_660),
.B(n_615),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_641),
.B(n_615),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_660),
.B(n_615),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_646),
.B(n_607),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_646),
.B(n_609),
.Y(n_693)
);

NAND2x1p5_ASAP7_75t_L g694 ( 
.A(n_652),
.B(n_619),
.Y(n_694)
);

AND2x2_ASAP7_75t_SL g695 ( 
.A(n_663),
.B(n_629),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_643),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_638),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_650),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_638),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_641),
.B(n_620),
.Y(n_700)
);

AOI21xp33_ASAP7_75t_SL g701 ( 
.A1(n_665),
.A2(n_596),
.B(n_602),
.Y(n_701)
);

AND2x2_ASAP7_75t_SL g702 ( 
.A(n_653),
.B(n_629),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_651),
.B(n_619),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_651),
.B(n_605),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_666),
.B(n_605),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_703),
.B(n_654),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_703),
.B(n_654),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_675),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_673),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_682),
.B(n_662),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_678),
.B(n_685),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_692),
.B(n_653),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_683),
.B(n_640),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_689),
.B(n_671),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_676),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_677),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_685),
.B(n_648),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_692),
.B(n_672),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_676),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_681),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_687),
.B(n_648),
.Y(n_721)
);

BUFx2_ASAP7_75t_SL g722 ( 
.A(n_684),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_680),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_687),
.B(n_658),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_717),
.B(n_686),
.Y(n_725)
);

NAND4xp75_ASAP7_75t_SL g726 ( 
.A(n_722),
.B(n_701),
.C(n_669),
.D(n_689),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_715),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_709),
.B(n_683),
.Y(n_728)
);

NOR3xp33_ASAP7_75t_L g729 ( 
.A(n_713),
.B(n_674),
.C(n_700),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_715),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_710),
.A2(n_695),
.B(n_661),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_708),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_706),
.B(n_691),
.Y(n_733)
);

AOI33xp33_ASAP7_75t_L g734 ( 
.A1(n_723),
.A2(n_691),
.A3(n_693),
.B1(n_696),
.B2(n_684),
.B3(n_637),
.Y(n_734)
);

AOI221xp5_ASAP7_75t_L g735 ( 
.A1(n_716),
.A2(n_637),
.B1(n_667),
.B2(n_661),
.C(n_693),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_721),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_719),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_736),
.B(n_711),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_728),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_729),
.B(n_706),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_728),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_735),
.A2(n_695),
.B1(n_702),
.B2(n_669),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_727),
.Y(n_743)
);

XOR2x2_ASAP7_75t_L g744 ( 
.A(n_726),
.B(n_702),
.Y(n_744)
);

AOI322xp5_ASAP7_75t_L g745 ( 
.A1(n_742),
.A2(n_735),
.A3(n_707),
.B1(n_712),
.B2(n_734),
.C1(n_733),
.C2(n_732),
.Y(n_745)
);

OAI222xp33_ASAP7_75t_L g746 ( 
.A1(n_742),
.A2(n_731),
.B1(n_679),
.B2(n_725),
.C1(n_724),
.C2(n_737),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_740),
.A2(n_688),
.B1(n_712),
.B2(n_707),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_739),
.Y(n_748)
);

OAI221xp5_ASAP7_75t_L g749 ( 
.A1(n_741),
.A2(n_730),
.B1(n_694),
.B2(n_657),
.C(n_719),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_748),
.Y(n_750)
);

NAND2xp33_ASAP7_75t_L g751 ( 
.A(n_747),
.B(n_595),
.Y(n_751)
);

NOR3x1_ASAP7_75t_L g752 ( 
.A(n_749),
.B(n_744),
.C(n_690),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_745),
.B(n_738),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_750),
.B(n_718),
.Y(n_754)
);

OAI21xp33_ASAP7_75t_L g755 ( 
.A1(n_753),
.A2(n_655),
.B(n_718),
.Y(n_755)
);

OAI211xp5_ASAP7_75t_SL g756 ( 
.A1(n_751),
.A2(n_746),
.B(n_668),
.C(n_655),
.Y(n_756)
);

OAI211xp5_ASAP7_75t_SL g757 ( 
.A1(n_755),
.A2(n_752),
.B(n_668),
.C(n_743),
.Y(n_757)
);

O2A1O1Ixp5_ASAP7_75t_L g758 ( 
.A1(n_754),
.A2(n_668),
.B(n_670),
.C(n_652),
.Y(n_758)
);

NOR3xp33_ASAP7_75t_L g759 ( 
.A(n_756),
.B(n_670),
.C(n_657),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_757),
.Y(n_760)
);

NOR2x1_ASAP7_75t_L g761 ( 
.A(n_758),
.B(n_759),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_758),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_758),
.Y(n_763)
);

NOR2x1_ASAP7_75t_L g764 ( 
.A(n_757),
.B(n_652),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_762),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_764),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_763),
.B(n_714),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_761),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_760),
.Y(n_769)
);

OAI221xp5_ASAP7_75t_L g770 ( 
.A1(n_762),
.A2(n_694),
.B1(n_664),
.B2(n_659),
.C(n_720),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_768),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_769),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_767),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_765),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_766),
.Y(n_775)
);

OA22x2_ASAP7_75t_L g776 ( 
.A1(n_775),
.A2(n_770),
.B1(n_672),
.B2(n_714),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_772),
.Y(n_777)
);

OAI21x1_ASAP7_75t_L g778 ( 
.A1(n_771),
.A2(n_611),
.B(n_704),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_775),
.B(n_606),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_773),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_780),
.A2(n_774),
.B1(n_714),
.B2(n_664),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_777),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_779),
.Y(n_783)
);

XNOR2xp5_ASAP7_75t_L g784 ( 
.A(n_782),
.B(n_776),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_783),
.A2(n_778),
.B1(n_606),
.B2(n_720),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_SL g786 ( 
.A1(n_784),
.A2(n_781),
.B1(n_705),
.B2(n_671),
.Y(n_786)
);

AOI21x1_ASAP7_75t_L g787 ( 
.A1(n_786),
.A2(n_785),
.B(n_704),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_787),
.A2(n_699),
.B1(n_697),
.B2(n_644),
.Y(n_788)
);

OR2x6_ASAP7_75t_L g789 ( 
.A(n_788),
.B(n_705),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_789),
.A2(n_650),
.B1(n_644),
.B2(n_698),
.Y(n_790)
);


endmodule