module fake_jpeg_23234_n_343 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_1),
.B(n_4),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_0),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_53),
.B(n_63),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_60),
.Y(n_82)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_47),
.B(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_39),
.B(n_26),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_35),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_37),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_69),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_42),
.A2(n_26),
.B1(n_20),
.B2(n_23),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_77),
.B1(n_23),
.B2(n_20),
.Y(n_108)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_36),
.A2(n_17),
.B1(n_21),
.B2(n_33),
.Y(n_77)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_34),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_84),
.A2(n_112),
.B(n_21),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_40),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_104),
.Y(n_121)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_19),
.B1(n_40),
.B2(n_36),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_61),
.B1(n_58),
.B2(n_55),
.Y(n_119)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_92),
.Y(n_138)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_99),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_15),
.C(n_9),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_101),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_57),
.A2(n_19),
.B(n_54),
.C(n_76),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_102),
.B1(n_109),
.B2(n_91),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_54),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_100),
.Y(n_141)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_19),
.B1(n_48),
.B2(n_44),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_30),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_103),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_28),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_28),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_28),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_24),
.B1(n_22),
.B2(n_18),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_50),
.A2(n_23),
.B1(n_20),
.B2(n_32),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g112 ( 
.A1(n_74),
.A2(n_46),
.B(n_35),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_28),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_66),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

AOI32xp33_ASAP7_75t_L g115 ( 
.A1(n_51),
.A2(n_48),
.A3(n_46),
.B1(n_44),
.B2(n_41),
.Y(n_115)
);

AOI32xp33_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_49),
.A3(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_116),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_17),
.B(n_33),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_135),
.B(n_78),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_119),
.A2(n_125),
.B1(n_126),
.B2(n_140),
.Y(n_173)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_142),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_95),
.A2(n_55),
.B1(n_17),
.B2(n_21),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_84),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_132),
.Y(n_148)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_84),
.B(n_41),
.CI(n_44),
.CON(n_131),
.SN(n_131)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_131),
.B(n_113),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_75),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_41),
.C(n_56),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_144),
.C(n_114),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_49),
.B1(n_32),
.B2(n_31),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_146),
.B1(n_30),
.B2(n_81),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_90),
.A2(n_31),
.B1(n_16),
.B2(n_24),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_81),
.B1(n_111),
.B2(n_92),
.Y(n_161)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_101),
.Y(n_147)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_79),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_94),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_104),
.B(n_25),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_147),
.B(n_150),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_121),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_162),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_152),
.A2(n_165),
.B(n_168),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_153),
.B(n_128),
.C(n_117),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_87),
.B1(n_102),
.B2(n_80),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_172),
.B1(n_177),
.B2(n_179),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_163),
.B(n_166),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_107),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_156),
.B(n_127),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_158),
.B(n_174),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_160),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_90),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_102),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_105),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_169),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_132),
.B(n_131),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_118),
.A2(n_136),
.B(n_145),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_167),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_126),
.B(n_80),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_110),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_170),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

AOI22x1_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_102),
.B1(n_106),
.B2(n_25),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_141),
.B(n_87),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_175),
.B(n_176),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_144),
.Y(n_176)
);

NAND2x1_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_103),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_129),
.B(n_127),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_141),
.B(n_22),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_180),
.B(n_18),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_178),
.A2(n_134),
.B1(n_133),
.B2(n_140),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_181),
.A2(n_196),
.B1(n_197),
.B2(n_205),
.Y(n_215)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_188),
.Y(n_217)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_178),
.A2(n_119),
.B1(n_144),
.B2(n_139),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_189),
.A2(n_148),
.B1(n_163),
.B2(n_154),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_16),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_192),
.A2(n_198),
.B(n_0),
.Y(n_234)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_195),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_93),
.B1(n_94),
.B2(n_129),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_93),
.B1(n_128),
.B2(n_117),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_199),
.B(n_206),
.Y(n_218)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_204),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_14),
.Y(n_232)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_173),
.A2(n_172),
.B1(n_176),
.B2(n_165),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_166),
.B(n_99),
.Y(n_206)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_211),
.C(n_152),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_153),
.B(n_98),
.C(n_18),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_150),
.B(n_16),
.Y(n_212)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_148),
.A2(n_98),
.B1(n_1),
.B2(n_2),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_214),
.A2(n_177),
.B1(n_175),
.B2(n_158),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_195),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_207),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_219),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_225),
.C(n_238),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_235),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

BUFx4f_ASAP7_75t_SL g249 ( 
.A(n_222),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_186),
.A2(n_155),
.B(n_163),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_224),
.A2(n_234),
.B(n_183),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_156),
.C(n_168),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_151),
.B1(n_174),
.B2(n_180),
.Y(n_226)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_230),
.B(n_233),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_181),
.A2(n_151),
.B1(n_170),
.B2(n_171),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_237),
.B1(n_206),
.B2(n_183),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_197),
.Y(n_259)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_185),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_182),
.B(n_14),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_2),
.C(n_3),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_9),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_241),
.C(n_211),
.Y(n_253)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_240),
.B(n_242),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_2),
.C(n_5),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_184),
.Y(n_244)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_263),
.Y(n_267)
);

O2A1O1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_190),
.B(n_198),
.C(n_214),
.Y(n_250)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_251),
.A2(n_254),
.B1(n_266),
.B2(n_210),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_184),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_252),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_253),
.B(n_192),
.Y(n_281)
);

INVxp33_ASAP7_75t_L g255 ( 
.A(n_217),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_264),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_204),
.C(n_186),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_225),
.C(n_239),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_246),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_261),
.B(n_265),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_224),
.A2(n_190),
.B(n_194),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_234),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_228),
.B(n_193),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g264 ( 
.A(n_229),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_191),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_231),
.A2(n_189),
.B1(n_200),
.B2(n_187),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_271),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_257),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_278),
.C(n_279),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_260),
.A2(n_200),
.B1(n_221),
.B2(n_237),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_275),
.A2(n_276),
.B1(n_285),
.B2(n_266),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_215),
.B1(n_235),
.B2(n_191),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_280),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_238),
.C(n_215),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_232),
.C(n_207),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_216),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_281),
.A2(n_252),
.B(n_244),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_254),
.B(n_192),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_282),
.B(n_259),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_253),
.B1(n_256),
.B2(n_243),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_250),
.A2(n_241),
.B1(n_213),
.B2(n_199),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_212),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_286),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_289),
.B(n_293),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_245),
.Y(n_290)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

XNOR2x1_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_261),
.Y(n_291)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_297),
.C(n_301),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_188),
.Y(n_292)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_292),
.Y(n_316)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_299),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_298),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_248),
.Y(n_299)
);

AO21x1_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_272),
.B(n_282),
.Y(n_300)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_300),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_249),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_256),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_279),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_291),
.A2(n_249),
.B1(n_274),
.B2(n_276),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_303),
.A2(n_313),
.B1(n_288),
.B2(n_7),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_269),
.Y(n_304)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_304),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_301),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_307),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_278),
.C(n_273),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_308),
.A2(n_312),
.B(n_6),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_10),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_249),
.C(n_7),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_299),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_297),
.B(n_294),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_317),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_307),
.A2(n_294),
.B(n_288),
.Y(n_319)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_320),
.A2(n_322),
.B1(n_11),
.B2(n_12),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_306),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_325),
.C(n_326),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_312),
.A2(n_10),
.B(n_11),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_12),
.C(n_13),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_11),
.Y(n_326)
);

AOI322xp5_ASAP7_75t_L g329 ( 
.A1(n_318),
.A2(n_310),
.A3(n_304),
.B1(n_314),
.B2(n_305),
.C1(n_309),
.C2(n_315),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_330),
.C(n_13),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_321),
.A2(n_316),
.B1(n_314),
.B2(n_305),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_331),
.A2(n_12),
.B(n_13),
.C(n_8),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_8),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_317),
.B(n_322),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_335),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_336),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_338),
.B(n_328),
.Y(n_340)
);

INVxp33_ASAP7_75t_L g341 ( 
.A(n_340),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_339),
.B(n_327),
.C(n_337),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_329),
.Y(n_343)
);


endmodule