module fake_jpeg_9759_n_277 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_24),
.Y(n_51)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_18),
.B1(n_21),
.B2(n_27),
.Y(n_68)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_47),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_R g96 ( 
.A(n_53),
.B(n_24),
.Y(n_96)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_56),
.Y(n_92)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_62),
.Y(n_106)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_23),
.B1(n_31),
.B2(n_30),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_65),
.A2(n_41),
.B1(n_40),
.B2(n_36),
.Y(n_103)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_66),
.B(n_29),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_19),
.B1(n_34),
.B2(n_31),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_67),
.A2(n_70),
.B1(n_44),
.B2(n_41),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_21),
.B1(n_18),
.B2(n_27),
.Y(n_83)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_69),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_75),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_30),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_73),
.B(n_80),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_33),
.B1(n_32),
.B2(n_35),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_83),
.B1(n_87),
.B2(n_89),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_17),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_22),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_82),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_70),
.A2(n_36),
.B(n_40),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g132 ( 
.A(n_84),
.Y(n_132)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_85),
.A2(n_94),
.B1(n_41),
.B2(n_40),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_48),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_104),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_33),
.B1(n_32),
.B2(n_24),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_55),
.A2(n_35),
.B1(n_24),
.B2(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_90),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_91),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_39),
.B1(n_37),
.B2(n_45),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_93),
.A2(n_98),
.B1(n_28),
.B2(n_26),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_36),
.Y(n_116)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_17),
.B1(n_20),
.B2(n_39),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_52),
.B(n_20),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_39),
.Y(n_102)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_124),
.B1(n_135),
.B2(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_113),
.B(n_125),
.Y(n_164)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_118),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_116),
.B(n_26),
.Y(n_156)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_84),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_133),
.Y(n_153)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_106),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_148),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_SL g138 ( 
.A1(n_116),
.A2(n_82),
.B(n_96),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_138),
.A2(n_139),
.B1(n_25),
.B2(n_118),
.Y(n_186)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_147),
.Y(n_170)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_79),
.C(n_81),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_142),
.B(n_149),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_127),
.A2(n_79),
.B1(n_100),
.B2(n_95),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_119),
.B1(n_125),
.B2(n_113),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_130),
.B1(n_108),
.B2(n_111),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_105),
.B1(n_95),
.B2(n_99),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_122),
.B1(n_117),
.B2(n_128),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_100),
.C(n_42),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_29),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_121),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_29),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_157),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_42),
.C(n_77),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_154),
.Y(n_188)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_155),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_115),
.Y(n_177)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_29),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_159),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_25),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_0),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_161),
.A2(n_157),
.B(n_148),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_85),
.B1(n_78),
.B2(n_72),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_163),
.A2(n_107),
.B1(n_72),
.B2(n_78),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_169),
.A2(n_183),
.B(n_185),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_174),
.B1(n_179),
.B2(n_161),
.Y(n_194)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_175),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_108),
.B1(n_111),
.B2(n_110),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_186),
.Y(n_203)
);

AO22x1_ASAP7_75t_SL g179 ( 
.A1(n_147),
.A2(n_110),
.B1(n_26),
.B2(n_88),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_180),
.B(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_107),
.B1(n_90),
.B2(n_114),
.Y(n_182)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

NOR2xp67_ASAP7_75t_SL g185 ( 
.A(n_151),
.B(n_131),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_160),
.B(n_42),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_159),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_190),
.B(n_3),
.Y(n_202)
);

NAND3xp33_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_158),
.C(n_137),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_202),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_150),
.C(n_146),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_195),
.C(n_197),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_204),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_156),
.C(n_140),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_145),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_136),
.C(n_155),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_201),
.C(n_172),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_187),
.Y(n_200)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_136),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_186),
.B1(n_165),
.B2(n_175),
.Y(n_221)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_173),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_121),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_209),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_162),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_210),
.A2(n_165),
.B1(n_183),
.B2(n_171),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_3),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_211),
.Y(n_217)
);

AO21x1_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_178),
.B(n_179),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_224),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_219),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_199),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_177),
.C(n_184),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_220),
.A2(n_221),
.B1(n_225),
.B2(n_194),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_167),
.C(n_42),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_198),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_196),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_210),
.A2(n_167),
.B1(n_5),
.B2(n_7),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_42),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_SL g229 ( 
.A(n_226),
.B(n_228),
.C(n_197),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_42),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_237),
.Y(n_248)
);

BUFx12_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_231),
.B(n_235),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_208),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_240),
.Y(n_251)
);

OAI321xp33_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_205),
.A3(n_201),
.B1(n_209),
.B2(n_206),
.C(n_193),
.Y(n_234)
);

NAND4xp25_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_227),
.C(n_214),
.D(n_228),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

XNOR2x1_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_206),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_225),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_242),
.Y(n_244)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_240),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_212),
.C(n_222),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_211),
.B(n_5),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_247),
.C(n_250),
.Y(n_254)
);

XOR2x1_ASAP7_75t_SL g258 ( 
.A(n_246),
.B(n_42),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_216),
.C(n_219),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_232),
.C(n_223),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_4),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_235),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_253),
.B(n_5),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_230),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_243),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_238),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_257),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_4),
.Y(n_257)
);

NAND3xp33_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_244),
.C(n_7),
.Y(n_262)
);

OAI221xp5_ASAP7_75t_L g264 ( 
.A1(n_259),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_254),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_252),
.C(n_244),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_263),
.Y(n_268)
);

OAI21x1_ASAP7_75t_SL g269 ( 
.A1(n_262),
.A2(n_264),
.B(n_8),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_266),
.A2(n_267),
.B(n_269),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_262),
.A2(n_258),
.B(n_255),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_268),
.A2(n_265),
.B(n_10),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_272),
.Y(n_273)
);

A2O1A1O1Ixp25_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_8),
.B(n_11),
.C(n_12),
.D(n_13),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_271),
.A2(n_13),
.B(n_14),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_15),
.C(n_16),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_273),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_15),
.Y(n_277)
);


endmodule