module fake_ibex_167_n_787 (n_85, n_128, n_84, n_64, n_3, n_73, n_65, n_103, n_95, n_55, n_130, n_63, n_98, n_129, n_29, n_106, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_88, n_133, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_50, n_11, n_92, n_101, n_113, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_91, n_54, n_19, n_787);

input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_103;
input n_95;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_106;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_133;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_50;
input n_11;
input n_92;
input n_101;
input n_113;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_787;

wire n_151;
wire n_599;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_738;
wire n_475;
wire n_166;
wire n_163;
wire n_753;
wire n_747;
wire n_500;
wire n_645;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_187;
wire n_667;
wire n_154;
wire n_682;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_723;
wire n_170;
wire n_144;
wire n_270;
wire n_383;
wire n_346;
wire n_561;
wire n_417;
wire n_471;
wire n_739;
wire n_755;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_598;
wire n_143;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_355;
wire n_767;
wire n_474;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_141;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_689;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_139;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_772;
wire n_768;
wire n_338;
wire n_173;
wire n_696;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_718;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_546;
wire n_199;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_138;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_332;
wire n_517;
wire n_211;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_164;
wire n_616;
wire n_782;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_728;
wire n_670;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_752;
wire n_668;
wire n_779;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_149;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_159;
wire n_231;
wire n_298;
wire n_202;
wire n_587;
wire n_760;
wire n_751;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_82),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_27),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_45),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_50),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_56),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_18),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_28),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_47),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_75),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_70),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_127),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_18),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_7),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_107),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_62),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_43),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_69),
.Y(n_159)
);

NOR2xp67_ASAP7_75t_L g160 ( 
.A(n_103),
.B(n_89),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_120),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_14),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_51),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_19),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_131),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_29),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_37),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_98),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_2),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_2),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_119),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_115),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_0),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_15),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_83),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_12),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_99),
.Y(n_187)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_97),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_29),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_38),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_72),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_25),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_90),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_100),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_L g196 ( 
.A(n_111),
.B(n_84),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_36),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_30),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_73),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_110),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_118),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_38),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_79),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_1),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_10),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_94),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_78),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_117),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_59),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_129),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_74),
.Y(n_213)
);

BUFx8_ASAP7_75t_SL g214 ( 
.A(n_71),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_86),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_46),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_22),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_11),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_48),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_77),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_122),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_87),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_124),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_114),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_39),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_123),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_95),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_130),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_76),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_49),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_67),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_66),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_40),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_39),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_0),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g236 ( 
.A(n_151),
.B(n_1),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_154),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_151),
.Y(n_238)
);

CKINVDCx6p67_ASAP7_75t_R g239 ( 
.A(n_143),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_146),
.B(n_174),
.Y(n_241)
);

CKINVDCx11_ASAP7_75t_R g242 ( 
.A(n_197),
.Y(n_242)
);

AND2x6_ASAP7_75t_L g243 ( 
.A(n_176),
.B(n_41),
.Y(n_243)
);

OAI21x1_ASAP7_75t_L g244 ( 
.A1(n_176),
.A2(n_68),
.B(n_135),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_188),
.B(n_3),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_201),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_188),
.B(n_4),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_180),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_154),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_169),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_169),
.Y(n_253)
);

BUFx8_ASAP7_75t_L g254 ( 
.A(n_180),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_156),
.B(n_4),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_197),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_256)
);

CKINVDCx11_ASAP7_75t_R g257 ( 
.A(n_199),
.Y(n_257)
);

AND2x4_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_5),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_169),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_180),
.Y(n_260)
);

BUFx8_ASAP7_75t_L g261 ( 
.A(n_180),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_215),
.B(n_8),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_185),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g264 ( 
.A(n_142),
.B(n_9),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_180),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_147),
.B(n_9),
.Y(n_266)
);

CKINVDCx11_ASAP7_75t_R g267 ( 
.A(n_199),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_140),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_203),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_224),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g271 ( 
.A(n_138),
.B(n_42),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_162),
.Y(n_272)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_185),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_198),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_180),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_149),
.B(n_13),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_198),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_148),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_163),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_163),
.Y(n_280)
);

OA21x2_ASAP7_75t_L g281 ( 
.A1(n_170),
.A2(n_80),
.B(n_134),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_172),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_175),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_185),
.B(n_16),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_210),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_178),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_155),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_198),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_142),
.B(n_173),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_165),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_210),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_170),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_198),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_166),
.B(n_17),
.Y(n_294)
);

NAND2xp33_ASAP7_75t_L g295 ( 
.A(n_192),
.B(n_44),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_173),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_171),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_184),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_186),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_200),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_200),
.Y(n_301)
);

BUFx8_ASAP7_75t_L g302 ( 
.A(n_231),
.Y(n_302)
);

AND2x4_ASAP7_75t_L g303 ( 
.A(n_179),
.B(n_20),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_157),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_189),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_L g306 ( 
.A(n_243),
.B(n_219),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_271),
.A2(n_203),
.B1(n_209),
.B2(n_181),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_236),
.Y(n_308)
);

NAND3xp33_ASAP7_75t_L g309 ( 
.A(n_245),
.B(n_206),
.C(n_183),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_254),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_236),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_258),
.A2(n_234),
.B1(n_190),
.B2(n_205),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_268),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_249),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_273),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_263),
.B(n_204),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_L g318 ( 
.A1(n_239),
.A2(n_195),
.B1(n_181),
.B2(n_209),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_258),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_243),
.Y(n_320)
);

AND2x2_ASAP7_75t_SL g321 ( 
.A(n_271),
.B(n_264),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_254),
.B(n_231),
.Y(n_322)
);

AND2x6_ASAP7_75t_L g323 ( 
.A(n_264),
.B(n_179),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_250),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_237),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_261),
.Y(n_327)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_285),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g329 ( 
.A(n_241),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_261),
.B(n_144),
.Y(n_330)
);

AND2x4_ASAP7_75t_L g331 ( 
.A(n_285),
.B(n_291),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_145),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_265),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_237),
.Y(n_334)
);

OR2x6_ASAP7_75t_L g335 ( 
.A(n_256),
.B(n_214),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_245),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_242),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_242),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_257),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_275),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_248),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_278),
.B(n_225),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_275),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_303),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_238),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_251),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_251),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_257),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_287),
.B(n_212),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_253),
.Y(n_350)
);

BUFx4f_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_253),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_240),
.B(n_139),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_259),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_259),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_303),
.B(n_152),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_289),
.B(n_141),
.Y(n_357)
);

AND2x6_ASAP7_75t_L g358 ( 
.A(n_284),
.B(n_212),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_290),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_247),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_279),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_279),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_252),
.A2(n_192),
.B1(n_164),
.B2(n_167),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_302),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_280),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_274),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_274),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_277),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_243),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_277),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_288),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_292),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_288),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_297),
.B(n_272),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_288),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_325),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_321),
.A2(n_262),
.B1(n_255),
.B2(n_284),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_364),
.B(n_302),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_255),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_321),
.A2(n_304),
.B1(n_235),
.B2(n_305),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_329),
.B(n_336),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_334),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_307),
.A2(n_283),
.B1(n_282),
.B2(n_299),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_374),
.A2(n_294),
.B1(n_276),
.B2(n_296),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_341),
.A2(n_243),
.B1(n_286),
.B2(n_298),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_331),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_266),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_345),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_331),
.Y(n_389)
);

NAND3xp33_ASAP7_75t_L g390 ( 
.A(n_309),
.B(n_294),
.C(n_270),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_313),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_306),
.A2(n_295),
.B(n_281),
.Y(n_392)
);

BUFx12f_ASAP7_75t_L g393 ( 
.A(n_337),
.Y(n_393)
);

INVx8_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_360),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_361),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_324),
.A2(n_269),
.B1(n_246),
.B2(n_300),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_310),
.B(n_244),
.Y(n_398)
);

A2O1A1Ixp33_ASAP7_75t_L g399 ( 
.A1(n_308),
.A2(n_301),
.B(n_300),
.C(n_244),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_362),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_317),
.B(n_150),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_349),
.B(n_153),
.Y(n_403)
);

AND2x4_ASAP7_75t_SL g404 ( 
.A(n_342),
.B(n_267),
.Y(n_404)
);

OR2x6_ASAP7_75t_L g405 ( 
.A(n_335),
.B(n_301),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_320),
.B(n_158),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_327),
.A2(n_182),
.B1(n_187),
.B2(n_191),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_312),
.A2(n_207),
.B1(n_208),
.B2(n_211),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_328),
.B(n_159),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_315),
.B(n_232),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_312),
.A2(n_220),
.B1(n_213),
.B2(n_216),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_332),
.B(n_161),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_332),
.B(n_168),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_323),
.A2(n_281),
.B1(n_193),
.B2(n_194),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_372),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_353),
.B(n_177),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_337),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_357),
.B(n_202),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_319),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_351),
.B(n_223),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_318),
.B(n_338),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_311),
.B(n_316),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_369),
.B(n_330),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_330),
.B(n_221),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_356),
.B(n_226),
.Y(n_425)
);

AO22x1_ASAP7_75t_L g426 ( 
.A1(n_339),
.A2(n_228),
.B1(n_233),
.B2(n_227),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_344),
.B(n_160),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_322),
.B(n_196),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_363),
.Y(n_430)
);

OR2x6_ASAP7_75t_L g431 ( 
.A(n_335),
.B(n_229),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g432 ( 
.A1(n_323),
.A2(n_293),
.B1(n_288),
.B2(n_24),
.Y(n_432)
);

OAI22xp33_ASAP7_75t_L g433 ( 
.A1(n_335),
.A2(n_293),
.B1(n_23),
.B2(n_24),
.Y(n_433)
);

INVx8_ASAP7_75t_L g434 ( 
.A(n_358),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_322),
.B(n_21),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_339),
.B(n_25),
.Y(n_436)
);

AND2x6_ASAP7_75t_L g437 ( 
.A(n_314),
.B(n_137),
.Y(n_437)
);

AO21x1_ASAP7_75t_L g438 ( 
.A1(n_398),
.A2(n_435),
.B(n_429),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_391),
.B(n_348),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_423),
.A2(n_422),
.B(n_399),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_387),
.B(n_348),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_381),
.B(n_326),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_381),
.B(n_333),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_414),
.A2(n_340),
.B(n_343),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_377),
.A2(n_340),
.B1(n_343),
.B2(n_371),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_26),
.Y(n_446)
);

O2A1O1Ixp33_ASAP7_75t_L g447 ( 
.A1(n_408),
.A2(n_411),
.B(n_383),
.C(n_380),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_383),
.A2(n_375),
.B1(n_373),
.B2(n_371),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_431),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_428),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_385),
.A2(n_354),
.B(n_346),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_390),
.B(n_30),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_394),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_386),
.B(n_31),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_389),
.B(n_31),
.Y(n_455)
);

O2A1O1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_408),
.A2(n_367),
.B(n_350),
.C(n_352),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_419),
.Y(n_457)
);

INVx3_ASAP7_75t_SL g458 ( 
.A(n_417),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_431),
.Y(n_459)
);

INVxp33_ASAP7_75t_SL g460 ( 
.A(n_421),
.Y(n_460)
);

AND2x2_ASAP7_75t_SL g461 ( 
.A(n_404),
.B(n_32),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_394),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_430),
.A2(n_355),
.B1(n_350),
.B2(n_366),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_403),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_382),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_434),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_393),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_384),
.B(n_33),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_405),
.B(n_33),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_378),
.B(n_34),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_396),
.B(n_400),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_411),
.B(n_34),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_434),
.Y(n_473)
);

BUFx2_ASAP7_75t_SL g474 ( 
.A(n_436),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_401),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_405),
.B(n_35),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_376),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_424),
.B(n_35),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_405),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_416),
.B(n_407),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_397),
.A2(n_370),
.B1(n_368),
.B2(n_347),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_415),
.B(n_36),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_426),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_388),
.Y(n_484)
);

BUFx12f_ASAP7_75t_L g485 ( 
.A(n_437),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_395),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_425),
.B(n_52),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_406),
.A2(n_53),
.B(n_54),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_427),
.B(n_55),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_412),
.A2(n_57),
.B(n_58),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_437),
.Y(n_491)
);

AO21x1_ASAP7_75t_L g492 ( 
.A1(n_433),
.A2(n_60),
.B(n_61),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_418),
.B(n_63),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_437),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_413),
.A2(n_64),
.B(n_65),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_410),
.B(n_402),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_420),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_409),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_453),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_453),
.Y(n_500)
);

A2O1A1Ixp33_ASAP7_75t_L g501 ( 
.A1(n_447),
.A2(n_496),
.B(n_480),
.C(n_452),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_486),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_464),
.B(n_432),
.Y(n_503)
);

NOR2x1_ASAP7_75t_L g504 ( 
.A(n_467),
.B(n_88),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_484),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_461),
.B(n_441),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_465),
.Y(n_507)
);

OA22x2_ASAP7_75t_L g508 ( 
.A1(n_479),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_458),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_462),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_442),
.B(n_443),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_460),
.B(n_102),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_473),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_473),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_457),
.B(n_497),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_477),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_466),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_482),
.Y(n_518)
);

AO31x2_ASAP7_75t_L g519 ( 
.A1(n_448),
.A2(n_133),
.A3(n_438),
.B(n_492),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_466),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_470),
.B(n_483),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_498),
.B(n_474),
.Y(n_522)
);

A2O1A1Ixp33_ASAP7_75t_L g523 ( 
.A1(n_487),
.A2(n_456),
.B(n_493),
.C(n_478),
.Y(n_523)
);

AO31x2_ASAP7_75t_L g524 ( 
.A1(n_445),
.A2(n_463),
.A3(n_495),
.B(n_490),
.Y(n_524)
);

A2O1A1Ixp33_ASAP7_75t_L g525 ( 
.A1(n_489),
.A2(n_455),
.B(n_454),
.C(n_450),
.Y(n_525)
);

AOI221x1_ASAP7_75t_L g526 ( 
.A1(n_494),
.A2(n_488),
.B1(n_446),
.B2(n_451),
.C(n_469),
.Y(n_526)
);

OAI22x1_ASAP7_75t_L g527 ( 
.A1(n_476),
.A2(n_449),
.B1(n_439),
.B2(n_459),
.Y(n_527)
);

BUFx8_ASAP7_75t_SL g528 ( 
.A(n_485),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_486),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_480),
.B(n_329),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_480),
.B(n_329),
.Y(n_531)
);

NAND3xp33_ASAP7_75t_SL g532 ( 
.A(n_447),
.B(n_338),
.C(n_337),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_480),
.B(n_329),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_440),
.A2(n_399),
.B(n_444),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_480),
.B(n_329),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_480),
.B(n_329),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_464),
.B(n_329),
.Y(n_537)
);

AOI221x1_ASAP7_75t_L g538 ( 
.A1(n_481),
.A2(n_440),
.B1(n_448),
.B2(n_452),
.C(n_399),
.Y(n_538)
);

AOI211x1_ASAP7_75t_L g539 ( 
.A1(n_468),
.A2(n_383),
.B(n_472),
.C(n_433),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_460),
.A2(n_307),
.B1(n_461),
.B2(n_269),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_453),
.B(n_462),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_480),
.B(n_329),
.Y(n_542)
);

OA21x2_ASAP7_75t_L g543 ( 
.A1(n_440),
.A2(n_399),
.B(n_392),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_475),
.Y(n_544)
);

A2O1A1Ixp33_ASAP7_75t_L g545 ( 
.A1(n_447),
.A2(n_496),
.B(n_480),
.C(n_452),
.Y(n_545)
);

AOI221x1_ASAP7_75t_L g546 ( 
.A1(n_481),
.A2(n_440),
.B1(n_448),
.B2(n_452),
.C(n_399),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_480),
.B(n_329),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_475),
.Y(n_548)
);

OAI21xp33_ASAP7_75t_SL g549 ( 
.A1(n_471),
.A2(n_321),
.B(n_271),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_440),
.A2(n_399),
.B(n_392),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_480),
.A2(n_321),
.B1(n_383),
.B2(n_460),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_SL g552 ( 
.A1(n_447),
.A2(n_307),
.B(n_383),
.Y(n_552)
);

OAI21x1_ASAP7_75t_SL g553 ( 
.A1(n_491),
.A2(n_447),
.B(n_471),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_480),
.B(n_329),
.Y(n_554)
);

BUFx12f_ASAP7_75t_L g555 ( 
.A(n_467),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_453),
.B(n_462),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_511),
.A2(n_525),
.B(n_523),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_543),
.Y(n_558)
);

AO21x2_ASAP7_75t_L g559 ( 
.A1(n_553),
.A2(n_550),
.B(n_534),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_502),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_530),
.B(n_531),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_509),
.Y(n_562)
);

OA21x2_ASAP7_75t_L g563 ( 
.A1(n_538),
.A2(n_546),
.B(n_550),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_537),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_533),
.B(n_535),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_549),
.A2(n_545),
.B(n_501),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_507),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_510),
.Y(n_568)
);

CKINVDCx11_ASAP7_75t_R g569 ( 
.A(n_555),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_529),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_516),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_536),
.B(n_542),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_517),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_547),
.B(n_554),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_522),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_505),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_506),
.B(n_551),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_513),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_544),
.Y(n_579)
);

BUFx12f_ASAP7_75t_L g580 ( 
.A(n_521),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_548),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_515),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_521),
.B(n_532),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_514),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_540),
.B(n_518),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_540),
.B(n_541),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_500),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_524),
.Y(n_588)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_508),
.A2(n_504),
.B(n_520),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g590 ( 
.A1(n_520),
.A2(n_514),
.B(n_519),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_503),
.B(n_556),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_499),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_539),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_528),
.Y(n_594)
);

CKINVDCx8_ASAP7_75t_R g595 ( 
.A(n_512),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_527),
.A2(n_511),
.B(n_525),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_511),
.A2(n_525),
.B(n_523),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_502),
.Y(n_598)
);

OA21x2_ASAP7_75t_L g599 ( 
.A1(n_538),
.A2(n_546),
.B(n_550),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_509),
.Y(n_600)
);

AO21x2_ASAP7_75t_L g601 ( 
.A1(n_553),
.A2(n_550),
.B(n_534),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_511),
.A2(n_525),
.B(n_523),
.Y(n_602)
);

OA21x2_ASAP7_75t_L g603 ( 
.A1(n_538),
.A2(n_546),
.B(n_550),
.Y(n_603)
);

OA21x2_ASAP7_75t_L g604 ( 
.A1(n_538),
.A2(n_546),
.B(n_550),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_502),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_502),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_509),
.Y(n_607)
);

AO31x2_ASAP7_75t_L g608 ( 
.A1(n_538),
.A2(n_546),
.A3(n_526),
.B(n_545),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_511),
.A2(n_525),
.B(n_523),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_543),
.Y(n_610)
);

CKINVDCx6p67_ASAP7_75t_R g611 ( 
.A(n_555),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_549),
.A2(n_545),
.B(n_501),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g613 ( 
.A1(n_549),
.A2(n_545),
.B(n_501),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_537),
.B(n_379),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_502),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_511),
.A2(n_525),
.B(n_523),
.Y(n_616)
);

A2O1A1Ixp33_ASAP7_75t_L g617 ( 
.A1(n_501),
.A2(n_545),
.B(n_549),
.C(n_552),
.Y(n_617)
);

NOR2x1_ASAP7_75t_SL g618 ( 
.A(n_511),
.B(n_453),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_593),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_614),
.B(n_561),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_587),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_558),
.Y(n_622)
);

CKINVDCx6p67_ASAP7_75t_R g623 ( 
.A(n_611),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_566),
.B(n_612),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_569),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_592),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_585),
.B(n_586),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_572),
.B(n_574),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_573),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_576),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_573),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_569),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_575),
.B(n_577),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_573),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_579),
.Y(n_635)
);

OR2x6_ASAP7_75t_L g636 ( 
.A(n_586),
.B(n_589),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_617),
.B(n_582),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_617),
.B(n_565),
.Y(n_638)
);

BUFx12f_ASAP7_75t_L g639 ( 
.A(n_562),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_568),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_571),
.B(n_613),
.Y(n_641)
);

BUFx12f_ASAP7_75t_L g642 ( 
.A(n_562),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_557),
.A2(n_616),
.B(n_609),
.Y(n_643)
);

OR2x6_ASAP7_75t_L g644 ( 
.A(n_586),
.B(n_589),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_581),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_560),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_L g647 ( 
.A1(n_597),
.A2(n_602),
.B(n_596),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_567),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_570),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_610),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_598),
.B(n_615),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_605),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_606),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_585),
.B(n_564),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_580),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_591),
.A2(n_583),
.B1(n_580),
.B2(n_607),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_618),
.B(n_590),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_578),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_595),
.B(n_584),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_559),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_563),
.B(n_604),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_563),
.B(n_604),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_629),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_622),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_629),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_631),
.Y(n_666)
);

INVxp67_ASAP7_75t_SL g667 ( 
.A(n_621),
.Y(n_667)
);

OAI211xp5_ASAP7_75t_L g668 ( 
.A1(n_656),
.A2(n_594),
.B(n_604),
.C(n_603),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_624),
.B(n_601),
.Y(n_669)
);

AND2x4_ASAP7_75t_SL g670 ( 
.A(n_623),
.B(n_594),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_624),
.B(n_563),
.Y(n_671)
);

HB1xp67_ASAP7_75t_SL g672 ( 
.A(n_625),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_630),
.A2(n_621),
.B1(n_638),
.B2(n_634),
.Y(n_673)
);

OR2x6_ASAP7_75t_L g674 ( 
.A(n_636),
.B(n_588),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_657),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_634),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_628),
.B(n_600),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_633),
.B(n_638),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_650),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_633),
.B(n_599),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_641),
.B(n_599),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_623),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_641),
.B(n_608),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_652),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_651),
.B(n_608),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_651),
.B(n_608),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_684),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_682),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_679),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_678),
.B(n_637),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_678),
.B(n_637),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_675),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_664),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_675),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_680),
.B(n_661),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_685),
.B(n_660),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_686),
.B(n_661),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_670),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_667),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_686),
.B(n_662),
.Y(n_700)
);

NAND2x1_ASAP7_75t_L g701 ( 
.A(n_666),
.B(n_644),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_665),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_671),
.B(n_662),
.Y(n_703)
);

OR2x6_ASAP7_75t_L g704 ( 
.A(n_701),
.B(n_674),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_689),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_702),
.Y(n_706)
);

AND2x4_ASAP7_75t_SL g707 ( 
.A(n_702),
.B(n_666),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_697),
.B(n_700),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_687),
.B(n_683),
.Y(n_709)
);

NOR2x1p5_ASAP7_75t_L g710 ( 
.A(n_701),
.B(n_666),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_697),
.B(n_669),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_693),
.Y(n_712)
);

NAND4xp25_ASAP7_75t_L g713 ( 
.A(n_690),
.B(n_627),
.C(n_668),
.D(n_654),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_695),
.B(n_680),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_703),
.B(n_669),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_691),
.B(n_699),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_703),
.B(n_681),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_692),
.Y(n_718)
);

NOR2x1_ASAP7_75t_L g719 ( 
.A(n_698),
.B(n_665),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_719),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_705),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_714),
.B(n_708),
.Y(n_722)
);

NAND2x1p5_ASAP7_75t_L g723 ( 
.A(n_710),
.B(n_666),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_705),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_719),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_708),
.B(n_717),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_717),
.B(n_696),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_714),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_712),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_709),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_716),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_704),
.B(n_692),
.Y(n_732)
);

OAI211xp5_ASAP7_75t_L g733 ( 
.A1(n_713),
.A2(n_694),
.B(n_688),
.C(n_626),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_726),
.B(n_728),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_729),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_726),
.B(n_711),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_727),
.B(n_715),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_730),
.B(n_731),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_722),
.Y(n_739)
);

OAI22xp33_ASAP7_75t_L g740 ( 
.A1(n_723),
.A2(n_704),
.B1(n_694),
.B2(n_673),
.Y(n_740)
);

INVx1_ASAP7_75t_SL g741 ( 
.A(n_722),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_721),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_721),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_724),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_727),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_733),
.A2(n_718),
.B1(n_644),
.B2(n_711),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_741),
.B(n_715),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_738),
.Y(n_748)
);

AOI21xp33_ASAP7_75t_L g749 ( 
.A1(n_740),
.A2(n_725),
.B(n_720),
.Y(n_749)
);

OAI222xp33_ASAP7_75t_L g750 ( 
.A1(n_746),
.A2(n_723),
.B1(n_725),
.B2(n_720),
.C1(n_732),
.C2(n_704),
.Y(n_750)
);

OAI211xp5_ASAP7_75t_SL g751 ( 
.A1(n_740),
.A2(n_677),
.B(n_659),
.C(n_626),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_742),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_739),
.A2(n_732),
.B1(n_718),
.B2(n_704),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_753),
.A2(n_723),
.B1(n_736),
.B2(n_745),
.Y(n_754)
);

OAI221xp5_ASAP7_75t_SL g755 ( 
.A1(n_748),
.A2(n_704),
.B1(n_640),
.B2(n_734),
.C(n_644),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_752),
.B(n_737),
.Y(n_756)
);

NAND3xp33_ASAP7_75t_L g757 ( 
.A(n_755),
.B(n_749),
.C(n_751),
.Y(n_757)
);

AOI211xp5_ASAP7_75t_L g758 ( 
.A1(n_754),
.A2(n_751),
.B(n_750),
.C(n_625),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_757),
.B(n_632),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_758),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_760),
.A2(n_756),
.B1(n_747),
.B2(n_672),
.Y(n_761)
);

NOR2xp67_ASAP7_75t_L g762 ( 
.A(n_759),
.B(n_632),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_761),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_762),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_763),
.B(n_737),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_764),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_764),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_766),
.Y(n_768)
);

XOR2xp5_ASAP7_75t_L g769 ( 
.A(n_767),
.B(n_600),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_SL g770 ( 
.A1(n_765),
.A2(n_642),
.B1(n_639),
.B2(n_640),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_766),
.A2(n_655),
.B(n_642),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_766),
.A2(n_655),
.B(n_639),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_768),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_769),
.Y(n_774)
);

OAI21x1_ASAP7_75t_L g775 ( 
.A1(n_771),
.A2(n_620),
.B(n_710),
.Y(n_775)
);

XOR2x2_ASAP7_75t_L g776 ( 
.A(n_772),
.B(n_732),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_SL g777 ( 
.A(n_770),
.B(n_643),
.C(n_635),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_769),
.A2(n_645),
.B(n_744),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_774),
.A2(n_663),
.B(n_653),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_773),
.A2(n_649),
.B(n_646),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_776),
.B(n_743),
.Y(n_781)
);

AOI222xp33_ASAP7_75t_L g782 ( 
.A1(n_777),
.A2(n_648),
.B1(n_735),
.B2(n_706),
.C1(n_665),
.C2(n_619),
.Y(n_782)
);

O2A1O1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_779),
.A2(n_778),
.B(n_775),
.C(n_663),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_781),
.A2(n_706),
.B1(n_735),
.B2(n_676),
.Y(n_784)
);

AO21x2_ASAP7_75t_L g785 ( 
.A1(n_780),
.A2(n_647),
.B(n_658),
.Y(n_785)
);

OAI21xp5_ASAP7_75t_SL g786 ( 
.A1(n_783),
.A2(n_782),
.B(n_707),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_786),
.A2(n_784),
.B(n_785),
.Y(n_787)
);


endmodule