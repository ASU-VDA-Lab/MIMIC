module real_aes_18011_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_835, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_835;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_756;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
AND2x4_ASAP7_75t_L g795 ( .A(n_0), .B(n_796), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_1), .A2(n_4), .B1(n_137), .B2(n_477), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g179 ( .A1(n_2), .A2(n_42), .B1(n_144), .B2(n_180), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_3), .A2(n_24), .B1(n_180), .B2(n_222), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_5), .A2(n_16), .B1(n_134), .B2(n_211), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_6), .A2(n_61), .B1(n_194), .B2(n_224), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_7), .A2(n_17), .B1(n_144), .B2(n_165), .Y(n_580) );
INVx1_ASAP7_75t_L g796 ( .A(n_8), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_9), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_10), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_11), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_12), .A2(n_18), .B1(n_193), .B2(n_196), .Y(n_192) );
OR2x2_ASAP7_75t_L g788 ( .A(n_13), .B(n_38), .Y(n_788) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_14), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_15), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_19), .A2(n_100), .B1(n_134), .B2(n_137), .Y(n_133) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_20), .A2(n_37), .B1(n_169), .B2(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_21), .B(n_135), .Y(n_166) );
OAI21x1_ASAP7_75t_L g152 ( .A1(n_22), .A2(n_57), .B(n_153), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_23), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_25), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_26), .B(n_141), .Y(n_500) );
INVx4_ASAP7_75t_R g548 ( .A(n_27), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_28), .A2(n_47), .B1(n_182), .B2(n_183), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_29), .A2(n_54), .B1(n_134), .B2(n_183), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_30), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_31), .B(n_169), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_32), .Y(n_245) );
INVx1_ASAP7_75t_L g479 ( .A(n_33), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_34), .B(n_180), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_SL g491 ( .A1(n_35), .A2(n_140), .B(n_144), .C(n_492), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_36), .A2(n_55), .B1(n_144), .B2(n_183), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_39), .A2(n_87), .B1(n_144), .B2(n_221), .Y(n_220) );
XOR2x2_ASAP7_75t_L g105 ( .A(n_40), .B(n_106), .Y(n_105) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_41), .A2(n_46), .B1(n_144), .B2(n_165), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_43), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_44), .A2(n_59), .B1(n_134), .B2(n_143), .Y(n_142) );
AOI22xp5_ASAP7_75t_L g106 ( .A1(n_45), .A2(n_72), .B1(n_107), .B2(n_108), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_45), .Y(n_108) );
INVx1_ASAP7_75t_L g503 ( .A(n_48), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_49), .B(n_144), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_50), .Y(n_520) );
INVx2_ASAP7_75t_L g794 ( .A(n_51), .Y(n_794) );
BUFx3_ASAP7_75t_L g787 ( .A(n_52), .Y(n_787) );
INVx1_ASAP7_75t_L g808 ( .A(n_52), .Y(n_808) );
OAI21xp5_ASAP7_75t_L g797 ( .A1(n_53), .A2(n_798), .B(n_810), .Y(n_797) );
AOI31xp33_ASAP7_75t_L g810 ( .A1(n_53), .A2(n_811), .A3(n_813), .B(n_814), .Y(n_810) );
INVx2_ASAP7_75t_L g833 ( .A(n_53), .Y(n_833) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_56), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_58), .A2(n_88), .B1(n_144), .B2(n_183), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_60), .A2(n_68), .B1(n_801), .B2(n_802), .Y(n_800) );
INVx1_ASAP7_75t_L g802 ( .A(n_60), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_62), .A2(n_76), .B1(n_143), .B2(n_182), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_63), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_64), .A2(n_78), .B1(n_144), .B2(n_165), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_65), .A2(n_99), .B1(n_134), .B2(n_196), .Y(n_242) );
AND2x4_ASAP7_75t_L g130 ( .A(n_66), .B(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g153 ( .A(n_67), .Y(n_153) );
INVx1_ASAP7_75t_L g801 ( .A(n_68), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_69), .A2(n_91), .B1(n_182), .B2(n_183), .Y(n_475) );
AO22x1_ASAP7_75t_L g537 ( .A1(n_70), .A2(n_77), .B1(n_208), .B2(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g131 ( .A(n_71), .Y(n_131) );
INVx1_ASAP7_75t_L g107 ( .A(n_72), .Y(n_107) );
AND2x2_ASAP7_75t_L g495 ( .A(n_73), .B(n_175), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_74), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_75), .B(n_224), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_79), .B(n_180), .Y(n_521) );
INVx2_ASAP7_75t_L g141 ( .A(n_80), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_81), .B(n_175), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_82), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_83), .A2(n_98), .B1(n_183), .B2(n_224), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_84), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_85), .B(n_151), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_86), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_89), .Y(n_815) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_90), .B(n_175), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_92), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_93), .B(n_175), .Y(n_517) );
INVx1_ASAP7_75t_L g116 ( .A(n_94), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_94), .B(n_807), .Y(n_806) );
NAND2xp33_ASAP7_75t_L g171 ( .A(n_95), .B(n_135), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_96), .A2(n_199), .B(n_224), .C(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g550 ( .A(n_97), .B(n_551), .Y(n_550) );
NAND2xp33_ASAP7_75t_L g525 ( .A(n_101), .B(n_170), .Y(n_525) );
AOI221xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_782), .B1(n_797), .B2(n_818), .C(n_822), .Y(n_102) );
AOI22xp33_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_105), .B1(n_109), .B2(n_781), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g781 ( .A(n_109), .Y(n_781) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OAI22xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_117), .B1(n_457), .B2(n_458), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_114), .Y(n_457) );
BUFx8_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g790 ( .A(n_115), .B(n_786), .Y(n_790) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
XOR2xp5_ASAP7_75t_L g799 ( .A(n_118), .B(n_800), .Y(n_799) );
OR2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_360), .Y(n_118) );
NAND4xp25_ASAP7_75t_L g119 ( .A(n_120), .B(n_284), .C(n_315), .D(n_344), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_251), .Y(n_120) );
OAI322xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_187), .A3(n_216), .B1(n_229), .B2(n_237), .C1(n_246), .C2(n_248), .Y(n_121) );
INVxp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_123), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_157), .Y(n_123) );
AND2x2_ASAP7_75t_L g281 ( .A(n_124), .B(n_282), .Y(n_281) );
INVx4_ASAP7_75t_L g317 ( .A(n_124), .Y(n_317) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g292 ( .A(n_125), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g295 ( .A(n_125), .B(n_189), .Y(n_295) );
AND2x2_ASAP7_75t_L g312 ( .A(n_125), .B(n_205), .Y(n_312) );
AND2x2_ASAP7_75t_L g410 ( .A(n_125), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g233 ( .A(n_126), .Y(n_233) );
AND2x4_ASAP7_75t_L g416 ( .A(n_126), .B(n_411), .Y(n_416) );
AO31x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_132), .A3(n_148), .B(n_154), .Y(n_126) );
AO31x2_ASAP7_75t_L g240 ( .A1(n_127), .A2(n_200), .A3(n_241), .B(n_244), .Y(n_240) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_128), .A2(n_543), .B(n_546), .Y(n_542) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AO31x2_ASAP7_75t_L g177 ( .A1(n_129), .A2(n_178), .A3(n_184), .B(n_185), .Y(n_177) );
AO31x2_ASAP7_75t_L g190 ( .A1(n_129), .A2(n_191), .A3(n_200), .B(n_202), .Y(n_190) );
AO31x2_ASAP7_75t_L g205 ( .A1(n_129), .A2(n_206), .A3(n_213), .B(n_214), .Y(n_205) );
AO31x2_ASAP7_75t_L g578 ( .A1(n_129), .A2(n_156), .A3(n_579), .B(n_582), .Y(n_578) );
BUFx10_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
BUFx10_ASAP7_75t_L g470 ( .A(n_130), .Y(n_470) );
INVx1_ASAP7_75t_L g494 ( .A(n_130), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_139), .B1(n_142), .B2(n_145), .Y(n_132) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVxp67_ASAP7_75t_SL g538 ( .A(n_135), .Y(n_538) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g138 ( .A(n_136), .Y(n_138) );
INVx3_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_136), .Y(n_170) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_136), .Y(n_180) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_136), .Y(n_183) );
INVx1_ASAP7_75t_L g195 ( .A(n_136), .Y(n_195) );
INVx1_ASAP7_75t_L g209 ( .A(n_136), .Y(n_209) );
INVx1_ASAP7_75t_L g212 ( .A(n_136), .Y(n_212) );
INVx2_ASAP7_75t_L g222 ( .A(n_136), .Y(n_222) );
INVx1_ASAP7_75t_L g224 ( .A(n_136), .Y(n_224) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_138), .B(n_488), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_139), .A2(n_168), .B(n_171), .Y(n_167) );
OAI22xp5_ASAP7_75t_L g178 ( .A1(n_139), .A2(n_145), .B1(n_179), .B2(n_181), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_139), .A2(n_192), .B1(n_197), .B2(n_198), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_139), .A2(n_145), .B1(n_207), .B2(n_210), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_139), .A2(n_220), .B1(n_223), .B2(n_225), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_139), .A2(n_198), .B1(n_242), .B2(n_243), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_139), .A2(n_145), .B1(n_261), .B2(n_262), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_139), .A2(n_467), .B1(n_468), .B2(n_469), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_139), .A2(n_225), .B1(n_475), .B2(n_476), .Y(n_474) );
OAI22x1_ASAP7_75t_L g579 ( .A1(n_139), .A2(n_225), .B1(n_580), .B2(n_581), .Y(n_579) );
INVx6_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
O2A1O1Ixp5_ASAP7_75t_L g163 ( .A1(n_140), .A2(n_164), .B(n_165), .C(n_166), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_140), .A2(n_525), .B(n_526), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_140), .B(n_537), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g594 ( .A1(n_140), .A2(n_533), .B(n_537), .C(n_540), .Y(n_594) );
BUFx8_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
INVx1_ASAP7_75t_L g199 ( .A(n_141), .Y(n_199) );
INVx1_ASAP7_75t_L g490 ( .A(n_141), .Y(n_490) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx4_ASAP7_75t_L g165 ( .A(n_144), .Y(n_165) );
INVx1_ASAP7_75t_L g196 ( .A(n_144), .Y(n_196) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g469 ( .A(n_146), .Y(n_469) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g523 ( .A(n_147), .Y(n_523) );
AO31x2_ASAP7_75t_L g259 ( .A1(n_148), .A2(n_226), .A3(n_260), .B(n_263), .Y(n_259) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_148), .A2(n_542), .B(n_550), .Y(n_541) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_SL g202 ( .A(n_150), .B(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_150), .B(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g156 ( .A(n_151), .Y(n_156) );
INVx2_ASAP7_75t_L g201 ( .A(n_151), .Y(n_201) );
OAI21xp33_ASAP7_75t_L g540 ( .A1(n_151), .A2(n_494), .B(n_535), .Y(n_540) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_152), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_156), .B(n_264), .Y(n_263) );
AND2x4_ASAP7_75t_L g421 ( .A(n_157), .B(n_322), .Y(n_421) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g250 ( .A(n_158), .Y(n_250) );
INVxp67_ASAP7_75t_SL g408 ( .A(n_158), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_176), .Y(n_158) );
AND2x2_ASAP7_75t_L g238 ( .A(n_159), .B(n_177), .Y(n_238) );
INVx1_ASAP7_75t_L g279 ( .A(n_159), .Y(n_279) );
OAI21x1_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_162), .B(n_174), .Y(n_159) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_160), .A2(n_162), .B(n_174), .Y(n_274) );
INVx2_ASAP7_75t_SL g160 ( .A(n_161), .Y(n_160) );
INVx4_ASAP7_75t_L g175 ( .A(n_161), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_161), .B(n_186), .Y(n_185) );
BUFx3_ASAP7_75t_L g213 ( .A(n_161), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_161), .B(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_161), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g507 ( .A(n_161), .B(n_470), .Y(n_507) );
OAI21x1_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_167), .B(n_172), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_165), .A2(n_520), .B(n_521), .C(n_522), .Y(n_519) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g182 ( .A(n_170), .Y(n_182) );
OAI22xp33_ASAP7_75t_L g547 ( .A1(n_170), .A2(n_212), .B1(n_548), .B2(n_549), .Y(n_547) );
INVx2_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_SL g226 ( .A(n_173), .Y(n_226) );
INVx2_ASAP7_75t_L g184 ( .A(n_175), .Y(n_184) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_175), .B(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g270 ( .A(n_176), .Y(n_270) );
AND2x2_ASAP7_75t_L g334 ( .A(n_176), .B(n_273), .Y(n_334) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g288 ( .A(n_177), .Y(n_288) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_177), .Y(n_341) );
OR2x2_ASAP7_75t_L g412 ( .A(n_177), .B(n_218), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_180), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g477 ( .A(n_183), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_183), .B(n_502), .Y(n_501) );
AO31x2_ASAP7_75t_L g465 ( .A1(n_184), .A2(n_466), .A3(n_470), .B(n_471), .Y(n_465) );
NAND4xp25_ASAP7_75t_L g290 ( .A(n_187), .B(n_291), .C(n_294), .D(n_296), .Y(n_290) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g428 ( .A(n_188), .B(n_416), .Y(n_428) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_204), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_189), .B(n_257), .Y(n_256) );
AND2x4_ASAP7_75t_L g282 ( .A(n_189), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g302 ( .A(n_189), .Y(n_302) );
INVx1_ASAP7_75t_L g319 ( .A(n_189), .Y(n_319) );
INVx1_ASAP7_75t_L g327 ( .A(n_189), .Y(n_327) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_189), .Y(n_441) );
INVx4_ASAP7_75t_SL g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_190), .B(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g359 ( .A(n_190), .B(n_259), .Y(n_359) );
AND2x2_ASAP7_75t_L g367 ( .A(n_190), .B(n_205), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_190), .B(n_390), .Y(n_389) );
BUFx2_ASAP7_75t_L g432 ( .A(n_190), .Y(n_432) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_195), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g225 ( .A(n_199), .Y(n_225) );
AO31x2_ASAP7_75t_L g473 ( .A1(n_200), .A2(n_226), .A3(n_474), .B(n_478), .Y(n_473) );
AOI21x1_ASAP7_75t_L g482 ( .A1(n_200), .A2(n_483), .B(n_495), .Y(n_482) );
BUFx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_201), .B(n_472), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_201), .B(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g551 ( .A(n_201), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_201), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g236 ( .A(n_205), .Y(n_236) );
OR2x2_ASAP7_75t_L g297 ( .A(n_205), .B(n_259), .Y(n_297) );
INVx2_ASAP7_75t_L g304 ( .A(n_205), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_205), .B(n_257), .Y(n_328) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_205), .Y(n_415) );
OAI21xp33_ASAP7_75t_SL g499 ( .A1(n_208), .A2(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AO31x2_ASAP7_75t_L g218 ( .A1(n_213), .A2(n_219), .A3(n_226), .B(n_227), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_216), .B(n_387), .Y(n_386) );
BUFx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g239 ( .A(n_218), .B(n_240), .Y(n_239) );
BUFx2_ASAP7_75t_L g249 ( .A(n_218), .Y(n_249) );
INVx2_ASAP7_75t_L g267 ( .A(n_218), .Y(n_267) );
AND2x4_ASAP7_75t_L g299 ( .A(n_218), .B(n_271), .Y(n_299) );
OR2x2_ASAP7_75t_L g379 ( .A(n_218), .B(n_279), .Y(n_379) );
INVx2_ASAP7_75t_SL g221 ( .A(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_222), .B(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_225), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_234), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_231), .B(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g296 ( .A(n_231), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_231), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_232), .B(n_302), .Y(n_310) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g255 ( .A(n_233), .Y(n_255) );
OR2x2_ASAP7_75t_L g348 ( .A(n_233), .B(n_258), .Y(n_348) );
INVx1_ASAP7_75t_L g275 ( .A(n_234), .Y(n_275) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g247 ( .A(n_235), .Y(n_247) );
INVx1_ASAP7_75t_L g283 ( .A(n_236), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
OAI322xp33_ASAP7_75t_L g251 ( .A1(n_238), .A2(n_252), .A3(n_265), .B1(n_268), .B2(n_275), .C1(n_276), .C2(n_280), .Y(n_251) );
AND2x4_ASAP7_75t_L g298 ( .A(n_238), .B(n_299), .Y(n_298) );
AOI211xp5_ASAP7_75t_SL g329 ( .A1(n_238), .A2(n_330), .B(n_331), .C(n_335), .Y(n_329) );
AND2x2_ASAP7_75t_L g349 ( .A(n_238), .B(n_239), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_238), .B(n_266), .Y(n_355) );
AND2x4_ASAP7_75t_SL g277 ( .A(n_239), .B(n_278), .Y(n_277) );
NAND3xp33_ASAP7_75t_L g368 ( .A(n_239), .B(n_295), .C(n_323), .Y(n_368) );
AND2x2_ASAP7_75t_L g399 ( .A(n_239), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g266 ( .A(n_240), .B(n_267), .Y(n_266) );
INVx3_ASAP7_75t_L g271 ( .A(n_240), .Y(n_271) );
BUFx2_ASAP7_75t_L g339 ( .A(n_240), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_249), .B(n_273), .Y(n_272) );
NAND2x1_ASAP7_75t_L g313 ( .A(n_249), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g332 ( .A(n_249), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_250), .B(n_266), .Y(n_397) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_256), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g340 ( .A(n_255), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_259), .Y(n_293) );
AND2x4_ASAP7_75t_L g303 ( .A(n_259), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g390 ( .A(n_259), .Y(n_390) );
INVx2_ASAP7_75t_L g411 ( .A(n_259), .Y(n_411) );
OAI22xp33_ASAP7_75t_L g423 ( .A1(n_265), .A2(n_424), .B1(n_426), .B2(n_427), .Y(n_423) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g335 ( .A(n_266), .B(n_336), .Y(n_335) );
AND2x4_ASAP7_75t_L g289 ( .A(n_267), .B(n_273), .Y(n_289) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
INVx1_ASAP7_75t_L g308 ( .A(n_269), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
AND2x4_ASAP7_75t_L g278 ( .A(n_270), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g400 ( .A(n_270), .Y(n_400) );
INVx2_ASAP7_75t_L g286 ( .A(n_271), .Y(n_286) );
AND2x2_ASAP7_75t_L g314 ( .A(n_271), .B(n_273), .Y(n_314) );
INVx3_ASAP7_75t_L g322 ( .A(n_271), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_271), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g307 ( .A(n_272), .Y(n_307) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
BUFx2_ASAP7_75t_L g323 ( .A(n_274), .Y(n_323) );
OAI222xp33_ASAP7_75t_L g446 ( .A1(n_276), .A2(n_436), .B1(n_447), .B2(n_450), .C1(n_452), .C2(n_454), .Y(n_446) );
INVx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g387 ( .A(n_278), .Y(n_387) );
AND2x2_ASAP7_75t_L g451 ( .A(n_278), .B(n_321), .Y(n_451) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_281), .B(n_372), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_290), .B1(n_298), .B2(n_300), .C(n_305), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g373 ( .A(n_286), .Y(n_373) );
INVx2_ASAP7_75t_L g435 ( .A(n_287), .Y(n_435) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx2_ASAP7_75t_L g336 ( .A(n_288), .Y(n_336) );
AND2x2_ASAP7_75t_L g372 ( .A(n_288), .B(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g338 ( .A(n_289), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g364 ( .A(n_289), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g453 ( .A(n_289), .Y(n_453) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g402 ( .A(n_293), .Y(n_402) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g425 ( .A(n_295), .B(n_303), .Y(n_425) );
AND2x2_ASAP7_75t_L g448 ( .A(n_295), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g309 ( .A(n_297), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g444 ( .A(n_297), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_298), .A2(n_352), .B1(n_386), .B2(n_388), .Y(n_385) );
OAI21xp5_ASAP7_75t_L g413 ( .A1(n_298), .A2(n_414), .B(n_417), .Y(n_413) );
INVxp67_ASAP7_75t_L g330 ( .A(n_299), .Y(n_330) );
INVx2_ASAP7_75t_SL g434 ( .A(n_299), .Y(n_434) );
AND2x4_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
OR2x2_ASAP7_75t_L g347 ( .A(n_301), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g445 ( .A(n_301), .B(n_444), .Y(n_445) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g318 ( .A(n_303), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_303), .B(n_327), .Y(n_343) );
INVx2_ASAP7_75t_L g370 ( .A(n_303), .Y(n_370) );
OAI22xp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_309), .B1(n_311), .B2(n_313), .Y(n_305) );
NOR2xp33_ASAP7_75t_SL g306 ( .A(n_307), .B(n_308), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_307), .A2(n_381), .B1(n_394), .B2(n_396), .Y(n_393) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g403 ( .A(n_312), .B(n_404), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_320), .B(n_324), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g384 ( .A(n_317), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_317), .B(n_367), .Y(n_395) );
INVx1_ASAP7_75t_L g353 ( .A(n_319), .Y(n_353) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_321), .B(n_334), .Y(n_426) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OAI21xp33_ASAP7_75t_L g439 ( .A1(n_322), .A2(n_440), .B(n_442), .Y(n_439) );
OAI21xp5_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_329), .B(n_337), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx1_ASAP7_75t_L g383 ( .A(n_328), .Y(n_383) );
INVx1_ASAP7_75t_L g449 ( .A(n_328), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g422 ( .A(n_332), .Y(n_422) );
OR2x2_ASAP7_75t_L g433 ( .A(n_333), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND3xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .C(n_342), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_338), .A2(n_399), .B1(n_401), .B2(n_403), .Y(n_398) );
INVx1_ASAP7_75t_L g365 ( .A(n_339), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_340), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g378 ( .A(n_341), .Y(n_378) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_343), .B(n_347), .Y(n_346) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_343), .A2(n_406), .B1(n_409), .B2(n_412), .C(n_413), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_349), .B(n_350), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g354 ( .A(n_348), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_355), .B1(n_356), .B2(n_835), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g437 ( .A(n_359), .B(n_415), .Y(n_437) );
NAND4xp25_ASAP7_75t_L g360 ( .A(n_361), .B(n_391), .C(n_418), .D(n_438), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_374), .Y(n_361) );
OAI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_366), .B1(n_368), .B2(n_369), .C(n_371), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_364), .A2(n_421), .B1(n_443), .B2(n_445), .Y(n_442) );
INVx1_ASAP7_75t_L g417 ( .A(n_366), .Y(n_417) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g401 ( .A(n_367), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_367), .B(n_410), .Y(n_409) );
NAND2x1_ASAP7_75t_L g454 ( .A(n_367), .B(n_455), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_369), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g376 ( .A(n_373), .B(n_377), .Y(n_376) );
OAI21xp33_ASAP7_75t_SL g374 ( .A1(n_375), .A2(n_380), .B(n_385), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NOR2x1_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g404 ( .A(n_390), .Y(n_404) );
AOI211xp5_ASAP7_75t_L g418 ( .A1(n_390), .A2(n_419), .B(n_423), .C(n_429), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_405), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_393), .B(n_398), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g452 ( .A(n_400), .B(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x4_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx3_ASAP7_75t_L g456 ( .A(n_416), .Y(n_456) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND2x1p5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI22xp33_ASAP7_75t_R g429 ( .A1(n_430), .A2(n_433), .B1(n_435), .B2(n_436), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g443 ( .A(n_432), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_439), .B(n_446), .Y(n_438) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_673), .Y(n_458) );
NOR2xp67_ASAP7_75t_L g459 ( .A(n_460), .B(n_615), .Y(n_459) );
NAND3xp33_ASAP7_75t_SL g460 ( .A(n_461), .B(n_552), .C(n_597), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_508), .B(n_529), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_462), .A2(n_553), .B1(n_572), .B2(n_584), .Y(n_552) );
AOI22x1_ASAP7_75t_L g677 ( .A1(n_462), .A2(n_678), .B1(n_682), .B2(n_683), .Y(n_677) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_480), .Y(n_463) );
OR2x2_ASAP7_75t_L g638 ( .A(n_464), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_473), .Y(n_464) );
OR2x2_ASAP7_75t_L g513 ( .A(n_465), .B(n_473), .Y(n_513) );
AND2x2_ASAP7_75t_L g556 ( .A(n_465), .B(n_557), .Y(n_556) );
INVx2_ASAP7_75t_SL g564 ( .A(n_465), .Y(n_564) );
BUFx2_ASAP7_75t_L g614 ( .A(n_465), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_469), .A2(n_505), .B(n_506), .Y(n_504) );
OAI21x1_ASAP7_75t_L g533 ( .A1(n_469), .A2(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g528 ( .A(n_470), .Y(n_528) );
AND2x2_ASAP7_75t_L g559 ( .A(n_473), .B(n_496), .Y(n_559) );
INVx1_ASAP7_75t_L g566 ( .A(n_473), .Y(n_566) );
INVx1_ASAP7_75t_L g571 ( .A(n_473), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_473), .B(n_564), .Y(n_633) );
INVx1_ASAP7_75t_L g654 ( .A(n_473), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_473), .B(n_557), .Y(n_724) );
INVx1_ASAP7_75t_L g617 ( .A(n_480), .Y(n_617) );
OR2x2_ASAP7_75t_L g669 ( .A(n_480), .B(n_633), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_496), .Y(n_480) );
AND2x2_ASAP7_75t_L g514 ( .A(n_481), .B(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g562 ( .A(n_481), .B(n_563), .Y(n_562) );
INVxp67_ASAP7_75t_L g568 ( .A(n_481), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_481), .B(n_511), .Y(n_645) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g557 ( .A(n_482), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_491), .B(n_494), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_487), .B(n_489), .Y(n_484) );
BUFx4f_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_490), .B(n_503), .Y(n_502) );
INVx3_ASAP7_75t_L g511 ( .A(n_496), .Y(n_511) );
INVx1_ASAP7_75t_L g611 ( .A(n_496), .Y(n_611) );
AND2x2_ASAP7_75t_L g613 ( .A(n_496), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g631 ( .A(n_496), .B(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g653 ( .A(n_496), .B(n_654), .Y(n_653) );
NAND2x1p5_ASAP7_75t_SL g664 ( .A(n_496), .B(n_640), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_496), .B(n_571), .Y(n_754) );
AND2x4_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_504), .B(n_507), .Y(n_498) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_514), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_509), .A2(n_693), .B1(n_694), .B2(n_696), .Y(n_692) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_512), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_510), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_510), .B(n_749), .Y(n_748) );
OR2x2_ASAP7_75t_L g771 ( .A(n_510), .B(n_629), .Y(n_771) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x4_ASAP7_75t_L g570 ( .A(n_511), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_511), .B(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g659 ( .A(n_511), .B(n_660), .Y(n_659) );
AND2x4_ASAP7_75t_L g610 ( .A(n_512), .B(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g700 ( .A(n_513), .Y(n_700) );
OR2x2_ASAP7_75t_L g774 ( .A(n_513), .B(n_701), .Y(n_774) );
INVx1_ASAP7_75t_L g605 ( .A(n_514), .Y(n_605) );
INVx3_ASAP7_75t_L g609 ( .A(n_515), .Y(n_609) );
BUFx2_ASAP7_75t_L g620 ( .A(n_515), .Y(n_620) );
BUFx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g590 ( .A(n_516), .B(n_541), .Y(n_590) );
INVx2_ASAP7_75t_L g636 ( .A(n_516), .Y(n_636) );
INVx1_ASAP7_75t_L g668 ( .A(n_516), .Y(n_668) );
AND2x2_ASAP7_75t_L g681 ( .A(n_516), .B(n_578), .Y(n_681) );
AND2x2_ASAP7_75t_L g703 ( .A(n_516), .B(n_602), .Y(n_703) );
NAND2x1p5_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
OAI21x1_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_524), .B(n_527), .Y(n_518) );
INVx2_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g694 ( .A(n_530), .B(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_530), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g719 ( .A(n_530), .B(n_587), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_530), .B(n_721), .Y(n_720) );
AND2x4_ASAP7_75t_L g530 ( .A(n_531), .B(n_541), .Y(n_530) );
INVx2_ASAP7_75t_L g576 ( .A(n_531), .Y(n_576) );
AND2x2_ASAP7_75t_L g603 ( .A(n_531), .B(n_604), .Y(n_603) );
AOI21x1_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_536), .B(n_539), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g577 ( .A(n_541), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g596 ( .A(n_541), .Y(n_596) );
INVx2_ASAP7_75t_L g604 ( .A(n_541), .Y(n_604) );
OR2x2_ASAP7_75t_L g624 ( .A(n_541), .B(n_578), .Y(n_624) );
AND2x2_ASAP7_75t_L g635 ( .A(n_541), .B(n_636), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_558), .B1(n_560), .B2(n_565), .C(n_567), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OAI32xp33_ASAP7_75t_L g665 ( .A1(n_555), .A2(n_569), .A3(n_666), .B1(n_669), .B2(n_670), .Y(n_665) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g655 ( .A(n_556), .Y(n_655) );
AND2x2_ASAP7_75t_L g691 ( .A(n_556), .B(n_570), .Y(n_691) );
INVx1_ASAP7_75t_L g755 ( .A(n_556), .Y(n_755) );
OR2x2_ASAP7_75t_L g629 ( .A(n_557), .B(n_564), .Y(n_629) );
INVx2_ASAP7_75t_L g640 ( .A(n_557), .Y(n_640) );
BUFx2_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g779 ( .A(n_559), .B(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVxp67_ASAP7_75t_L g766 ( .A(n_562), .Y(n_766) );
INVx1_ASAP7_75t_L g780 ( .A(n_562), .Y(n_780) );
OR2x2_ASAP7_75t_L g660 ( .A(n_563), .B(n_640), .Y(n_660) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_565), .B(n_660), .Y(n_682) );
INVx1_ASAP7_75t_L g713 ( .A(n_565), .Y(n_713) );
BUFx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g747 ( .A(n_566), .Y(n_747) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2x1_ASAP7_75t_L g716 ( .A(n_568), .B(n_717), .Y(n_716) );
OAI21xp5_ASAP7_75t_SL g738 ( .A1(n_569), .A2(n_739), .B(n_744), .Y(n_738) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_577), .Y(n_573) );
AND2x2_ASAP7_75t_L g648 ( .A(n_574), .B(n_590), .Y(n_648) );
INVxp67_ASAP7_75t_SL g778 ( .A(n_574), .Y(n_778) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g680 ( .A(n_575), .Y(n_680) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g662 ( .A(n_576), .B(n_636), .Y(n_662) );
AND2x2_ASAP7_75t_L g733 ( .A(n_576), .B(n_604), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_577), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g661 ( .A(n_577), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g740 ( .A(n_577), .B(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g589 ( .A(n_578), .Y(n_589) );
INVx2_ASAP7_75t_L g602 ( .A(n_578), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_578), .B(n_593), .Y(n_650) );
AND2x2_ASAP7_75t_L g710 ( .A(n_578), .B(n_604), .Y(n_710) );
NAND2xp33_ASAP7_75t_SL g584 ( .A(n_585), .B(n_591), .Y(n_584) );
INVx2_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g685 ( .A(n_588), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_588), .B(n_668), .Y(n_760) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g592 ( .A(n_589), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g721 ( .A(n_589), .B(n_636), .Y(n_721) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
OR2x2_ASAP7_75t_L g666 ( .A(n_592), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g623 ( .A(n_593), .Y(n_623) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g649 ( .A(n_596), .B(n_650), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_610), .B1(n_612), .B2(n_613), .Y(n_597) );
OAI21xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_605), .B(n_606), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g612 ( .A(n_600), .B(n_609), .Y(n_612) );
BUFx2_ASAP7_75t_L g630 ( .A(n_600), .Y(n_630) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVx1_ASAP7_75t_L g641 ( .A(n_601), .Y(n_641) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g656 ( .A(n_603), .B(n_620), .Y(n_656) );
INVx2_ASAP7_75t_L g672 ( .A(n_603), .Y(n_672) );
AND2x2_ASAP7_75t_L g714 ( .A(n_603), .B(n_636), .Y(n_714) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g689 ( .A(n_609), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g736 ( .A(n_610), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g767 ( .A(n_611), .Y(n_767) );
INVx2_ASAP7_75t_L g706 ( .A(n_614), .Y(n_706) );
NAND4xp25_ASAP7_75t_L g615 ( .A(n_616), .B(n_625), .C(n_642), .D(n_657), .Y(n_615) );
NAND2xp33_ASAP7_75t_SL g616 ( .A(n_617), .B(n_618), .Y(n_616) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_618), .A2(n_696), .B1(n_712), .B2(n_714), .C(n_715), .Y(n_711) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2x1_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g693 ( .A(n_622), .Y(n_693) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx2_ASAP7_75t_L g686 ( .A(n_623), .Y(n_686) );
INVx2_ASAP7_75t_L g758 ( .A(n_624), .Y(n_758) );
AOI222xp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_630), .B1(n_631), .B2(n_634), .C1(n_637), .C2(n_641), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g712 ( .A(n_628), .B(n_713), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_628), .A2(n_740), .B(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g751 ( .A(n_629), .B(n_695), .Y(n_751) );
OAI21xp33_ASAP7_75t_SL g725 ( .A1(n_630), .A2(n_651), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g644 ( .A(n_633), .B(n_645), .Y(n_644) );
INVxp67_ASAP7_75t_SL g696 ( .A(n_633), .Y(n_696) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
BUFx2_ASAP7_75t_L g695 ( .A(n_636), .Y(n_695) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g701 ( .A(n_640), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g642 ( .A1(n_643), .A2(n_646), .B1(n_651), .B2(n_656), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_648), .A2(n_658), .B1(n_661), .B2(n_663), .C(n_665), .Y(n_657) );
INVx3_ASAP7_75t_R g772 ( .A(n_649), .Y(n_772) );
INVx1_ASAP7_75t_L g690 ( .A(n_650), .Y(n_690) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVxp67_ASAP7_75t_SL g707 ( .A(n_653), .Y(n_707) );
INVx1_ASAP7_75t_L g717 ( .A(n_653), .Y(n_717) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_662), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g735 ( .A(n_662), .Y(n_735) );
AND2x2_ASAP7_75t_L g763 ( .A(n_662), .B(n_710), .Y(n_763) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g757 ( .A(n_667), .B(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx3_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NOR2x1_ASAP7_75t_L g673 ( .A(n_674), .B(n_729), .Y(n_673) );
NAND3xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_711), .C(n_725), .Y(n_674) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_687), .C(n_697), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI21xp33_ASAP7_75t_L g688 ( .A1(n_678), .A2(n_689), .B(n_691), .Y(n_688) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx1_ASAP7_75t_L g728 ( .A(n_680), .Y(n_728) );
AND2x2_ASAP7_75t_L g769 ( .A(n_680), .B(n_758), .Y(n_769) );
NAND2x1_ASAP7_75t_L g727 ( .A(n_681), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g749 ( .A(n_686), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_692), .Y(n_687) );
INVx1_ASAP7_75t_L g741 ( .A(n_695), .Y(n_741) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_702), .B1(n_704), .B2(n_708), .Y(n_697) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g737 ( .A(n_701), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_703), .B(n_733), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g776 ( .A(n_709), .Y(n_776) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
OAI22xp33_ASAP7_75t_SL g715 ( .A1(n_716), .A2(n_718), .B1(n_720), .B2(n_722), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_756), .Y(n_729) );
O2A1O1Ixp33_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_734), .B(n_736), .C(n_738), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI21xp33_ASAP7_75t_L g745 ( .A1(n_732), .A2(n_746), .B(n_748), .Y(n_745) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
O2A1O1Ixp5_ASAP7_75t_SL g756 ( .A1(n_736), .A2(n_757), .B(n_759), .C(n_761), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_740), .A2(n_745), .B1(n_750), .B2(n_752), .Y(n_744) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
OR2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OAI211xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_764), .B(n_768), .C(n_775), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_770), .B1(n_772), .B2(n_773), .Y(n_768) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OAI21xp5_ASAP7_75t_SL g775 ( .A1(n_776), .A2(n_777), .B(n_779), .Y(n_775) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
BUFx4f_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx3_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
OR2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_789), .Y(n_784) );
BUFx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NOR2x1_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g809 ( .A(n_788), .Y(n_809) );
OR2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
AND2x2_ASAP7_75t_L g824 ( .A(n_790), .B(n_825), .Y(n_824) );
NOR2xp33_ASAP7_75t_L g825 ( .A(n_791), .B(n_826), .Y(n_825) );
NAND2xp5_ASAP7_75t_SL g791 ( .A(n_792), .B(n_795), .Y(n_791) );
BUFx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_793), .B(n_820), .Y(n_819) );
INVx3_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_794), .B(n_804), .Y(n_832) );
INVx2_ASAP7_75t_SL g821 ( .A(n_795), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_803), .Y(n_798) );
INVx1_ASAP7_75t_L g813 ( .A(n_799), .Y(n_813) );
BUFx2_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
INVx3_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx5_ASAP7_75t_L g812 ( .A(n_805), .Y(n_812) );
INVx5_ASAP7_75t_L g817 ( .A(n_805), .Y(n_817) );
CKINVDCx8_ASAP7_75t_R g827 ( .A(n_805), .Y(n_827) );
AND2x6_ASAP7_75t_SL g805 ( .A(n_806), .B(n_809), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
BUFx2_ASAP7_75t_SL g811 ( .A(n_812), .Y(n_811) );
NOR2xp67_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
BUFx3_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
BUFx3_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
OR2x4_ASAP7_75t_L g831 ( .A(n_820), .B(n_832), .Y(n_831) );
BUFx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_828), .B1(n_829), .B2(n_833), .Y(n_822) );
INVx3_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx3_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx6_ASAP7_75t_SL g829 ( .A(n_830), .Y(n_829) );
BUFx10_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
endmodule