module fake_netlist_5_1792_n_1733 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1733);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1733;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_696;
wire n_550;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1587;
wire n_1473;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_12),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_27),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_7),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_66),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_15),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_68),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_57),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_77),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_78),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_47),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_89),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_47),
.Y(n_173)
);

INVxp67_ASAP7_75t_SL g174 ( 
.A(n_46),
.Y(n_174)
);

INVx4_ASAP7_75t_R g175 ( 
.A(n_71),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_107),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_123),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_90),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_105),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_65),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_50),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_111),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_52),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_97),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_31),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_55),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_35),
.Y(n_189)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_33),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_85),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_72),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_21),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_54),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_126),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_45),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_79),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_29),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_17),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_23),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_51),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_114),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_9),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_129),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_2),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_110),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_59),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_147),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_8),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_141),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_82),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_38),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_83),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_38),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_3),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_14),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_70),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_21),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_104),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_153),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_143),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_17),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_49),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_96),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_24),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_60),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_0),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_127),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_122),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_80),
.Y(n_233)
);

BUFx8_ASAP7_75t_SL g234 ( 
.A(n_148),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_119),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_41),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_32),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_50),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_28),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_62),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_128),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_92),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_86),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_135),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_109),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_61),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_48),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_26),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_88),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_56),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_132),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_117),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_155),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_102),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_74),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_8),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_58),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_37),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_30),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_48),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_115),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_91),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_34),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_151),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_63),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_154),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_136),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_131),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_41),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_39),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_28),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_4),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_64),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_43),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_15),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_46),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_12),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_125),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_84),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_75),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_149),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_20),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_2),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_42),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_69),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_121),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_106),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_26),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_6),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_24),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_142),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_100),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_45),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_36),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_53),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_43),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_6),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_16),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_22),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_23),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_25),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_120),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_25),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_37),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_31),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_95),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_19),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_140),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_9),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_10),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_219),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_200),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_252),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_179),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_190),
.B(n_0),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_200),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_200),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_228),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_234),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_200),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_200),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_205),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_186),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_193),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_205),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_193),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_205),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_205),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_205),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_203),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_173),
.B(n_1),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_204),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_196),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_241),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_206),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_163),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_212),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_282),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_215),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_221),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_222),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_260),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_223),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_182),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_235),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_240),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_289),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_242),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_260),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_239),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_243),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_263),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_169),
.B(n_1),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_263),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_183),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_246),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_239),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_250),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_310),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_251),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_182),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_257),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_169),
.B(n_3),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_187),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_156),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_261),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_201),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_262),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_266),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_267),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_217),
.B(n_4),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_239),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_216),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_241),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_273),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_213),
.B(n_5),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_218),
.Y(n_378)
);

BUFx6f_ASAP7_75t_SL g379 ( 
.A(n_281),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_281),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_305),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_305),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_312),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_366),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_345),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_312),
.B(n_213),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_366),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_345),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_316),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_362),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_317),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_317),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_320),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_311),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_320),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_321),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_321),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_322),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_322),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_325),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_325),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_327),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_327),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_315),
.B(n_185),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_328),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_328),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_329),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_329),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_338),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_338),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_341),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_377),
.B(n_233),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_356),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_356),
.Y(n_417)
);

AND2x6_ASAP7_75t_L g418 ( 
.A(n_354),
.B(n_233),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_334),
.B(n_249),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_377),
.B(n_249),
.Y(n_420)
);

OA21x2_ASAP7_75t_L g421 ( 
.A1(n_360),
.A2(n_247),
.B(n_220),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_360),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_365),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_334),
.B(n_195),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_336),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_334),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_368),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_368),
.Y(n_429)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_375),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_324),
.B(n_162),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_326),
.B(n_380),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_364),
.B(n_157),
.Y(n_433)
);

BUFx12f_ASAP7_75t_L g434 ( 
.A(n_319),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_374),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_374),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_378),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_375),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_378),
.Y(n_439)
);

NAND3xp33_ASAP7_75t_L g440 ( 
.A(n_331),
.B(n_296),
.C(n_283),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_375),
.Y(n_441)
);

BUFx8_ASAP7_75t_L g442 ( 
.A(n_379),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_343),
.Y(n_443)
);

OAI21x1_ASAP7_75t_L g444 ( 
.A1(n_331),
.A2(n_161),
.B(n_160),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_343),
.B(n_162),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_350),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_350),
.Y(n_447)
);

NAND2xp33_ASAP7_75t_L g448 ( 
.A(n_418),
.B(n_323),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_401),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_406),
.B(n_330),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_385),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_385),
.Y(n_452)
);

AOI21x1_ASAP7_75t_L g453 ( 
.A1(n_433),
.A2(n_420),
.B(n_415),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_441),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_430),
.B(n_332),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_427),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_419),
.B(n_441),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_401),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_401),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_391),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_430),
.B(n_337),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_406),
.B(n_339),
.Y(n_463)
);

INVx5_ASAP7_75t_L g464 ( 
.A(n_391),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_385),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_391),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_427),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_401),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_403),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_388),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_418),
.A2(n_314),
.B1(n_269),
.B2(n_259),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_391),
.Y(n_472)
);

BUFx8_ASAP7_75t_SL g473 ( 
.A(n_434),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_388),
.Y(n_474)
);

OAI22xp33_ASAP7_75t_L g475 ( 
.A1(n_433),
.A2(n_387),
.B1(n_432),
.B2(n_318),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_388),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_403),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_387),
.B(n_373),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_419),
.B(n_353),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_388),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_432),
.B(n_340),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_431),
.B(n_344),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_403),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_431),
.B(n_346),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_430),
.B(n_347),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_433),
.A2(n_352),
.B1(n_349),
.B2(n_335),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_430),
.B(n_357),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_418),
.A2(n_348),
.B1(n_372),
.B2(n_300),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_391),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_403),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_394),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_391),
.Y(n_493)
);

OAI22x1_ASAP7_75t_L g494 ( 
.A1(n_387),
.A2(n_384),
.B1(n_425),
.B2(n_358),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_438),
.Y(n_495)
);

OR2x6_ASAP7_75t_L g496 ( 
.A(n_434),
.B(n_372),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_442),
.B(n_359),
.Y(n_497)
);

OAI22xp33_ASAP7_75t_L g498 ( 
.A1(n_440),
.A2(n_293),
.B1(n_373),
.B2(n_211),
.Y(n_498)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_424),
.B(n_195),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_L g500 ( 
.A(n_418),
.B(n_363),
.Y(n_500)
);

BUFx10_ASAP7_75t_L g501 ( 
.A(n_418),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_394),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_438),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_430),
.B(n_367),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_419),
.B(n_353),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_424),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_430),
.B(n_369),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_441),
.B(n_370),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_443),
.Y(n_509)
);

OAI22xp33_ASAP7_75t_L g510 ( 
.A1(n_440),
.A2(n_415),
.B1(n_420),
.B2(n_445),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_418),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_394),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_443),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_391),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_424),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_445),
.B(n_371),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_397),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_442),
.B(n_376),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_443),
.Y(n_519)
);

BUFx10_ASAP7_75t_L g520 ( 
.A(n_418),
.Y(n_520)
);

BUFx6f_ASAP7_75t_SL g521 ( 
.A(n_418),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_391),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_384),
.B(n_342),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_442),
.B(n_361),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_397),
.Y(n_525)
);

AND2x6_ASAP7_75t_L g526 ( 
.A(n_424),
.B(n_195),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_442),
.B(n_333),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_418),
.B(n_208),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_397),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_440),
.B(n_379),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_397),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_418),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_419),
.B(n_355),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_447),
.B(n_355),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_396),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_399),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_399),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_421),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_421),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_399),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_396),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_391),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_421),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_418),
.B(n_255),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_399),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_408),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_424),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_418),
.B(n_292),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_408),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_408),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_421),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_421),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_421),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_423),
.B(n_379),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_408),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_421),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_390),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_393),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_396),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_383),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_442),
.B(n_351),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_393),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_444),
.A2(n_307),
.B1(n_297),
.B2(n_301),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_390),
.Y(n_564)
);

INVx8_ASAP7_75t_L g565 ( 
.A(n_434),
.Y(n_565)
);

INVxp67_ASAP7_75t_SL g566 ( 
.A(n_390),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_383),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_424),
.B(n_306),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_393),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_423),
.B(n_381),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_383),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_393),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_442),
.B(n_382),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_389),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_389),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_415),
.B(n_165),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_389),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_395),
.B(n_400),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_395),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_423),
.B(n_313),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_395),
.B(n_278),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_447),
.B(n_174),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_390),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_400),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_390),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_434),
.B(n_164),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_400),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_402),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_390),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_444),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_392),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_402),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_402),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_423),
.B(n_425),
.Y(n_594)
);

BUFx4f_ASAP7_75t_L g595 ( 
.A(n_446),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_SL g596 ( 
.A(n_565),
.B(n_197),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_481),
.B(n_444),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_516),
.B(n_444),
.Y(n_598)
);

OAI221xp5_ASAP7_75t_L g599 ( 
.A1(n_471),
.A2(n_420),
.B1(n_417),
.B2(n_437),
.C(n_436),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_463),
.B(n_423),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_580),
.A2(n_280),
.B1(n_279),
.B2(n_177),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_570),
.B(n_423),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_547),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_528),
.B(n_182),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_458),
.B(n_446),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_458),
.B(n_446),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_451),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_547),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_479),
.B(n_447),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_471),
.A2(n_232),
.B1(n_167),
.B2(n_168),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_451),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_538),
.A2(n_417),
.B1(n_437),
.B2(n_436),
.Y(n_612)
);

OAI22xp33_ASAP7_75t_SL g613 ( 
.A1(n_450),
.A2(n_170),
.B1(n_159),
.B2(n_158),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_452),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_560),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_510),
.B(n_446),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_538),
.A2(n_417),
.B1(n_437),
.B2(n_436),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_594),
.B(n_446),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_478),
.Y(n_619)
);

BUFx8_ASAP7_75t_L g620 ( 
.A(n_478),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_467),
.B(n_422),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_475),
.B(n_165),
.Y(n_622)
);

OR2x6_ASAP7_75t_L g623 ( 
.A(n_565),
.B(n_166),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_523),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_467),
.B(n_422),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_454),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_520),
.B(n_446),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_520),
.B(n_446),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_560),
.Y(n_629)
);

INVx8_ASAP7_75t_L g630 ( 
.A(n_565),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_453),
.B(n_446),
.Y(n_631)
);

NAND2x1_ASAP7_75t_L g632 ( 
.A(n_539),
.B(n_175),
.Y(n_632)
);

A2O1A1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_539),
.A2(n_447),
.B(n_426),
.C(n_435),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_453),
.B(n_446),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_567),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_582),
.B(n_386),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_452),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_534),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_455),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_520),
.B(n_195),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_520),
.B(n_195),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_532),
.B(n_291),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_582),
.B(n_386),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_566),
.B(n_386),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_495),
.B(n_156),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_509),
.B(n_386),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_509),
.B(n_386),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_543),
.A2(n_552),
.B1(n_553),
.B2(n_551),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_534),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_473),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_449),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_543),
.A2(n_422),
.B1(n_435),
.B2(n_429),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_565),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_567),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_495),
.B(n_167),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_449),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_503),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_455),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_503),
.B(n_426),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_506),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_513),
.B(n_386),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_513),
.B(n_413),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_532),
.B(n_291),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_459),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_457),
.B(n_426),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_459),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_460),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_519),
.B(n_413),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_519),
.B(n_413),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_465),
.Y(n_670)
);

INVxp67_ASAP7_75t_SL g671 ( 
.A(n_557),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_535),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_479),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_504),
.B(n_413),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_505),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_465),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_505),
.B(n_413),
.Y(n_677)
);

OAI221xp5_ASAP7_75t_L g678 ( 
.A1(n_489),
.A2(n_428),
.B1(n_435),
.B2(n_429),
.C(n_209),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_460),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_532),
.B(n_291),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_533),
.B(n_413),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_533),
.B(n_407),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_506),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_508),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_532),
.B(n_291),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_470),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_551),
.A2(n_429),
.B(n_428),
.C(n_412),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_468),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_469),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_469),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_501),
.B(n_291),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_482),
.A2(n_171),
.B1(n_172),
.B2(n_168),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_535),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_541),
.B(n_428),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_515),
.B(n_407),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_484),
.B(n_171),
.Y(n_696)
);

NOR3xp33_ASAP7_75t_L g697 ( 
.A(n_487),
.B(n_202),
.C(n_207),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_501),
.B(n_511),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_515),
.B(n_407),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_576),
.B(n_172),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_498),
.B(n_176),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_590),
.A2(n_409),
.B(n_439),
.Y(n_702)
);

NOR2x1p5_ASAP7_75t_L g703 ( 
.A(n_541),
.B(n_559),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_563),
.A2(n_199),
.B1(n_178),
.B2(n_184),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_544),
.A2(n_244),
.B1(n_188),
.B2(n_192),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_477),
.B(n_409),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_477),
.B(n_409),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_501),
.B(n_182),
.Y(n_708)
);

AO22x2_ASAP7_75t_L g709 ( 
.A1(n_561),
.A2(n_264),
.B1(n_210),
.B2(n_226),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_559),
.B(n_158),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_568),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_552),
.A2(n_284),
.B1(n_237),
.B2(n_182),
.Y(n_712)
);

OAI22xp33_ASAP7_75t_L g713 ( 
.A1(n_553),
.A2(n_556),
.B1(n_496),
.B2(n_586),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_556),
.A2(n_412),
.B(n_439),
.C(n_416),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_SL g715 ( 
.A(n_573),
.B(n_159),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_511),
.B(n_182),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_483),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_530),
.B(n_176),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_483),
.B(n_398),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_491),
.B(n_398),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_491),
.B(n_558),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_574),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_511),
.B(n_182),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_493),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_574),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_558),
.B(n_398),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_SL g727 ( 
.A(n_565),
.B(n_177),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_494),
.B(n_496),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_448),
.A2(n_285),
.B1(n_181),
.B2(n_231),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_496),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_494),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_470),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_548),
.B(n_590),
.Y(n_733)
);

O2A1O1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_500),
.A2(n_439),
.B(n_416),
.C(n_412),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_586),
.Y(n_735)
);

INVxp67_ASAP7_75t_SL g736 ( 
.A(n_557),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_557),
.B(n_182),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_581),
.B(n_180),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_562),
.B(n_398),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_474),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_562),
.B(n_398),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_586),
.B(n_416),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_569),
.B(n_398),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_474),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_569),
.B(n_404),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_456),
.B(n_180),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_564),
.B(n_254),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_462),
.B(n_181),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_586),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_575),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_572),
.B(n_404),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_577),
.B(n_404),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_577),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_579),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_476),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_579),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_584),
.B(n_404),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_571),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_584),
.B(n_404),
.Y(n_759)
);

OR2x6_ASAP7_75t_L g760 ( 
.A(n_586),
.B(n_496),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_587),
.B(n_404),
.Y(n_761)
);

INVx8_ASAP7_75t_L g762 ( 
.A(n_496),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_521),
.A2(n_254),
.B1(n_227),
.B2(n_229),
.Y(n_763)
);

OAI21xp33_ASAP7_75t_L g764 ( 
.A1(n_622),
.A2(n_288),
.B(n_170),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_711),
.B(n_485),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_684),
.B(n_488),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_600),
.B(n_507),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_621),
.B(n_625),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_657),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_657),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_673),
.B(n_524),
.Y(n_771)
);

O2A1O1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_599),
.A2(n_593),
.B(n_592),
.C(n_588),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_L g773 ( 
.A1(n_597),
.A2(n_598),
.B(n_616),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_762),
.B(n_527),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_683),
.B(n_564),
.Y(n_775)
);

AOI21xp33_ASAP7_75t_L g776 ( 
.A1(n_622),
.A2(n_701),
.B(n_718),
.Y(n_776)
);

AOI22x1_ASAP7_75t_L g777 ( 
.A1(n_671),
.A2(n_593),
.B1(n_592),
.B2(n_588),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_698),
.A2(n_595),
.B(n_490),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_712),
.A2(n_521),
.B1(n_499),
.B2(n_526),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_619),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_615),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_672),
.Y(n_782)
);

O2A1O1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_687),
.A2(n_578),
.B(n_497),
.C(n_518),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_698),
.A2(n_595),
.B(n_490),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_615),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_636),
.A2(n_595),
.B(n_490),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_648),
.A2(n_712),
.B1(n_660),
.B2(n_718),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_624),
.B(n_564),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_694),
.B(n_305),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_683),
.B(n_583),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_643),
.A2(n_514),
.B(n_493),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_683),
.B(n_583),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_659),
.B(n_554),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_687),
.A2(n_571),
.B(n_268),
.C(n_295),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_683),
.B(n_583),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_631),
.A2(n_493),
.B(n_514),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_648),
.A2(n_521),
.B1(n_589),
.B2(n_585),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_713),
.B(n_585),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_701),
.B(n_585),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_713),
.B(n_589),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_634),
.A2(n_514),
.B(n_493),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_627),
.A2(n_514),
.B(n_493),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_627),
.A2(n_514),
.B(n_461),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_629),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_665),
.B(n_461),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_675),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_738),
.B(n_461),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_628),
.A2(n_522),
.B(n_466),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_693),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_629),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_738),
.B(n_466),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_609),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_628),
.A2(n_522),
.B(n_466),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_609),
.B(n_472),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_733),
.A2(n_472),
.B(n_542),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_696),
.A2(n_253),
.B(n_265),
.C(n_245),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_645),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_655),
.B(n_416),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_696),
.A2(n_700),
.B(n_748),
.C(n_746),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_653),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_677),
.B(n_542),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_635),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_746),
.B(n_542),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_638),
.A2(n_198),
.B1(n_308),
.B2(n_232),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_733),
.A2(n_464),
.B(n_591),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_681),
.B(n_591),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_635),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_748),
.B(n_476),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_603),
.A2(n_499),
.B1(n_526),
.B2(n_591),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_655),
.B(n_710),
.Y(n_830)
);

O2A1O1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_633),
.A2(n_555),
.B(n_550),
.C(n_549),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_714),
.A2(n_480),
.B(n_550),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_605),
.A2(n_464),
.B(n_480),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_742),
.B(n_486),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_606),
.A2(n_464),
.B(n_549),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_703),
.B(n_439),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_654),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_654),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_731),
.B(n_189),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_618),
.A2(n_464),
.B(n_546),
.Y(n_840)
);

NOR3xp33_ASAP7_75t_L g841 ( 
.A(n_613),
.B(n_231),
.C(n_285),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_722),
.Y(n_842)
);

NOR2xp67_ASAP7_75t_L g843 ( 
.A(n_601),
.B(n_286),
.Y(n_843)
);

OR2x2_ASAP7_75t_L g844 ( 
.A(n_610),
.B(n_288),
.Y(n_844)
);

AO21x1_ASAP7_75t_L g845 ( 
.A1(n_704),
.A2(n_555),
.B(n_546),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_742),
.B(n_486),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_758),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_644),
.A2(n_464),
.B(n_540),
.Y(n_848)
);

NAND2x1_ASAP7_75t_L g849 ( 
.A(n_724),
.B(n_499),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_674),
.A2(n_464),
.B(n_540),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_649),
.B(n_725),
.Y(n_851)
);

AO21x1_ASAP7_75t_L g852 ( 
.A1(n_715),
.A2(n_545),
.B(n_537),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_714),
.A2(n_545),
.B(n_537),
.Y(n_853)
);

AO21x1_ASAP7_75t_L g854 ( 
.A1(n_700),
.A2(n_536),
.B(n_531),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_736),
.A2(n_536),
.B(n_531),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_620),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_750),
.B(n_492),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_753),
.B(n_492),
.Y(n_858)
);

O2A1O1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_633),
.A2(n_529),
.B(n_502),
.C(n_525),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_754),
.A2(n_286),
.B1(n_287),
.B2(n_302),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_608),
.A2(n_526),
.B1(n_499),
.B2(n_302),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_602),
.A2(n_529),
.B(n_502),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_756),
.B(n_512),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_724),
.A2(n_525),
.B(n_517),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_620),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_709),
.A2(n_499),
.B1(n_526),
.B2(n_254),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_697),
.B(n_290),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_651),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_724),
.A2(n_405),
.B(n_414),
.Y(n_869)
);

NAND2x1p5_ASAP7_75t_L g870 ( 
.A(n_653),
.B(n_405),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_705),
.A2(n_405),
.B(n_414),
.C(n_411),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_656),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_724),
.A2(n_405),
.B(n_414),
.Y(n_873)
);

NAND2x1p5_ASAP7_75t_L g874 ( 
.A(n_626),
.B(n_405),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_678),
.A2(n_682),
.B(n_679),
.C(n_664),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_758),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_666),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_596),
.B(n_735),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_728),
.B(n_290),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_667),
.B(n_526),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_612),
.A2(n_309),
.B(n_304),
.C(n_303),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_692),
.B(n_294),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_708),
.A2(n_499),
.B1(n_526),
.B2(n_287),
.Y(n_883)
);

OAI21xp33_ASAP7_75t_L g884 ( 
.A1(n_612),
.A2(n_309),
.B(n_304),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_688),
.B(n_499),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_708),
.A2(n_414),
.B(n_411),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_734),
.A2(n_411),
.B(n_271),
.C(n_270),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_716),
.A2(n_411),
.B(n_410),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_689),
.B(n_191),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_690),
.B(n_194),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_716),
.A2(n_410),
.B(n_392),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_717),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_723),
.A2(n_410),
.B(n_392),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_617),
.A2(n_303),
.B(n_299),
.C(n_298),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_749),
.B(n_730),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_607),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_646),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_617),
.B(n_526),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_721),
.B(n_214),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_723),
.A2(n_410),
.B(n_392),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_647),
.A2(n_410),
.B(n_392),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_650),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_611),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_652),
.B(n_410),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_661),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_709),
.A2(n_254),
.B1(n_294),
.B2(n_299),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_652),
.B(n_410),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_702),
.A2(n_258),
.B(n_225),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_760),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_662),
.B(n_254),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_695),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_709),
.B(n_298),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_729),
.B(n_224),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_762),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_L g915 ( 
.A(n_630),
.B(n_254),
.Y(n_915)
);

INVx4_ASAP7_75t_L g916 ( 
.A(n_630),
.Y(n_916)
);

INVx5_ASAP7_75t_L g917 ( 
.A(n_630),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_614),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_699),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_763),
.A2(n_272),
.B(n_236),
.C(n_277),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_760),
.A2(n_256),
.B1(n_238),
.B2(n_276),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_668),
.B(n_410),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_706),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_691),
.A2(n_410),
.B(n_392),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_760),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_707),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_669),
.B(n_392),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_691),
.A2(n_392),
.B(n_275),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_637),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_762),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_640),
.A2(n_392),
.B(n_274),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_639),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_640),
.A2(n_248),
.B(n_230),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_752),
.B(n_254),
.Y(n_934)
);

AO21x1_ASAP7_75t_L g935 ( 
.A1(n_604),
.A2(n_254),
.B(n_7),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_623),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_641),
.A2(n_663),
.B(n_642),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_623),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_737),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_641),
.A2(n_146),
.B(n_137),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_642),
.A2(n_134),
.B(n_130),
.Y(n_941)
);

INVx4_ASAP7_75t_L g942 ( 
.A(n_623),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_658),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_727),
.B(n_5),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_670),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_663),
.A2(n_118),
.B(n_116),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_676),
.Y(n_947)
);

AO22x1_ASAP7_75t_L g948 ( 
.A1(n_719),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_948)
);

NOR3xp33_ASAP7_75t_L g949 ( 
.A(n_776),
.B(n_737),
.C(n_747),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_768),
.B(n_911),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_773),
.A2(n_680),
.B(n_685),
.Y(n_951)
);

BUFx4f_ASAP7_75t_L g952 ( 
.A(n_930),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_930),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_819),
.A2(n_763),
.B1(n_680),
.B2(n_685),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_SL g955 ( 
.A1(n_782),
.A2(n_632),
.B1(n_720),
.B2(n_757),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_823),
.A2(n_761),
.B(n_759),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_842),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_868),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_809),
.Y(n_959)
);

INVxp67_ASAP7_75t_L g960 ( 
.A(n_769),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_872),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_816),
.A2(n_747),
.B(n_751),
.C(n_741),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_767),
.A2(n_811),
.B(n_807),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_789),
.B(n_740),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_816),
.A2(n_739),
.B(n_745),
.C(n_726),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_769),
.Y(n_966)
);

INVxp67_ASAP7_75t_SL g967 ( 
.A(n_812),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_793),
.A2(n_743),
.B(n_744),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_787),
.A2(n_755),
.B1(n_732),
.B2(n_686),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_830),
.B(n_11),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_791),
.A2(n_93),
.B(n_108),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_930),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_766),
.B(n_13),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_881),
.A2(n_14),
.B(n_16),
.C(n_18),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_809),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_770),
.B(n_18),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_919),
.B(n_19),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_902),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_770),
.Y(n_979)
);

NAND2x1p5_ASAP7_75t_L g980 ( 
.A(n_916),
.B(n_112),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_786),
.A2(n_81),
.B(n_98),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_812),
.B(n_99),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_799),
.A2(n_94),
.B1(n_87),
.B2(n_76),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_771),
.B(n_73),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_820),
.Y(n_985)
);

BUFx12f_ASAP7_75t_L g986 ( 
.A(n_856),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_796),
.A2(n_67),
.B(n_22),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_801),
.A2(n_20),
.B(n_27),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_913),
.A2(n_783),
.B(n_799),
.C(n_899),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_930),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_876),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_877),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_771),
.B(n_29),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_R g994 ( 
.A(n_820),
.B(n_49),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_923),
.B(n_926),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_876),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_780),
.B(n_30),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_780),
.Y(n_998)
);

BUFx12f_ASAP7_75t_L g999 ( 
.A(n_865),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_828),
.A2(n_32),
.B(n_33),
.Y(n_1000)
);

AOI21x1_ASAP7_75t_L g1001 ( 
.A1(n_821),
.A2(n_34),
.B(n_35),
.Y(n_1001)
);

AND3x1_ASAP7_75t_L g1002 ( 
.A(n_841),
.B(n_36),
.C(n_39),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_897),
.A2(n_40),
.B(n_42),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_817),
.B(n_879),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_899),
.B(n_40),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_836),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_779),
.A2(n_44),
.B1(n_905),
.B2(n_939),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_781),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_765),
.B(n_44),
.Y(n_1009)
);

INVx5_ASAP7_75t_L g1010 ( 
.A(n_917),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_937),
.A2(n_875),
.B(n_784),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_878),
.B(n_851),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_788),
.B(n_818),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_895),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_779),
.A2(n_939),
.B1(n_805),
.B2(n_898),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_SL g1016 ( 
.A1(n_906),
.A2(n_913),
.B1(n_844),
.B2(n_774),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_785),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_798),
.A2(n_800),
.B1(n_788),
.B2(n_797),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_778),
.A2(n_798),
.B(n_800),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_806),
.B(n_892),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_914),
.B(n_909),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_820),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_925),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_820),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_909),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_804),
.Y(n_1026)
);

O2A1O1Ixp5_ASAP7_75t_L g1027 ( 
.A1(n_854),
.A2(n_852),
.B(n_845),
.C(n_887),
.Y(n_1027)
);

INVx3_ASAP7_75t_SL g1028 ( 
.A(n_774),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_944),
.Y(n_1029)
);

AO21x1_ASAP7_75t_L g1030 ( 
.A1(n_794),
.A2(n_910),
.B(n_772),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_882),
.B(n_867),
.Y(n_1031)
);

OA21x2_ASAP7_75t_L g1032 ( 
.A1(n_853),
.A2(n_832),
.B(n_815),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_810),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_822),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_849),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_936),
.Y(n_1036)
);

INVx4_ASAP7_75t_L g1037 ( 
.A(n_916),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_912),
.B(n_889),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_870),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_827),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_821),
.A2(n_826),
.B(n_915),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_938),
.B(n_843),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_764),
.B(n_889),
.Y(n_1043)
);

AO21x2_ASAP7_75t_L g1044 ( 
.A1(n_934),
.A2(n_850),
.B(n_862),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_774),
.A2(n_814),
.B1(n_834),
.B2(n_846),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_938),
.B(n_890),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_837),
.Y(n_1047)
);

CKINVDCx20_ASAP7_75t_R g1048 ( 
.A(n_938),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_942),
.B(n_938),
.Y(n_1049)
);

BUFx12f_ASAP7_75t_L g1050 ( 
.A(n_942),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_881),
.A2(n_894),
.B(n_920),
.C(n_910),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_890),
.B(n_894),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_917),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_884),
.B(n_838),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_826),
.A2(n_922),
.B(n_927),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_841),
.A2(n_839),
.B1(n_834),
.B2(n_846),
.Y(n_1056)
);

AO22x1_ASAP7_75t_L g1057 ( 
.A1(n_839),
.A2(n_921),
.B1(n_908),
.B2(n_824),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_847),
.B(n_903),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_903),
.Y(n_1059)
);

INVxp33_ASAP7_75t_SL g1060 ( 
.A(n_860),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_904),
.A2(n_907),
.B(n_835),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_814),
.A2(n_906),
.B1(n_929),
.B2(n_945),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_920),
.B(n_943),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_896),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_935),
.A2(n_932),
.B1(n_918),
.B2(n_947),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_SL g1066 ( 
.A1(n_775),
.A2(n_790),
.B(n_792),
.C(n_795),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_857),
.B(n_858),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_L g1068 ( 
.A(n_917),
.B(n_790),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_777),
.A2(n_917),
.B1(n_863),
.B2(n_792),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_874),
.Y(n_1070)
);

AOI22x1_ASAP7_75t_L g1071 ( 
.A1(n_848),
.A2(n_840),
.B1(n_874),
.B2(n_802),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_R g1072 ( 
.A(n_880),
.B(n_885),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_870),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_831),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_933),
.B(n_795),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_833),
.A2(n_803),
.B(n_855),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_948),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_866),
.B(n_808),
.Y(n_1078)
);

CKINVDCx14_ASAP7_75t_R g1079 ( 
.A(n_883),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_866),
.B(n_813),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_859),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_829),
.B(n_825),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_931),
.B(n_928),
.Y(n_1083)
);

NAND3xp33_ASAP7_75t_SL g1084 ( 
.A(n_940),
.B(n_946),
.C(n_941),
.Y(n_1084)
);

BUFx2_ASAP7_75t_R g1085 ( 
.A(n_861),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_864),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_901),
.B(n_886),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_888),
.A2(n_891),
.B(n_893),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_871),
.Y(n_1089)
);

NOR3xp33_ASAP7_75t_L g1090 ( 
.A(n_869),
.B(n_873),
.C(n_900),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_924),
.A2(n_819),
.B1(n_776),
.B2(n_787),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_819),
.A2(n_776),
.B1(n_787),
.B2(n_799),
.Y(n_1092)
);

NAND2x1_ASAP7_75t_L g1093 ( 
.A(n_916),
.B(n_683),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_1043),
.A2(n_989),
.B(n_1052),
.C(n_1005),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_SL g1095 ( 
.A1(n_1092),
.A2(n_982),
.B(n_984),
.C(n_995),
.Y(n_1095)
);

AO31x2_ASAP7_75t_L g1096 ( 
.A1(n_1091),
.A2(n_1011),
.A3(n_1018),
.B(n_1030),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_1038),
.A2(n_970),
.B(n_1056),
.C(n_973),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_SL g1098 ( 
.A1(n_1063),
.A2(n_1046),
.B(n_954),
.C(n_1078),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_975),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_1076),
.A2(n_1088),
.B(n_1071),
.Y(n_1100)
);

AOI221x1_ASAP7_75t_L g1101 ( 
.A1(n_1016),
.A2(n_1007),
.B1(n_1019),
.B2(n_1000),
.C(n_988),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_963),
.A2(n_951),
.B(n_1041),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_1051),
.A2(n_1031),
.B(n_1012),
.C(n_950),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_978),
.Y(n_1104)
);

OR2x2_ASAP7_75t_L g1105 ( 
.A(n_1029),
.B(n_998),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_951),
.A2(n_1041),
.B(n_1067),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_1053),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_958),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_979),
.Y(n_1109)
);

INVx4_ASAP7_75t_L g1110 ( 
.A(n_952),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_1061),
.A2(n_1076),
.A3(n_1055),
.B(n_1015),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_1060),
.B(n_1006),
.Y(n_1112)
);

OA21x2_ASAP7_75t_L g1113 ( 
.A1(n_1027),
.A2(n_1061),
.B(n_1055),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_964),
.B(n_1013),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1051),
.A2(n_949),
.B(n_977),
.C(n_1062),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_1048),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_1053),
.Y(n_1117)
);

AO31x2_ASAP7_75t_L g1118 ( 
.A1(n_1069),
.A2(n_969),
.A3(n_1074),
.B(n_1089),
.Y(n_1118)
);

CKINVDCx11_ASAP7_75t_R g1119 ( 
.A(n_986),
.Y(n_1119)
);

NAND2x1p5_ASAP7_75t_L g1120 ( 
.A(n_952),
.B(n_1037),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_961),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_968),
.A2(n_1087),
.B(n_1086),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_953),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_959),
.B(n_1004),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_993),
.A2(n_1009),
.B(n_974),
.C(n_1042),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_1023),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_SL g1127 ( 
.A(n_1085),
.B(n_999),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1080),
.A2(n_1083),
.B(n_1032),
.Y(n_1128)
);

AO22x2_ASAP7_75t_L g1129 ( 
.A1(n_1000),
.A2(n_1045),
.B1(n_1003),
.B2(n_988),
.Y(n_1129)
);

CKINVDCx11_ASAP7_75t_R g1130 ( 
.A(n_1050),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1032),
.A2(n_1084),
.B(n_968),
.Y(n_1131)
);

CKINVDCx11_ASAP7_75t_R g1132 ( 
.A(n_1036),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_992),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_1014),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_1028),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1057),
.B(n_967),
.Y(n_1136)
);

AO31x2_ASAP7_75t_L g1137 ( 
.A1(n_987),
.A2(n_981),
.A3(n_971),
.B(n_1075),
.Y(n_1137)
);

OAI22x1_ASAP7_75t_L g1138 ( 
.A1(n_1077),
.A2(n_976),
.B1(n_997),
.B2(n_1025),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_949),
.A2(n_1027),
.B(n_962),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1017),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_966),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_960),
.B(n_1020),
.Y(n_1142)
);

NAND3xp33_ASAP7_75t_L g1143 ( 
.A(n_1002),
.B(n_974),
.C(n_1003),
.Y(n_1143)
);

BUFx10_ASAP7_75t_L g1144 ( 
.A(n_1021),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_960),
.B(n_1021),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1084),
.A2(n_1066),
.B(n_1010),
.Y(n_1146)
);

AO31x2_ASAP7_75t_L g1147 ( 
.A1(n_987),
.A2(n_981),
.A3(n_971),
.B(n_983),
.Y(n_1147)
);

INVx4_ASAP7_75t_L g1148 ( 
.A(n_953),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1010),
.A2(n_1081),
.B(n_1044),
.Y(n_1149)
);

NAND3xp33_ASAP7_75t_SL g1150 ( 
.A(n_994),
.B(n_1065),
.C(n_980),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1026),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_962),
.A2(n_965),
.B(n_1081),
.C(n_1079),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_1054),
.A2(n_1047),
.A3(n_1040),
.B(n_991),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_967),
.B(n_1064),
.Y(n_1154)
);

NAND3xp33_ASAP7_75t_L g1155 ( 
.A(n_1090),
.B(n_965),
.C(n_1059),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1010),
.A2(n_1044),
.B(n_1086),
.Y(n_1156)
);

INVx5_ASAP7_75t_L g1157 ( 
.A(n_1053),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1082),
.A2(n_1058),
.B(n_1090),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1008),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_1049),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_956),
.A2(n_1068),
.B(n_1093),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1033),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1034),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1082),
.A2(n_980),
.B(n_1070),
.C(n_996),
.Y(n_1164)
);

INVx8_ASAP7_75t_L g1165 ( 
.A(n_953),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1010),
.A2(n_955),
.B(n_1068),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1049),
.B(n_985),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_972),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1085),
.B(n_985),
.Y(n_1169)
);

INVx4_ASAP7_75t_L g1170 ( 
.A(n_972),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_972),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1022),
.B(n_1024),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_990),
.Y(n_1173)
);

O2A1O1Ixp5_ASAP7_75t_L g1174 ( 
.A1(n_1001),
.A2(n_1073),
.B(n_1039),
.C(n_1035),
.Y(n_1174)
);

NAND3xp33_ASAP7_75t_L g1175 ( 
.A(n_1022),
.B(n_1024),
.C(n_990),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1039),
.A2(n_1073),
.B(n_1035),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1024),
.B(n_1072),
.Y(n_1177)
);

NOR2xp67_ASAP7_75t_L g1178 ( 
.A(n_1037),
.B(n_990),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_957),
.Y(n_1179)
);

AO21x1_ASAP7_75t_L g1180 ( 
.A1(n_1092),
.A2(n_776),
.B(n_1091),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_995),
.B(n_950),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_SL g1182 ( 
.A1(n_989),
.A2(n_819),
.B(n_776),
.C(n_1092),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_989),
.A2(n_776),
.B(n_819),
.C(n_1043),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_995),
.B(n_950),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_975),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_975),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_989),
.A2(n_819),
.B(n_776),
.Y(n_1187)
);

XOR2xp5_ASAP7_75t_L g1188 ( 
.A(n_978),
.B(n_902),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_995),
.B(n_950),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_975),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_957),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1016),
.A2(n_776),
.B1(n_1043),
.B2(n_913),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_963),
.A2(n_1011),
.B(n_989),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_953),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1060),
.B(n_624),
.Y(n_1195)
);

AOI221xp5_ASAP7_75t_L g1196 ( 
.A1(n_1043),
.A2(n_776),
.B1(n_475),
.B2(n_622),
.C(n_1092),
.Y(n_1196)
);

BUFx8_ASAP7_75t_L g1197 ( 
.A(n_986),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_SL g1198 ( 
.A(n_978),
.B(n_672),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1092),
.A2(n_854),
.A3(n_989),
.B(n_1091),
.Y(n_1199)
);

AOI221x1_ASAP7_75t_L g1200 ( 
.A1(n_1092),
.A2(n_776),
.B1(n_819),
.B2(n_989),
.C(n_1091),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_1092),
.A2(n_854),
.A3(n_989),
.B(n_1091),
.Y(n_1201)
);

INVx5_ASAP7_75t_L g1202 ( 
.A(n_1053),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_963),
.A2(n_1011),
.B(n_989),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1092),
.A2(n_854),
.A3(n_989),
.B(n_1091),
.Y(n_1204)
);

INVx5_ASAP7_75t_L g1205 ( 
.A(n_1053),
.Y(n_1205)
);

OR2x6_ASAP7_75t_L g1206 ( 
.A(n_986),
.B(n_565),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_SL g1207 ( 
.A1(n_1016),
.A2(n_1060),
.B1(n_672),
.B2(n_1079),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_963),
.A2(n_1011),
.B(n_989),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_978),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_963),
.A2(n_1011),
.B(n_989),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_963),
.A2(n_1011),
.B(n_989),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1076),
.A2(n_1088),
.B(n_1071),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1049),
.B(n_914),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1076),
.A2(n_1088),
.B(n_1071),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_963),
.A2(n_1011),
.B(n_989),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_963),
.A2(n_1011),
.B(n_989),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1076),
.A2(n_1088),
.B(n_1071),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1076),
.A2(n_1088),
.B(n_1071),
.Y(n_1218)
);

AOI21x1_ASAP7_75t_L g1219 ( 
.A1(n_951),
.A2(n_1041),
.B(n_1011),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_953),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_963),
.A2(n_1011),
.B(n_989),
.Y(n_1221)
);

AOI221x1_ASAP7_75t_L g1222 ( 
.A1(n_1092),
.A2(n_776),
.B1(n_819),
.B2(n_989),
.C(n_1091),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1076),
.A2(n_1088),
.B(n_1071),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_975),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_957),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1076),
.A2(n_1088),
.B(n_1071),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_963),
.A2(n_1011),
.B(n_989),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_957),
.Y(n_1228)
);

INVxp67_ASAP7_75t_L g1229 ( 
.A(n_975),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1049),
.B(n_914),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1076),
.A2(n_1088),
.B(n_1071),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1076),
.A2(n_1088),
.B(n_1071),
.Y(n_1232)
);

INVx3_ASAP7_75t_SL g1233 ( 
.A(n_1104),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1110),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1158),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1120),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1192),
.A2(n_1196),
.B1(n_1195),
.B2(n_1207),
.Y(n_1237)
);

BUFx4f_ASAP7_75t_SL g1238 ( 
.A(n_1209),
.Y(n_1238)
);

BUFx8_ASAP7_75t_SL g1239 ( 
.A(n_1116),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1133),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1225),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1187),
.A2(n_1143),
.B1(n_1127),
.B2(n_1139),
.Y(n_1242)
);

CKINVDCx11_ASAP7_75t_R g1243 ( 
.A(n_1119),
.Y(n_1243)
);

INVx6_ASAP7_75t_L g1244 ( 
.A(n_1157),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1228),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1108),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1179),
.Y(n_1247)
);

BUFx10_ASAP7_75t_L g1248 ( 
.A(n_1112),
.Y(n_1248)
);

BUFx8_ASAP7_75t_L g1249 ( 
.A(n_1186),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1191),
.Y(n_1250)
);

CKINVDCx11_ASAP7_75t_R g1251 ( 
.A(n_1130),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1180),
.A2(n_1150),
.B1(n_1138),
.B2(n_1189),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1140),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1151),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1165),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1162),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1114),
.B(n_1103),
.Y(n_1257)
);

BUFx8_ASAP7_75t_SL g1258 ( 
.A(n_1134),
.Y(n_1258)
);

INVx4_ASAP7_75t_L g1259 ( 
.A(n_1157),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1097),
.A2(n_1152),
.B1(n_1094),
.B2(n_1105),
.Y(n_1260)
);

INVx8_ASAP7_75t_L g1261 ( 
.A(n_1165),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1162),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_SL g1263 ( 
.A1(n_1135),
.A2(n_1169),
.B1(n_1188),
.B2(n_1142),
.Y(n_1263)
);

CKINVDCx12_ASAP7_75t_R g1264 ( 
.A(n_1206),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1129),
.A2(n_1216),
.B1(n_1210),
.B2(n_1211),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_SL g1266 ( 
.A1(n_1129),
.A2(n_1198),
.B1(n_1203),
.B2(n_1193),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1159),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1163),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1099),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1154),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1208),
.A2(n_1215),
.B1(n_1221),
.B2(n_1227),
.Y(n_1271)
);

OAI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1200),
.A2(n_1222),
.B1(n_1101),
.B2(n_1136),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1183),
.A2(n_1109),
.B1(n_1177),
.B2(n_1229),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1124),
.B(n_1145),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1123),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1185),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_1190),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1182),
.A2(n_1141),
.B1(n_1197),
.B2(n_1113),
.Y(n_1278)
);

BUFx2_ASAP7_75t_SL g1279 ( 
.A(n_1202),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1153),
.Y(n_1280)
);

BUFx4f_ASAP7_75t_L g1281 ( 
.A(n_1206),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1197),
.A2(n_1113),
.B1(n_1146),
.B2(n_1155),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1106),
.A2(n_1102),
.B1(n_1128),
.B2(n_1160),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1153),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1224),
.A2(n_1115),
.B1(n_1164),
.B2(n_1125),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1167),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1213),
.A2(n_1230),
.B1(n_1166),
.B2(n_1132),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1144),
.Y(n_1288)
);

BUFx4_ASAP7_75t_SL g1289 ( 
.A(n_1175),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1118),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1213),
.A2(n_1230),
.B1(n_1178),
.B2(n_1205),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1219),
.A2(n_1131),
.B(n_1172),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1144),
.A2(n_1095),
.B1(n_1149),
.B2(n_1117),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1096),
.A2(n_1202),
.B1(n_1205),
.B2(n_1098),
.Y(n_1294)
);

OAI22xp33_ASAP7_75t_R g1295 ( 
.A1(n_1096),
.A2(n_1204),
.B1(n_1199),
.B2(n_1201),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_1202),
.Y(n_1296)
);

INVx6_ASAP7_75t_L g1297 ( 
.A(n_1205),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_SL g1298 ( 
.A1(n_1096),
.A2(n_1201),
.B1(n_1199),
.B2(n_1204),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1107),
.A2(n_1117),
.B1(n_1122),
.B2(n_1156),
.Y(n_1299)
);

OAI22x1_ASAP7_75t_SL g1300 ( 
.A1(n_1148),
.A2(n_1170),
.B1(n_1220),
.B2(n_1171),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1176),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1123),
.Y(n_1302)
);

BUFx12f_ASAP7_75t_L g1303 ( 
.A(n_1168),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1171),
.Y(n_1304)
);

INVx8_ASAP7_75t_L g1305 ( 
.A(n_1171),
.Y(n_1305)
);

OAI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1148),
.A2(n_1170),
.B1(n_1194),
.B2(n_1173),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1174),
.A2(n_1161),
.B(n_1100),
.Y(n_1307)
);

INVx4_ASAP7_75t_L g1308 ( 
.A(n_1194),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1199),
.B(n_1201),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1137),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_1147),
.Y(n_1311)
);

BUFx12f_ASAP7_75t_L g1312 ( 
.A(n_1147),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1212),
.A2(n_1218),
.B1(n_1231),
.B2(n_1214),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1111),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1217),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1223),
.A2(n_776),
.B1(n_1196),
.B2(n_1192),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1226),
.B(n_1232),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1121),
.Y(n_1318)
);

OAI21xp33_ASAP7_75t_L g1319 ( 
.A1(n_1192),
.A2(n_776),
.B(n_1043),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1192),
.A2(n_819),
.B1(n_1060),
.B2(n_1195),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1181),
.B(n_1184),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1121),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1196),
.A2(n_776),
.B1(n_1192),
.B2(n_1016),
.Y(n_1323)
);

OAI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1196),
.A2(n_776),
.B1(n_596),
.B2(n_1200),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1134),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1192),
.A2(n_819),
.B1(n_1060),
.B2(n_1195),
.Y(n_1326)
);

OAI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1196),
.A2(n_776),
.B1(n_596),
.B2(n_1200),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1121),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1121),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1181),
.B(n_1184),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1126),
.Y(n_1331)
);

OAI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1187),
.A2(n_1005),
.B1(n_596),
.B2(n_1043),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1126),
.Y(n_1333)
);

NAND2x1p5_ASAP7_75t_L g1334 ( 
.A(n_1157),
.B(n_1010),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1126),
.Y(n_1335)
);

INVx6_ASAP7_75t_L g1336 ( 
.A(n_1157),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1196),
.A2(n_776),
.B1(n_1192),
.B2(n_1016),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_1209),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_SL g1339 ( 
.A1(n_1207),
.A2(n_1016),
.B1(n_1038),
.B2(n_1043),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_1209),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1196),
.A2(n_776),
.B1(n_1192),
.B2(n_1016),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1126),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1196),
.A2(n_776),
.B1(n_1192),
.B2(n_1016),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1110),
.B(n_1160),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1196),
.A2(n_776),
.B1(n_1192),
.B2(n_1016),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1134),
.Y(n_1346)
);

AND2x2_ASAP7_75t_SL g1347 ( 
.A(n_1265),
.B(n_1323),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1280),
.Y(n_1348)
);

OR2x6_ASAP7_75t_L g1349 ( 
.A(n_1312),
.B(n_1292),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1309),
.B(n_1235),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1284),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1323),
.A2(n_1345),
.B1(n_1337),
.B2(n_1343),
.Y(n_1352)
);

OAI21xp33_ASAP7_75t_SL g1353 ( 
.A1(n_1337),
.A2(n_1343),
.B(n_1341),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1281),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1321),
.B(n_1330),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1235),
.B(n_1298),
.Y(n_1356)
);

NOR2x1_ASAP7_75t_SL g1357 ( 
.A(n_1285),
.B(n_1260),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1324),
.A2(n_1327),
.B(n_1319),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1281),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1290),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1298),
.B(n_1242),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1320),
.B(n_1326),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1239),
.Y(n_1363)
);

AO21x2_ASAP7_75t_L g1364 ( 
.A1(n_1307),
.A2(n_1313),
.B(n_1272),
.Y(n_1364)
);

INVxp67_ASAP7_75t_L g1365 ( 
.A(n_1269),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1271),
.A2(n_1283),
.B(n_1317),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1242),
.B(n_1310),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1311),
.B(n_1256),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1295),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1271),
.A2(n_1283),
.B(n_1315),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1314),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1301),
.B(n_1299),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1262),
.Y(n_1373)
);

BUFx4f_ASAP7_75t_SL g1374 ( 
.A(n_1338),
.Y(n_1374)
);

AO21x2_ASAP7_75t_L g1375 ( 
.A1(n_1272),
.A2(n_1324),
.B(n_1327),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1246),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1247),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1266),
.B(n_1316),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1250),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1253),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1265),
.A2(n_1299),
.B(n_1293),
.Y(n_1381)
);

BUFx2_ASAP7_75t_SL g1382 ( 
.A(n_1296),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1254),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1267),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1257),
.B(n_1286),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1266),
.B(n_1316),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_1276),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1252),
.B(n_1341),
.Y(n_1388)
);

AO21x2_ASAP7_75t_L g1389 ( 
.A1(n_1237),
.A2(n_1270),
.B(n_1306),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1268),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1240),
.B(n_1241),
.Y(n_1391)
);

AO21x2_ASAP7_75t_L g1392 ( 
.A1(n_1306),
.A2(n_1318),
.B(n_1245),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1244),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1274),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1252),
.B(n_1345),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1273),
.B(n_1329),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1328),
.Y(n_1397)
);

BUFx4f_ASAP7_75t_SL g1398 ( 
.A(n_1340),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1322),
.B(n_1339),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1249),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1282),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1334),
.Y(n_1402)
);

OR2x6_ASAP7_75t_L g1403 ( 
.A(n_1279),
.B(n_1291),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1282),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1294),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1294),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1278),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1278),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1249),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1297),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1297),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1293),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1332),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1300),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1339),
.A2(n_1287),
.B(n_1234),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1289),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1277),
.B(n_1346),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1336),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1264),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1263),
.A2(n_1248),
.B1(n_1325),
.B2(n_1344),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1289),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1259),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1352),
.A2(n_1233),
.B1(n_1236),
.B2(n_1238),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1347),
.A2(n_1233),
.B1(n_1238),
.B2(n_1288),
.Y(n_1424)
);

INVxp67_ASAP7_75t_L g1425 ( 
.A(n_1417),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1368),
.B(n_1248),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1355),
.B(n_1258),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1369),
.B(n_1304),
.Y(n_1428)
);

NOR2xp67_ASAP7_75t_L g1429 ( 
.A(n_1419),
.B(n_1308),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1366),
.A2(n_1344),
.B(n_1305),
.Y(n_1430)
);

NOR2x1_ASAP7_75t_SL g1431 ( 
.A(n_1349),
.B(n_1389),
.Y(n_1431)
);

INVx2_ASAP7_75t_SL g1432 ( 
.A(n_1374),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1362),
.A2(n_1261),
.B(n_1335),
.C(n_1333),
.Y(n_1433)
);

NOR2x1_ASAP7_75t_SL g1434 ( 
.A(n_1349),
.B(n_1303),
.Y(n_1434)
);

CKINVDCx20_ASAP7_75t_R g1435 ( 
.A(n_1398),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1369),
.B(n_1304),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1353),
.A2(n_1261),
.B(n_1342),
.C(n_1331),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1357),
.A2(n_1305),
.B(n_1261),
.Y(n_1438)
);

AO21x1_ASAP7_75t_L g1439 ( 
.A1(n_1358),
.A2(n_1308),
.B(n_1305),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1391),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_SL g1441 ( 
.A1(n_1357),
.A2(n_1243),
.B(n_1251),
.Y(n_1441)
);

NOR3xp33_ASAP7_75t_SL g1442 ( 
.A(n_1363),
.B(n_1255),
.C(n_1302),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1376),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1365),
.B(n_1387),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1377),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1347),
.A2(n_1255),
.B1(n_1275),
.B2(n_1358),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1353),
.A2(n_1275),
.B(n_1388),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1350),
.B(n_1394),
.Y(n_1448)
);

A2O1A1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1388),
.A2(n_1395),
.B(n_1386),
.C(n_1378),
.Y(n_1449)
);

AO32x2_ASAP7_75t_L g1450 ( 
.A1(n_1393),
.A2(n_1411),
.A3(n_1410),
.B1(n_1375),
.B2(n_1350),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1413),
.B(n_1379),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1413),
.B(n_1367),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1395),
.A2(n_1386),
.B(n_1378),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1356),
.B(n_1361),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_SL g1455 ( 
.A1(n_1415),
.A2(n_1396),
.B(n_1385),
.Y(n_1455)
);

NOR2x1_ASAP7_75t_SL g1456 ( 
.A(n_1349),
.B(n_1389),
.Y(n_1456)
);

INVx5_ASAP7_75t_SL g1457 ( 
.A(n_1403),
.Y(n_1457)
);

AOI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1401),
.A2(n_1404),
.B1(n_1375),
.B2(n_1412),
.C(n_1399),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1356),
.B(n_1383),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1416),
.B(n_1421),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1383),
.B(n_1373),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1418),
.Y(n_1462)
);

A2O1A1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1381),
.A2(n_1404),
.B(n_1401),
.C(n_1407),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1414),
.A2(n_1405),
.B1(n_1406),
.B2(n_1420),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1373),
.B(n_1384),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1412),
.A2(n_1370),
.B(n_1407),
.Y(n_1466)
);

AO21x1_ASAP7_75t_L g1467 ( 
.A1(n_1408),
.A2(n_1406),
.B(n_1405),
.Y(n_1467)
);

AO32x2_ASAP7_75t_L g1468 ( 
.A1(n_1393),
.A2(n_1411),
.A3(n_1410),
.B1(n_1375),
.B2(n_1364),
.Y(n_1468)
);

AOI21xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1419),
.A2(n_1414),
.B(n_1409),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1382),
.B(n_1354),
.Y(n_1470)
);

AOI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1375),
.A2(n_1408),
.B1(n_1389),
.B2(n_1364),
.C(n_1397),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1384),
.B(n_1380),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1382),
.B(n_1359),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1348),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1390),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_SL g1476 ( 
.A1(n_1402),
.A2(n_1422),
.B(n_1397),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1448),
.B(n_1451),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1459),
.B(n_1364),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1474),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1450),
.B(n_1364),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1445),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1450),
.B(n_1468),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1430),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1465),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1430),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1461),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1472),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1450),
.B(n_1372),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1468),
.B(n_1372),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1468),
.B(n_1372),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1472),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1454),
.B(n_1351),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1466),
.B(n_1371),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1471),
.B(n_1360),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1475),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1440),
.Y(n_1496)
);

INVxp67_ASAP7_75t_L g1497 ( 
.A(n_1476),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1443),
.Y(n_1498)
);

CKINVDCx16_ASAP7_75t_R g1499 ( 
.A(n_1426),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1431),
.Y(n_1500)
);

INVx5_ASAP7_75t_L g1501 ( 
.A(n_1485),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1496),
.Y(n_1502)
);

AOI221xp5_ASAP7_75t_L g1503 ( 
.A1(n_1494),
.A2(n_1464),
.B1(n_1458),
.B2(n_1453),
.C(n_1449),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1499),
.A2(n_1437),
.B1(n_1424),
.B2(n_1423),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1492),
.B(n_1452),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1478),
.B(n_1456),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1492),
.B(n_1452),
.Y(n_1507)
);

OR2x6_ASAP7_75t_L g1508 ( 
.A(n_1500),
.B(n_1349),
.Y(n_1508)
);

OAI31xp33_ASAP7_75t_L g1509 ( 
.A1(n_1494),
.A2(n_1423),
.A3(n_1464),
.B(n_1424),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1478),
.B(n_1457),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1485),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1478),
.B(n_1457),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1495),
.Y(n_1513)
);

INVxp67_ASAP7_75t_SL g1514 ( 
.A(n_1498),
.Y(n_1514)
);

NAND4xp25_ASAP7_75t_L g1515 ( 
.A(n_1480),
.B(n_1453),
.C(n_1463),
.D(n_1444),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1500),
.B(n_1434),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1477),
.B(n_1425),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1479),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1477),
.B(n_1467),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1487),
.B(n_1389),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1479),
.Y(n_1521)
);

NAND4xp25_ASAP7_75t_L g1522 ( 
.A(n_1480),
.B(n_1447),
.C(n_1460),
.D(n_1469),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1486),
.B(n_1462),
.Y(n_1523)
);

NAND4xp25_ASAP7_75t_L g1524 ( 
.A(n_1480),
.B(n_1447),
.C(n_1427),
.D(n_1433),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1481),
.Y(n_1525)
);

AOI221xp5_ASAP7_75t_L g1526 ( 
.A1(n_1482),
.A2(n_1455),
.B1(n_1446),
.B2(n_1428),
.C(n_1436),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1499),
.B(n_1409),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1493),
.A2(n_1349),
.B1(n_1439),
.B2(n_1446),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1487),
.B(n_1428),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1491),
.B(n_1436),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1491),
.B(n_1392),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1518),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1506),
.B(n_1488),
.Y(n_1533)
);

NOR2xp67_ASAP7_75t_L g1534 ( 
.A(n_1501),
.B(n_1497),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1506),
.B(n_1488),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1519),
.B(n_1498),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1501),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1514),
.B(n_1484),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1501),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1518),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1521),
.Y(n_1541)
);

NAND2xp33_ASAP7_75t_R g1542 ( 
.A(n_1527),
.B(n_1442),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1521),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1501),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1529),
.B(n_1484),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1515),
.B(n_1497),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1530),
.B(n_1484),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1511),
.B(n_1489),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1511),
.B(n_1489),
.Y(n_1549)
);

NOR2xp67_ASAP7_75t_L g1550 ( 
.A(n_1501),
.B(n_1500),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1511),
.B(n_1490),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1501),
.B(n_1483),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1511),
.B(n_1490),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1525),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1502),
.Y(n_1555)
);

NAND2x1_ASAP7_75t_SL g1556 ( 
.A(n_1516),
.B(n_1482),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1513),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1523),
.B(n_1490),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1508),
.Y(n_1559)
);

OAI31xp33_ASAP7_75t_L g1560 ( 
.A1(n_1546),
.A2(n_1509),
.A3(n_1522),
.B(n_1504),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1557),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1546),
.B(n_1526),
.Y(n_1562)
);

INVxp67_ASAP7_75t_SL g1563 ( 
.A(n_1556),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1536),
.B(n_1400),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1559),
.B(n_1516),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1554),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1554),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1559),
.B(n_1516),
.Y(n_1568)
);

NAND2x1p5_ASAP7_75t_L g1569 ( 
.A(n_1534),
.B(n_1483),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1559),
.B(n_1516),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1542),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1533),
.B(n_1510),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1532),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1537),
.B(n_1508),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1536),
.B(n_1503),
.Y(n_1575)
);

OR2x6_ASAP7_75t_L g1576 ( 
.A(n_1537),
.B(n_1508),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1532),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1538),
.B(n_1520),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1557),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1556),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1533),
.B(n_1510),
.Y(n_1581)
);

INVxp67_ASAP7_75t_SL g1582 ( 
.A(n_1556),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1545),
.B(n_1515),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1540),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1557),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1545),
.B(n_1517),
.Y(n_1586)
);

OAI31xp33_ASAP7_75t_L g1587 ( 
.A1(n_1555),
.A2(n_1509),
.A3(n_1522),
.B(n_1524),
.Y(n_1587)
);

OAI221xp5_ASAP7_75t_L g1588 ( 
.A1(n_1542),
.A2(n_1524),
.B1(n_1528),
.B2(n_1508),
.C(n_1470),
.Y(n_1588)
);

INVxp67_ASAP7_75t_L g1589 ( 
.A(n_1538),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1533),
.B(n_1535),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1557),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1540),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1535),
.B(n_1512),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1547),
.B(n_1531),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1534),
.B(n_1483),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1537),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1555),
.Y(n_1597)
);

INVxp67_ASAP7_75t_L g1598 ( 
.A(n_1547),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1535),
.B(n_1512),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1558),
.B(n_1505),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1558),
.B(n_1507),
.Y(n_1601)
);

NOR2xp67_ASAP7_75t_SL g1602 ( 
.A(n_1588),
.B(n_1400),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1562),
.B(n_1558),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1563),
.B(n_1582),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1590),
.B(n_1548),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1590),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1560),
.B(n_1548),
.Y(n_1607)
);

OAI31xp33_ASAP7_75t_L g1608 ( 
.A1(n_1560),
.A2(n_1552),
.A3(n_1482),
.B(n_1551),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1583),
.B(n_1541),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1587),
.A2(n_1441),
.B(n_1552),
.Y(n_1610)
);

INVx1_ASAP7_75t_SL g1611 ( 
.A(n_1597),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1575),
.B(n_1548),
.Y(n_1612)
);

INVx2_ASAP7_75t_SL g1613 ( 
.A(n_1565),
.Y(n_1613)
);

NAND2x1p5_ASAP7_75t_L g1614 ( 
.A(n_1580),
.B(n_1537),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1587),
.B(n_1549),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1578),
.B(n_1541),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1571),
.B(n_1435),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1578),
.B(n_1600),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1572),
.B(n_1549),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1572),
.B(n_1549),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1573),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1573),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1580),
.B(n_1550),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1581),
.B(n_1551),
.Y(n_1624)
);

AOI21xp33_ASAP7_75t_SL g1625 ( 
.A1(n_1564),
.A2(n_1432),
.B(n_1473),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1581),
.B(n_1551),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1596),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1601),
.B(n_1586),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1577),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1577),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1596),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1589),
.B(n_1553),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1594),
.B(n_1543),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1594),
.B(n_1543),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1584),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1561),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1622),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1622),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1629),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1611),
.B(n_1598),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1603),
.B(n_1566),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1629),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1630),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1614),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1607),
.B(n_1593),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1630),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1615),
.B(n_1593),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1604),
.B(n_1565),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1635),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1612),
.B(n_1599),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1635),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1610),
.B(n_1569),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1614),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1614),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1604),
.B(n_1568),
.Y(n_1655)
);

AOI32xp33_ASAP7_75t_L g1656 ( 
.A1(n_1613),
.A2(n_1570),
.A3(n_1568),
.B1(n_1599),
.B2(n_1552),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1608),
.A2(n_1569),
.B(n_1595),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_L g1658 ( 
.A(n_1613),
.B(n_1570),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1609),
.B(n_1566),
.Y(n_1659)
);

AND2x2_ASAP7_75t_SL g1660 ( 
.A(n_1617),
.B(n_1539),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1621),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1648),
.B(n_1619),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1656),
.A2(n_1625),
.B(n_1569),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1648),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1640),
.B(n_1602),
.Y(n_1665)
);

OAI21xp33_ASAP7_75t_L g1666 ( 
.A1(n_1647),
.A2(n_1632),
.B(n_1609),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1645),
.B(n_1602),
.Y(n_1667)
);

OAI211xp5_ASAP7_75t_SL g1668 ( 
.A1(n_1652),
.A2(n_1618),
.B(n_1628),
.C(n_1627),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1642),
.Y(n_1669)
);

NOR2x1_ASAP7_75t_L g1670 ( 
.A(n_1652),
.B(n_1658),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1660),
.A2(n_1606),
.B1(n_1628),
.B2(n_1618),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1655),
.A2(n_1606),
.B1(n_1576),
.B2(n_1574),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1642),
.Y(n_1673)
);

NAND2xp33_ASAP7_75t_SL g1674 ( 
.A(n_1655),
.B(n_1641),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1660),
.A2(n_1574),
.B1(n_1576),
.B2(n_1619),
.Y(n_1675)
);

INVx1_ASAP7_75t_SL g1676 ( 
.A(n_1641),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1659),
.Y(n_1677)
);

OAI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1657),
.A2(n_1576),
.B1(n_1574),
.B2(n_1508),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1650),
.B(n_1623),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1644),
.A2(n_1574),
.B1(n_1576),
.B2(n_1620),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1669),
.Y(n_1681)
);

XNOR2xp5_ASAP7_75t_L g1682 ( 
.A(n_1664),
.B(n_1359),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1663),
.A2(n_1574),
.B1(n_1576),
.B2(n_1644),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1670),
.A2(n_1653),
.B1(n_1654),
.B2(n_1620),
.Y(n_1684)
);

OAI21xp33_ASAP7_75t_L g1685 ( 
.A1(n_1667),
.A2(n_1661),
.B(n_1638),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1677),
.B(n_1665),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1662),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1673),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1671),
.A2(n_1654),
.B1(n_1653),
.B2(n_1624),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1676),
.B(n_1637),
.Y(n_1690)
);

AO22x1_ASAP7_75t_L g1691 ( 
.A1(n_1675),
.A2(n_1623),
.B1(n_1649),
.B2(n_1643),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1687),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1690),
.B(n_1674),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_SL g1694 ( 
.A(n_1684),
.B(n_1672),
.C(n_1679),
.Y(n_1694)
);

NOR3xp33_ASAP7_75t_L g1695 ( 
.A(n_1686),
.B(n_1668),
.C(n_1666),
.Y(n_1695)
);

OAI321xp33_ASAP7_75t_L g1696 ( 
.A1(n_1683),
.A2(n_1668),
.A3(n_1678),
.B1(n_1680),
.B2(n_1651),
.C(n_1646),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1681),
.Y(n_1697)
);

AOI211x1_ASAP7_75t_L g1698 ( 
.A1(n_1691),
.A2(n_1639),
.B(n_1643),
.C(n_1649),
.Y(n_1698)
);

AOI211xp5_ASAP7_75t_L g1699 ( 
.A1(n_1689),
.A2(n_1623),
.B(n_1631),
.C(n_1627),
.Y(n_1699)
);

AOI21xp33_ASAP7_75t_L g1700 ( 
.A1(n_1685),
.A2(n_1631),
.B(n_1636),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1688),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1682),
.B(n_1624),
.Y(n_1702)
);

NOR2x1_ASAP7_75t_L g1703 ( 
.A(n_1693),
.B(n_1567),
.Y(n_1703)
);

AOI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1696),
.A2(n_1567),
.B1(n_1636),
.B2(n_1626),
.C(n_1544),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1692),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1695),
.A2(n_1694),
.B(n_1699),
.C(n_1700),
.Y(n_1706)
);

OAI21xp33_ASAP7_75t_L g1707 ( 
.A1(n_1702),
.A2(n_1626),
.B(n_1605),
.Y(n_1707)
);

AOI211xp5_ASAP7_75t_L g1708 ( 
.A1(n_1706),
.A2(n_1705),
.B(n_1707),
.C(n_1704),
.Y(n_1708)
);

NAND4xp25_ASAP7_75t_SL g1709 ( 
.A(n_1703),
.B(n_1701),
.C(n_1697),
.D(n_1698),
.Y(n_1709)
);

AOI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1706),
.A2(n_1539),
.B1(n_1544),
.B2(n_1605),
.C(n_1595),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1703),
.Y(n_1711)
);

AOI211x1_ASAP7_75t_SL g1712 ( 
.A1(n_1706),
.A2(n_1544),
.B(n_1539),
.C(n_1561),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1705),
.Y(n_1713)
);

XNOR2x1_ASAP7_75t_L g1714 ( 
.A(n_1711),
.B(n_1359),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1713),
.Y(n_1715)
);

NAND4xp75_ASAP7_75t_L g1716 ( 
.A(n_1710),
.B(n_1550),
.C(n_1544),
.D(n_1539),
.Y(n_1716)
);

OA22x2_ASAP7_75t_L g1717 ( 
.A1(n_1709),
.A2(n_1712),
.B1(n_1708),
.B2(n_1595),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1711),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1718),
.B(n_1616),
.Y(n_1719)
);

A2O1A1Ixp33_ASAP7_75t_L g1720 ( 
.A1(n_1715),
.A2(n_1717),
.B(n_1595),
.C(n_1714),
.Y(n_1720)
);

NOR2x1p5_ASAP7_75t_L g1721 ( 
.A(n_1716),
.B(n_1616),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1720),
.A2(n_1634),
.B1(n_1633),
.B2(n_1592),
.Y(n_1722)
);

OAI22x1_ASAP7_75t_L g1723 ( 
.A1(n_1722),
.A2(n_1719),
.B1(n_1721),
.B2(n_1552),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1723),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1724),
.Y(n_1725)
);

INVxp67_ASAP7_75t_SL g1726 ( 
.A(n_1725),
.Y(n_1726)
);

AO221x1_ASAP7_75t_L g1727 ( 
.A1(n_1726),
.A2(n_1579),
.B1(n_1561),
.B2(n_1591),
.C(n_1585),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_SL g1728 ( 
.A1(n_1726),
.A2(n_1552),
.B1(n_1591),
.B2(n_1585),
.Y(n_1728)
);

OAI21xp5_ASAP7_75t_SL g1729 ( 
.A1(n_1728),
.A2(n_1727),
.B(n_1634),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1728),
.B(n_1633),
.Y(n_1730)
);

AOI22x1_ASAP7_75t_L g1731 ( 
.A1(n_1729),
.A2(n_1591),
.B1(n_1585),
.B2(n_1579),
.Y(n_1731)
);

AOI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1731),
.A2(n_1730),
.B1(n_1579),
.B2(n_1584),
.C(n_1592),
.Y(n_1732)
);

AOI211xp5_ASAP7_75t_L g1733 ( 
.A1(n_1732),
.A2(n_1429),
.B(n_1438),
.C(n_1422),
.Y(n_1733)
);


endmodule