module fake_jpeg_16161_n_185 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_185);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx12f_ASAP7_75t_SL g36 ( 
.A(n_23),
.Y(n_36)
);

NOR3xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_23),
.C(n_16),
.Y(n_57)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_61),
.B1(n_31),
.B2(n_19),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_49),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_22),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_28),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_30),
.Y(n_77)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_16),
.B1(n_29),
.B2(n_22),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_20),
.C(n_21),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_31),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_32),
.A2(n_29),
.B1(n_20),
.B2(n_21),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_72),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_32),
.B1(n_34),
.B2(n_38),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_75),
.B1(n_76),
.B2(n_59),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_67),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_51),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_68),
.A2(n_71),
.B1(n_44),
.B2(n_60),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_23),
.C(n_15),
.Y(n_70)
);

XNOR2x1_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_15),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_78),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_53),
.B(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_52),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_27),
.B1(n_17),
.B2(n_23),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_53),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_85),
.B(n_90),
.Y(n_110)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_66),
.B(n_45),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_69),
.B(n_70),
.Y(n_104)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_68),
.C(n_79),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_72),
.B1(n_64),
.B2(n_67),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_68),
.B1(n_66),
.B2(n_47),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_50),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_62),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_109),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_112),
.B(n_87),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_93),
.C(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_43),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_89),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_15),
.B(n_44),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_118),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_132),
.Y(n_135)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_107),
.C(n_109),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_125),
.B1(n_128),
.B2(n_131),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_90),
.B(n_92),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_124),
.A2(n_115),
.B1(n_108),
.B2(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_126),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_130),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_88),
.B1(n_81),
.B2(n_59),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_99),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_88),
.B(n_91),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_144),
.C(n_131),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_103),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_136),
.B(n_139),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_103),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_141),
.A2(n_143),
.B1(n_106),
.B2(n_101),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_113),
.B1(n_108),
.B2(n_105),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_114),
.C(n_106),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_125),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_147),
.C(n_149),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_120),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_123),
.B1(n_126),
.B2(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_140),
.Y(n_151)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

NAND2xp33_ASAP7_75t_R g161 ( 
.A(n_153),
.B(n_154),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_141),
.A2(n_14),
.B(n_12),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_155),
.A2(n_9),
.B(n_12),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_156),
.A2(n_142),
.B(n_135),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_160),
.B1(n_164),
.B2(n_152),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_135),
.C(n_30),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_146),
.C(n_149),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_8),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_166),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_164),
.B(n_148),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_168),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_156),
.Y(n_168)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_170),
.A3(n_171),
.B1(n_80),
.B2(n_1),
.C1(n_2),
.C2(n_3),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_158),
.B(n_153),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_173),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_165),
.A2(n_55),
.B1(n_80),
.B2(n_3),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_168),
.A2(n_0),
.B(n_1),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_0),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_166),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_174),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_181),
.A2(n_1),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.C1(n_152),
.C2(n_153),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_180),
.A2(n_177),
.B1(n_173),
.B2(n_5),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_183),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_4),
.Y(n_185)
);


endmodule