module real_aes_2636_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_733;
wire n_552;
wire n_402;
wire n_617;
wire n_602;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_286;
wire n_416;
wire n_410;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_397;
wire n_293;
wire n_358;
wire n_275;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_300;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_312;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_762;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_475;
wire n_554;
wire n_668;
NAND2xp5_ASAP7_75t_L g366 ( .A(n_0), .B(n_367), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_1), .A2(n_240), .B1(n_423), .B2(n_424), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_2), .A2(n_203), .B1(n_418), .B2(n_419), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_3), .A2(n_250), .B1(n_387), .B2(n_433), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_4), .A2(n_149), .B1(n_323), .B2(n_652), .Y(n_651) );
XNOR2x1_ASAP7_75t_L g648 ( .A(n_5), .B(n_649), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_6), .A2(n_93), .B1(n_603), .B2(n_604), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_7), .A2(n_29), .B1(n_376), .B2(n_381), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_8), .A2(n_122), .B1(n_397), .B2(n_398), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_9), .A2(n_220), .B1(n_550), .B2(n_552), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_10), .A2(n_178), .B1(n_357), .B2(n_740), .Y(n_739) );
AO22x2_ASAP7_75t_L g305 ( .A1(n_11), .A2(n_187), .B1(n_295), .B2(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g731 ( .A(n_11), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_12), .A2(n_188), .B1(n_419), .B2(n_454), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_13), .A2(n_120), .B1(n_361), .B2(n_426), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_14), .A2(n_190), .B1(n_341), .B2(n_768), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_15), .A2(n_56), .B1(n_552), .B2(n_643), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_16), .A2(n_735), .B1(n_751), .B2(n_752), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_16), .Y(n_752) );
INVx1_ASAP7_75t_L g621 ( .A(n_17), .Y(n_621) );
INVx1_ASAP7_75t_L g638 ( .A(n_18), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_19), .A2(n_237), .B1(n_423), .B2(n_424), .Y(n_688) );
INVx1_ASAP7_75t_L g617 ( .A(n_20), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g678 ( .A(n_21), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_22), .A2(n_88), .B1(n_395), .B2(n_712), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_23), .A2(n_78), .B1(n_535), .B2(n_536), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_24), .A2(n_180), .B1(n_426), .B2(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_SL g591 ( .A1(n_25), .A2(n_210), .B1(n_375), .B2(n_592), .Y(n_591) );
AO22x2_ASAP7_75t_L g302 ( .A1(n_26), .A2(n_68), .B1(n_295), .B2(n_303), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_26), .B(n_730), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_27), .A2(n_224), .B1(n_345), .B2(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_SL g765 ( .A1(n_28), .A2(n_223), .B1(n_542), .B2(n_748), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_30), .A2(n_126), .B1(n_357), .B2(n_360), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_31), .A2(n_143), .B1(n_375), .B2(n_457), .Y(n_456) );
AO222x2_ASAP7_75t_SL g484 ( .A1(n_32), .A2(n_49), .B1(n_159), .B2(n_411), .C1(n_463), .C2(n_464), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_33), .A2(n_160), .B1(n_353), .B2(n_354), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_34), .A2(n_222), .B1(n_431), .B2(n_450), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_35), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_36), .A2(n_89), .B1(n_426), .B2(n_427), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_37), .A2(n_164), .B1(n_473), .B2(n_476), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_38), .A2(n_151), .B1(n_454), .B2(n_467), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_39), .A2(n_48), .B1(n_384), .B2(n_386), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_40), .A2(n_69), .B1(n_384), .B2(n_604), .Y(n_710) );
AOI22xp33_ASAP7_75t_SL g588 ( .A1(n_41), .A2(n_63), .B1(n_373), .B2(n_589), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g317 ( .A1(n_42), .A2(n_166), .B1(n_318), .B2(n_323), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_43), .A2(n_154), .B1(n_427), .B2(n_433), .Y(n_685) );
OA22x2_ASAP7_75t_L g755 ( .A1(n_44), .A2(n_756), .B1(n_757), .B2(n_775), .Y(n_755) );
INVx1_ASAP7_75t_L g775 ( .A(n_44), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_45), .A2(n_137), .B1(n_360), .B2(n_663), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_46), .A2(n_85), .B1(n_313), .B2(n_380), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_47), .A2(n_134), .B1(n_423), .B2(n_424), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_50), .A2(n_182), .B1(n_431), .B2(n_450), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_51), .A2(n_79), .B1(n_424), .B2(n_515), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_52), .A2(n_146), .B1(n_394), .B2(n_606), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_53), .A2(n_115), .B1(n_703), .B2(n_704), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_54), .A2(n_227), .B1(n_594), .B2(n_595), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_55), .A2(n_251), .B1(n_536), .B2(n_599), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_57), .A2(n_99), .B1(n_415), .B2(n_488), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_58), .A2(n_135), .B1(n_389), .B2(n_392), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_59), .A2(n_116), .B1(n_419), .B2(n_454), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_60), .A2(n_179), .B1(n_535), .B2(n_743), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_61), .A2(n_244), .B1(n_529), .B2(n_531), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_62), .A2(n_248), .B1(n_355), .B2(n_426), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_64), .A2(n_167), .B1(n_430), .B2(n_431), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_65), .A2(n_129), .B1(n_415), .B2(n_488), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_66), .A2(n_74), .B1(n_663), .B2(n_743), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_67), .A2(n_147), .B1(n_411), .B2(n_464), .Y(n_671) );
AOI22xp33_ASAP7_75t_SL g466 ( .A1(n_70), .A2(n_112), .B1(n_418), .B2(n_467), .Y(n_466) );
AO222x2_ASAP7_75t_SL g462 ( .A1(n_71), .A2(n_183), .B1(n_199), .B2(n_411), .C1(n_463), .C2(n_464), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_72), .A2(n_157), .B1(n_357), .B2(n_386), .Y(n_533) );
OA22x2_ASAP7_75t_L g666 ( .A1(n_73), .A2(n_667), .B1(n_668), .B2(n_689), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_73), .Y(n_667) );
INVx3_ASAP7_75t_L g295 ( .A(n_75), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_76), .A2(n_106), .B1(n_389), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_77), .A2(n_256), .B1(n_339), .B2(n_341), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_80), .A2(n_140), .B1(n_430), .B2(n_431), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_81), .A2(n_193), .B1(n_427), .B2(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_82), .A2(n_231), .B1(n_411), .B2(n_464), .Y(n_510) );
INVx1_ASAP7_75t_L g630 ( .A(n_83), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_84), .A2(n_185), .B1(n_542), .B2(n_748), .Y(n_747) );
AOI222xp33_ASAP7_75t_L g571 ( .A1(n_86), .A2(n_104), .B1(n_189), .B2(n_412), .C1(n_572), .C2(n_573), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_87), .A2(n_96), .B1(n_329), .B2(n_333), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_90), .A2(n_118), .B1(n_524), .B2(n_527), .Y(n_523) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_91), .A2(n_699), .B1(n_714), .B2(n_715), .Y(n_698) );
INVx1_ASAP7_75t_L g714 ( .A(n_91), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_92), .A2(n_158), .B1(n_595), .B2(n_643), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_94), .A2(n_162), .B1(n_370), .B2(n_373), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_95), .A2(n_123), .B1(n_419), .B2(n_454), .Y(n_453) );
INVx1_ASAP7_75t_SL g296 ( .A(n_97), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_97), .B(n_131), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_98), .A2(n_103), .B1(n_426), .B2(n_427), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_100), .A2(n_133), .B1(n_329), .B2(n_333), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_101), .A2(n_175), .B1(n_654), .B2(n_655), .Y(n_653) );
INVx2_ASAP7_75t_L g280 ( .A(n_102), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_105), .A2(n_266), .B1(n_444), .B2(n_560), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_107), .A2(n_214), .B1(n_415), .B2(n_416), .Y(n_468) );
AOI222xp33_ASAP7_75t_L g759 ( .A1(n_108), .A2(n_125), .B1(n_249), .B2(n_376), .C1(n_760), .C2(n_762), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_109), .A2(n_136), .B1(n_411), .B2(n_412), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_110), .A2(n_144), .B1(n_430), .B2(n_431), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_111), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_113), .A2(n_139), .B1(n_329), .B2(n_592), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_114), .A2(n_181), .B1(n_529), .B2(n_531), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_117), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_119), .A2(n_236), .B1(n_372), .B2(n_373), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_121), .A2(n_238), .B1(n_333), .B2(n_550), .Y(n_570) );
XNOR2x1_ASAP7_75t_SL g581 ( .A(n_124), .B(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_SL g422 ( .A1(n_127), .A2(n_176), .B1(n_423), .B2(n_424), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_128), .A2(n_243), .B1(n_308), .B2(n_313), .Y(n_307) );
INVx1_ASAP7_75t_L g554 ( .A(n_130), .Y(n_554) );
AO22x2_ASAP7_75t_L g298 ( .A1(n_131), .A2(n_202), .B1(n_295), .B2(n_299), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_132), .A2(n_152), .B1(n_542), .B2(n_544), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_138), .A2(n_219), .B1(n_427), .B2(n_433), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_141), .A2(n_263), .B1(n_345), .B2(n_348), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_142), .A2(n_184), .B1(n_373), .B2(n_589), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_145), .A2(n_268), .B1(n_390), .B2(n_560), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_148), .A2(n_255), .B1(n_625), .B2(n_770), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_150), .A2(n_213), .B1(n_375), .B2(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g297 ( .A(n_153), .Y(n_297) );
INVx1_ASAP7_75t_L g640 ( .A(n_155), .Y(n_640) );
CKINVDCx20_ASAP7_75t_R g674 ( .A(n_156), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_161), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_163), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_165), .A2(n_221), .B1(n_565), .B2(n_566), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_168), .A2(n_246), .B1(n_345), .B2(n_660), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_169), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_170), .A2(n_253), .B1(n_643), .B2(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_171), .B(n_368), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_172), .B(n_368), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_173), .A2(n_254), .B1(n_547), .B2(n_548), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_174), .B(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_177), .A2(n_232), .B1(n_394), .B2(n_395), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_186), .A2(n_252), .B1(n_341), .B2(n_444), .Y(n_443) );
XNOR2x1_ASAP7_75t_L g612 ( .A(n_191), .B(n_613), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_192), .A2(n_197), .B1(n_433), .B2(n_476), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_194), .A2(n_217), .B1(n_361), .B2(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_195), .B(n_367), .Y(n_749) );
AOI22xp33_ASAP7_75t_SL g414 ( .A1(n_196), .A2(n_204), .B1(n_415), .B2(n_416), .Y(n_414) );
AOI221x1_ASAP7_75t_L g624 ( .A1(n_198), .A2(n_225), .B1(n_536), .B2(n_625), .C(n_626), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_200), .A2(n_201), .B1(n_547), .B2(n_548), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_205), .B(n_586), .Y(n_657) );
INVx1_ASAP7_75t_L g616 ( .A(n_206), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_207), .A2(n_269), .B1(n_536), .B2(n_603), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_208), .A2(n_257), .B1(n_562), .B2(n_773), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_209), .A2(n_212), .B1(n_526), .B2(n_660), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_211), .A2(n_234), .B1(n_389), .B2(n_392), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_215), .A2(n_265), .B1(n_426), .B2(n_427), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_216), .B(n_368), .Y(n_706) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_218), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g727 ( .A(n_218), .Y(n_727) );
INVx1_ASAP7_75t_L g276 ( .A(n_226), .Y(n_276) );
AND2x2_ASAP7_75t_R g754 ( .A(n_226), .B(n_727), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_228), .B(n_572), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_229), .B(n_289), .Y(n_288) );
XNOR2xp5_ASAP7_75t_L g363 ( .A(n_230), .B(n_364), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_233), .A2(n_264), .B1(n_433), .B2(n_434), .Y(n_432) );
INVxp67_ASAP7_75t_L g278 ( .A(n_235), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_239), .Y(n_680) );
INVx1_ASAP7_75t_L g629 ( .A(n_241), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_242), .A2(n_262), .B1(n_430), .B2(n_431), .Y(n_477) );
INVx1_ASAP7_75t_L g620 ( .A(n_245), .Y(n_620) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_247), .A2(n_271), .B(n_281), .C(n_733), .Y(n_270) );
INVx1_ASAP7_75t_L g633 ( .A(n_258), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_259), .B(n_368), .Y(n_409) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_260), .A2(n_557), .B(n_575), .Y(n_556) );
INVx1_ASAP7_75t_L g577 ( .A(n_260), .Y(n_577) );
INVx1_ASAP7_75t_L g362 ( .A(n_261), .Y(n_362) );
AOI22x1_ASAP7_75t_L g459 ( .A1(n_267), .A2(n_460), .B1(n_478), .B2(n_479), .Y(n_459) );
INVx1_ASAP7_75t_L g479 ( .A(n_267), .Y(n_479) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_273), .Y(n_272) );
AND2x4_ASAP7_75t_SL g273 ( .A(n_274), .B(n_277), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g781 ( .A(n_275), .B(n_277), .Y(n_781) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_276), .B(n_727), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_501), .B1(n_722), .B2(n_723), .C(n_724), .Y(n_281) );
INVx1_ASAP7_75t_L g723 ( .A(n_282), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_403), .B1(n_499), .B2(n_500), .Y(n_282) );
CKINVDCx11_ASAP7_75t_R g499 ( .A(n_283), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_363), .B1(n_401), .B2(n_402), .Y(n_283) );
INVx1_ASAP7_75t_L g401 ( .A(n_284), .Y(n_401) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
XNOR2x1_ASAP7_75t_L g285 ( .A(n_286), .B(n_362), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_337), .Y(n_286) );
NAND4xp25_ASAP7_75t_L g287 ( .A(n_288), .B(n_307), .C(n_317), .D(n_328), .Y(n_287) );
INVx3_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx4_ASAP7_75t_SL g368 ( .A(n_290), .Y(n_368) );
BUFx2_ASAP7_75t_L g540 ( .A(n_290), .Y(n_540) );
INVx4_ASAP7_75t_SL g586 ( .A(n_290), .Y(n_586) );
INVx3_ASAP7_75t_SL g636 ( .A(n_290), .Y(n_636) );
INVx6_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_300), .Y(n_291) );
AND2x4_ASAP7_75t_L g315 ( .A(n_292), .B(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g334 ( .A(n_292), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g416 ( .A(n_292), .B(n_335), .Y(n_416) );
AND2x2_ASAP7_75t_L g419 ( .A(n_292), .B(n_316), .Y(n_419) );
AND2x4_ASAP7_75t_L g463 ( .A(n_292), .B(n_300), .Y(n_463) );
AND2x2_ASAP7_75t_L g467 ( .A(n_292), .B(n_316), .Y(n_467) );
AND2x2_ASAP7_75t_L g488 ( .A(n_292), .B(n_335), .Y(n_488) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_298), .Y(n_292) );
INVx2_ASAP7_75t_L g312 ( .A(n_293), .Y(n_312) );
AND2x2_ASAP7_75t_L g321 ( .A(n_293), .B(n_322), .Y(n_321) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_293), .Y(n_327) );
OAI22x1_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_295), .B1(n_296), .B2(n_297), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g299 ( .A(n_295), .Y(n_299) );
INVx2_ASAP7_75t_L g303 ( .A(n_295), .Y(n_303) );
INVx1_ASAP7_75t_L g306 ( .A(n_295), .Y(n_306) );
AND2x2_ASAP7_75t_L g311 ( .A(n_298), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g322 ( .A(n_298), .Y(n_322) );
BUFx2_ASAP7_75t_L g343 ( .A(n_298), .Y(n_343) );
AND2x2_ASAP7_75t_L g347 ( .A(n_300), .B(n_311), .Y(n_347) );
AND2x4_ASAP7_75t_L g353 ( .A(n_300), .B(n_321), .Y(n_353) );
AND2x4_ASAP7_75t_L g359 ( .A(n_300), .B(n_351), .Y(n_359) );
AND2x2_ASAP7_75t_L g430 ( .A(n_300), .B(n_321), .Y(n_430) );
AND2x6_ASAP7_75t_L g433 ( .A(n_300), .B(n_311), .Y(n_433) );
AND2x2_ASAP7_75t_L g450 ( .A(n_300), .B(n_321), .Y(n_450) );
AND2x2_ASAP7_75t_L g473 ( .A(n_300), .B(n_351), .Y(n_473) );
AND2x4_ASAP7_75t_L g300 ( .A(n_301), .B(n_304), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x4_ASAP7_75t_L g310 ( .A(n_302), .B(n_304), .Y(n_310) );
AND2x2_ASAP7_75t_L g326 ( .A(n_302), .B(n_305), .Y(n_326) );
INVx1_ASAP7_75t_L g332 ( .A(n_302), .Y(n_332) );
INVxp67_ASAP7_75t_L g316 ( .A(n_304), .Y(n_316) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g331 ( .A(n_305), .B(n_332), .Y(n_331) );
BUFx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_309), .Y(n_381) );
BUFx3_ASAP7_75t_L g654 ( .A(n_309), .Y(n_654) );
BUFx2_ASAP7_75t_L g703 ( .A(n_309), .Y(n_703) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AND2x2_ASAP7_75t_L g320 ( .A(n_310), .B(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g361 ( .A(n_310), .B(n_351), .Y(n_361) );
AND2x4_ASAP7_75t_L g411 ( .A(n_310), .B(n_321), .Y(n_411) );
AND2x2_ASAP7_75t_L g418 ( .A(n_310), .B(n_311), .Y(n_418) );
AND2x2_ASAP7_75t_L g454 ( .A(n_310), .B(n_311), .Y(n_454) );
AND2x2_ASAP7_75t_L g476 ( .A(n_310), .B(n_351), .Y(n_476) );
AND2x2_ASAP7_75t_L g340 ( .A(n_311), .B(n_331), .Y(n_340) );
AND2x2_ASAP7_75t_SL g423 ( .A(n_311), .B(n_331), .Y(n_423) );
AND2x2_ASAP7_75t_L g515 ( .A(n_311), .B(n_331), .Y(n_515) );
AND2x4_ASAP7_75t_L g351 ( .A(n_312), .B(n_322), .Y(n_351) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g548 ( .A(n_314), .Y(n_548) );
INVx2_ASAP7_75t_L g595 ( .A(n_314), .Y(n_595) );
INVx2_ASAP7_75t_L g655 ( .A(n_314), .Y(n_655) );
INVx2_ASAP7_75t_SL g704 ( .A(n_314), .Y(n_704) );
INVx2_ASAP7_75t_SL g746 ( .A(n_314), .Y(n_746) );
INVx6_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g639 ( .A(n_318), .Y(n_639) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g652 ( .A(n_319), .Y(n_652) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx3_ASAP7_75t_L g372 ( .A(n_320), .Y(n_372) );
BUFx3_ASAP7_75t_L g543 ( .A(n_320), .Y(n_543) );
BUFx5_ASAP7_75t_L g589 ( .A(n_320), .Y(n_589) );
AND2x2_ASAP7_75t_L g330 ( .A(n_321), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g415 ( .A(n_321), .B(n_331), .Y(n_415) );
BUFx2_ASAP7_75t_L g748 ( .A(n_323), .Y(n_748) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx3_ASAP7_75t_L g545 ( .A(n_324), .Y(n_545) );
INVx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx12f_ASAP7_75t_L g373 ( .A(n_325), .Y(n_373) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x4_ASAP7_75t_L g342 ( .A(n_326), .B(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g355 ( .A(n_326), .B(n_351), .Y(n_355) );
AND2x2_ASAP7_75t_SL g412 ( .A(n_326), .B(n_327), .Y(n_412) );
AND2x4_ASAP7_75t_L g424 ( .A(n_326), .B(n_343), .Y(n_424) );
AND2x4_ASAP7_75t_L g431 ( .A(n_326), .B(n_351), .Y(n_431) );
AND2x2_ASAP7_75t_SL g464 ( .A(n_326), .B(n_327), .Y(n_464) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_330), .Y(n_375) );
INVx3_ASAP7_75t_L g551 ( .A(n_330), .Y(n_551) );
AND2x4_ASAP7_75t_L g350 ( .A(n_331), .B(n_351), .Y(n_350) );
AND2x6_ASAP7_75t_L g427 ( .A(n_331), .B(n_351), .Y(n_427) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_332), .Y(n_336) );
BUFx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g378 ( .A(n_334), .Y(n_378) );
BUFx6f_ASAP7_75t_SL g457 ( .A(n_334), .Y(n_457) );
INVx1_ASAP7_75t_L g553 ( .A(n_334), .Y(n_553) );
BUFx4f_ASAP7_75t_L g592 ( .A(n_334), .Y(n_592) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND4xp25_ASAP7_75t_L g337 ( .A(n_338), .B(n_344), .C(n_352), .D(n_356), .Y(n_337) );
BUFx2_ASAP7_75t_L g768 ( .A(n_339), .Y(n_768) );
BUFx3_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g391 ( .A(n_340), .Y(n_391) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_340), .Y(n_444) );
BUFx3_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx2_ASAP7_75t_L g392 ( .A(n_342), .Y(n_392) );
INVx5_ASAP7_75t_SL g532 ( .A(n_342), .Y(n_532) );
BUFx2_ASAP7_75t_L g709 ( .A(n_342), .Y(n_709) );
INVx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_SL g394 ( .A(n_346), .Y(n_394) );
INVx2_ASAP7_75t_SL g712 ( .A(n_346), .Y(n_712) );
INVx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx2_ASAP7_75t_L g526 ( .A(n_347), .Y(n_526) );
BUFx2_ASAP7_75t_L g774 ( .A(n_347), .Y(n_774) );
INVx2_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g395 ( .A(n_349), .Y(n_395) );
INVx2_ASAP7_75t_L g527 ( .A(n_349), .Y(n_527) );
INVx2_ASAP7_75t_L g562 ( .A(n_349), .Y(n_562) );
INVx2_ASAP7_75t_SL g606 ( .A(n_349), .Y(n_606) );
INVx2_ASAP7_75t_L g660 ( .A(n_349), .Y(n_660) );
INVx8_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx6_ASAP7_75t_L g385 ( .A(n_353), .Y(n_385) );
BUFx3_ASAP7_75t_L g565 ( .A(n_353), .Y(n_565) );
BUFx6f_ASAP7_75t_L g743 ( .A(n_354), .Y(n_743) );
BUFx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_SL g397 ( .A(n_355), .Y(n_397) );
BUFx2_ASAP7_75t_SL g536 ( .A(n_355), .Y(n_536) );
BUFx3_ASAP7_75t_L g665 ( .A(n_355), .Y(n_665) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx4_ASAP7_75t_L g400 ( .A(n_358), .Y(n_400) );
INVx3_ASAP7_75t_L g426 ( .A(n_358), .Y(n_426) );
INVx3_ASAP7_75t_SL g625 ( .A(n_358), .Y(n_625) );
INVx8_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_361), .Y(n_387) );
INVx2_ASAP7_75t_L g435 ( .A(n_361), .Y(n_435) );
BUFx3_ASAP7_75t_L g604 ( .A(n_361), .Y(n_604) );
INVxp67_ASAP7_75t_SL g402 ( .A(n_363), .Y(n_402) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_382), .Y(n_364) );
NAND4xp25_ASAP7_75t_L g365 ( .A(n_366), .B(n_369), .C(n_374), .D(n_379), .Y(n_365) );
BUFx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g637 ( .A(n_373), .Y(n_637) );
BUFx6f_ASAP7_75t_SL g643 ( .A(n_375), .Y(n_643) );
INVx1_ASAP7_75t_L g675 ( .A(n_375), .Y(n_675) );
INVx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx2_ASAP7_75t_L g547 ( .A(n_381), .Y(n_547) );
BUFx4f_ASAP7_75t_SL g594 ( .A(n_381), .Y(n_594) );
NAND4xp25_ASAP7_75t_L g382 ( .A(n_383), .B(n_388), .C(n_393), .D(n_396), .Y(n_382) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g535 ( .A(n_385), .Y(n_535) );
INVx2_ASAP7_75t_L g599 ( .A(n_385), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_385), .A2(n_620), .B1(n_621), .B2(n_622), .Y(n_619) );
INVx3_ASAP7_75t_L g663 ( .A(n_385), .Y(n_663) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g628 ( .A(n_390), .Y(n_628) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g530 ( .A(n_391), .Y(n_530) );
INVx1_ASAP7_75t_L g618 ( .A(n_395), .Y(n_618) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_400), .Y(n_603) );
INVx1_ASAP7_75t_L g500 ( .A(n_403), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_437), .B2(n_498), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
XOR2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_436), .Y(n_405) );
NAND2x1_ASAP7_75t_L g406 ( .A(n_407), .B(n_420), .Y(n_406) );
NOR2x1_ASAP7_75t_L g407 ( .A(n_408), .B(n_413), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_SL g574 ( .A(n_411), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_417), .Y(n_413) );
NOR2x1_ASAP7_75t_L g420 ( .A(n_421), .B(n_428), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_425), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_432), .Y(n_428) );
INVx1_ASAP7_75t_L g448 ( .A(n_433), .Y(n_448) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g566 ( .A(n_435), .Y(n_566) );
INVx1_ASAP7_75t_L g770 ( .A(n_435), .Y(n_770) );
INVx1_ASAP7_75t_L g498 ( .A(n_437), .Y(n_498) );
XNOR2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_458), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
XNOR2x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_451), .Y(n_441) );
NAND4xp25_ASAP7_75t_L g442 ( .A(n_443), .B(n_445), .C(n_446), .D(n_449), .Y(n_442) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND4xp25_ASAP7_75t_SL g451 ( .A(n_452), .B(n_453), .C(n_455), .D(n_456), .Y(n_451) );
INVxp67_ASAP7_75t_L g679 ( .A(n_454), .Y(n_679) );
AO22x2_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_480), .B1(n_481), .B2(n_497), .Y(n_458) );
INVx1_ASAP7_75t_L g497 ( .A(n_459), .Y(n_497) );
INVx1_ASAP7_75t_L g478 ( .A(n_460), .Y(n_478) );
NAND2x1_ASAP7_75t_SL g460 ( .A(n_461), .B(n_469), .Y(n_460) );
NOR2xp67_ASAP7_75t_L g461 ( .A(n_462), .B(n_465), .Y(n_461) );
BUFx2_ASAP7_75t_L g572 ( .A(n_463), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .Y(n_465) );
INVxp67_ASAP7_75t_L g681 ( .A(n_467), .Y(n_681) );
NOR2x1_ASAP7_75t_L g469 ( .A(n_470), .B(n_474), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .Y(n_474) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
XOR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_496), .Y(n_481) );
NAND2x1_ASAP7_75t_L g482 ( .A(n_483), .B(n_489), .Y(n_482) );
NOR2x1_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
NOR2x1_ASAP7_75t_L g489 ( .A(n_490), .B(n_493), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g722 ( .A(n_501), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_609), .B1(n_720), .B2(n_721), .Y(n_501) );
INVx1_ASAP7_75t_L g720 ( .A(n_502), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_580), .B1(n_607), .B2(n_608), .Y(n_502) );
INVx1_ASAP7_75t_L g608 ( .A(n_503), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_555), .B1(n_578), .B2(n_579), .Y(n_503) );
INVx1_ASAP7_75t_L g578 ( .A(n_504), .Y(n_578) );
XOR2x1_ASAP7_75t_L g504 ( .A(n_505), .B(n_520), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
XNOR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_519), .Y(n_506) );
NOR2x1_ASAP7_75t_L g507 ( .A(n_508), .B(n_513), .Y(n_507) );
NAND4xp25_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .C(n_511), .D(n_512), .Y(n_508) );
NAND4xp25_ASAP7_75t_L g513 ( .A(n_514), .B(n_516), .C(n_517), .D(n_518), .Y(n_513) );
XOR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_554), .Y(n_520) );
NOR2x1_ASAP7_75t_L g521 ( .A(n_522), .B(n_537), .Y(n_521) );
NAND4xp25_ASAP7_75t_L g522 ( .A(n_523), .B(n_528), .C(n_533), .D(n_534), .Y(n_522) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_525), .A2(n_616), .B1(n_617), .B2(n_618), .Y(n_615) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g560 ( .A(n_532), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_532), .A2(n_627), .B1(n_629), .B2(n_630), .Y(n_626) );
NAND4xp25_ASAP7_75t_L g537 ( .A(n_538), .B(n_541), .C(n_546), .D(n_549), .Y(n_537) );
INVx2_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx4_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_553), .A2(n_674), .B1(n_675), .B2(n_676), .Y(n_673) );
INVx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_556), .Y(n_579) );
NOR2x1_ASAP7_75t_SL g575 ( .A(n_557), .B(n_576), .Y(n_575) );
NAND4xp75_ASAP7_75t_L g557 ( .A(n_558), .B(n_563), .C(n_568), .D(n_571), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_567), .Y(n_563) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_566), .Y(n_740) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g607 ( .A(n_580), .Y(n_607) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_596), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_590), .Y(n_583) );
OAI21xp33_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_587), .B(n_588), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_601), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_605), .Y(n_601) );
BUFx2_ASAP7_75t_L g623 ( .A(n_604), .Y(n_623) );
INVx1_ASAP7_75t_L g721 ( .A(n_609), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_693), .B1(n_718), .B2(n_719), .Y(n_609) );
INVx1_ASAP7_75t_L g719 ( .A(n_610), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_645), .B1(n_646), .B2(n_691), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g692 ( .A(n_612), .Y(n_692) );
NAND3xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_624), .C(n_631), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_619), .Y(n_614) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_641), .Y(n_631) );
OAI222xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B1(n_637), .B2(n_638), .C1(n_639), .C2(n_640), .Y(n_632) );
INVx3_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g761 ( .A(n_636), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AO22x2_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B1(n_666), .B2(n_690), .Y(n_646) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_658), .Y(n_649) );
NAND4xp25_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .C(n_656), .D(n_657), .Y(n_650) );
INVx1_ASAP7_75t_L g763 ( .A(n_654), .Y(n_763) );
NAND4xp25_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .C(n_662), .D(n_664), .Y(n_658) );
INVx2_ASAP7_75t_L g690 ( .A(n_666), .Y(n_690) );
INVx1_ASAP7_75t_L g717 ( .A(n_666), .Y(n_717) );
INVx1_ASAP7_75t_L g689 ( .A(n_668), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_682), .Y(n_668) );
NOR3xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_673), .C(n_677), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_671), .B(n_672), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_680), .B2(n_681), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_683), .B(n_686), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
INVx2_ASAP7_75t_L g695 ( .A(n_690), .Y(n_695) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g718 ( .A(n_693), .Y(n_718) );
OA21x2_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B(n_716), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_698), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g715 ( .A(n_699), .Y(n_715) );
NOR2xp67_ASAP7_75t_L g699 ( .A(n_700), .B(n_707), .Y(n_699) );
NAND4xp25_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .C(n_705), .D(n_706), .Y(n_700) );
NAND4xp25_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .C(n_711), .D(n_713), .Y(n_707) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_726), .B(n_729), .Y(n_778) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
OAI222xp33_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_753), .B1(n_755), .B2(n_775), .C1(n_776), .C2(n_779), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_735), .Y(n_751) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NOR2xp67_ASAP7_75t_L g736 ( .A(n_737), .B(n_744), .Y(n_736) );
NAND4xp25_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .C(n_741), .D(n_742), .Y(n_737) );
NAND4xp25_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .C(n_749), .D(n_750), .Y(n_744) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
OR2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_766), .Y(n_757) );
NAND3xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_764), .C(n_765), .Y(n_758) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NAND4xp25_ASAP7_75t_L g766 ( .A(n_767), .B(n_769), .C(n_771), .D(n_772), .Y(n_766) );
BUFx3_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
CKINVDCx6p67_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_780), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_781), .Y(n_780) );
endmodule