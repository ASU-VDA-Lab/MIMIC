module fake_jpeg_19920_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_15),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_48),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_22),
.B1(n_23),
.B2(n_32),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_38),
.B1(n_39),
.B2(n_23),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_22),
.B1(n_33),
.B2(n_32),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_64),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_22),
.B1(n_23),
.B2(n_34),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_52),
.B1(n_64),
.B2(n_53),
.Y(n_83)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_26),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_66),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_25),
.B(n_20),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_38),
.B1(n_43),
.B2(n_35),
.Y(n_81)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_33),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_69),
.B(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_46),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_75),
.B(n_78),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_39),
.B1(n_38),
.B2(n_21),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_42),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_79),
.B(n_80),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_46),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_20),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_42),
.B(n_41),
.C(n_37),
.Y(n_82)
);

AO21x1_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_45),
.B(n_51),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_85),
.B1(n_61),
.B2(n_63),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_86),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_43),
.B1(n_35),
.B2(n_27),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_69),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_42),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_90),
.C(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_42),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_53),
.A2(n_55),
.B1(n_64),
.B2(n_57),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_95),
.B1(n_97),
.B2(n_28),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_41),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_41),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_49),
.C(n_20),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_53),
.A2(n_41),
.B1(n_31),
.B2(n_34),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_55),
.A2(n_21),
.B1(n_27),
.B2(n_31),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_99),
.A2(n_91),
.B(n_95),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_100),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_103),
.A2(n_67),
.B1(n_51),
.B2(n_24),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_111),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_105),
.A2(n_114),
.B(n_20),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_76),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_112),
.B(n_119),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_26),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_30),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_117),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_93),
.Y(n_148)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_97),
.B1(n_83),
.B2(n_114),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_89),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_121),
.B(n_80),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_124),
.A2(n_84),
.B1(n_68),
.B2(n_125),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_126),
.A2(n_133),
.B1(n_139),
.B2(n_150),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_128),
.B(n_135),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_119),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_131),
.B(n_142),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_68),
.B1(n_79),
.B2(n_82),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_71),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_154),
.B1(n_156),
.B2(n_16),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_137),
.B(n_144),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_106),
.A2(n_82),
.B1(n_88),
.B2(n_78),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_75),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_140),
.B(n_149),
.C(n_16),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_81),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_141),
.A2(n_146),
.B(n_155),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_102),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_18),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_17),
.B(n_30),
.C(n_28),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_12),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_123),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_92),
.C(n_90),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_87),
.B1(n_61),
.B2(n_49),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_116),
.B(n_18),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_152),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_102),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_67),
.B1(n_24),
.B2(n_17),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_105),
.A2(n_20),
.B1(n_29),
.B2(n_3),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_99),
.B(n_114),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_158),
.A2(n_133),
.B(n_144),
.Y(n_197)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_165),
.Y(n_198)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_105),
.B(n_112),
.Y(n_161)
);

AO22x1_ASAP7_75t_L g204 ( 
.A1(n_161),
.A2(n_150),
.B1(n_134),
.B2(n_149),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_128),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_162),
.B(n_163),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_120),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_164),
.Y(n_202)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_168),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_121),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_169),
.B(n_176),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_107),
.B(n_98),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_170),
.A2(n_184),
.B(n_0),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_98),
.B(n_20),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_171),
.A2(n_138),
.B1(n_152),
.B2(n_155),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_172),
.B(n_6),
.Y(n_219)
);

AO22x2_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_136),
.B1(n_139),
.B2(n_141),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_180),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_174),
.A2(n_182),
.B1(n_177),
.B2(n_154),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_132),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_181),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_148),
.A2(n_117),
.B1(n_101),
.B2(n_108),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_188),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_16),
.B(n_0),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_0),
.C(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_186),
.Y(n_191)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_193),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_218),
.B1(n_170),
.B2(n_160),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_197),
.A2(n_212),
.B(n_161),
.Y(n_237)
);

NOR2x1_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_147),
.Y(n_200)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_140),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_208),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_209),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_151),
.Y(n_208)
);

OAI32xp33_ASAP7_75t_L g209 ( 
.A1(n_175),
.A2(n_117),
.A3(n_101),
.B1(n_4),
.B2(n_5),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_217),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_158),
.A2(n_178),
.B(n_188),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_8),
.B1(n_2),
.B2(n_5),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_214),
.A2(n_163),
.B1(n_177),
.B2(n_167),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_166),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_215),
.B(n_216),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_181),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_15),
.C(n_6),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_219),
.B(n_184),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_207),
.B(n_180),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_SL g261 ( 
.A(n_220),
.B(n_240),
.C(n_210),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_221),
.A2(n_222),
.B1(n_193),
.B2(n_204),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_192),
.A2(n_189),
.B1(n_173),
.B2(n_157),
.Y(n_223)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_237),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_194),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_231),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_189),
.B1(n_161),
.B2(n_187),
.Y(n_227)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_235),
.Y(n_255)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_191),
.B(n_179),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_236),
.B(n_239),
.Y(n_259)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_238),
.Y(n_254)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

NOR3xp33_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_173),
.C(n_190),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_203),
.B(n_182),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_226),
.Y(n_245)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_195),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_243),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_192),
.B(n_159),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_213),
.B1(n_218),
.B2(n_205),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_252),
.Y(n_272)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

OA22x2_ASAP7_75t_L g248 ( 
.A1(n_229),
.A2(n_204),
.B1(n_209),
.B2(n_196),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_248),
.A2(n_257),
.B(n_7),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_226),
.C(n_208),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_258),
.C(n_241),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_212),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_253),
.A2(n_228),
.B1(n_221),
.B2(n_233),
.Y(n_265)
);

XOR2x2_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_200),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_219),
.C(n_197),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_211),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_262),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_234),
.B(n_243),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_205),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_265),
.A2(n_276),
.B1(n_248),
.B2(n_262),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_266),
.B(n_278),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_228),
.C(n_241),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_260),
.C(n_250),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_259),
.B(n_258),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_270),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_257),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_231),
.Y(n_273)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_264),
.A2(n_195),
.B1(n_183),
.B2(n_168),
.Y(n_275)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_251),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_248),
.B(n_263),
.Y(n_284)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_279),
.B(n_280),
.Y(n_293)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_249),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_282),
.A2(n_284),
.B1(n_8),
.B2(n_11),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_286),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_266),
.C(n_269),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_269),
.C(n_272),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_294),
.Y(n_299)
);

INVxp33_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_275),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_265),
.B(n_246),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_287),
.C(n_285),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_289),
.A2(n_267),
.B(n_277),
.Y(n_296)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_296),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_290),
.B(n_246),
.Y(n_297)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_297),
.Y(n_313)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_292),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_300),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_252),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_291),
.B(n_13),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_272),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_303),
.Y(n_310)
);

NOR2x1_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_11),
.Y(n_305)
);

NOR2x1_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_284),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_SL g315 ( 
.A1(n_306),
.A2(n_305),
.B(n_299),
.C(n_302),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_311),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_281),
.C(n_288),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_312),
.A2(n_309),
.B(n_306),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_313),
.A2(n_298),
.B1(n_295),
.B2(n_304),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_314),
.A2(n_315),
.B(n_317),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_318)
);

NOR3xp33_ASAP7_75t_SL g320 ( 
.A(n_318),
.B(n_309),
.C(n_15),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_315),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_319),
.C(n_316),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_310),
.C(n_14),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_14),
.Y(n_324)
);


endmodule