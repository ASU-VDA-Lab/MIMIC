module fake_jpeg_28517_n_541 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_541);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_541;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_17),
.B(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_52),
.B(n_53),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_0),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_55),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_35),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_81),
.Y(n_107)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_1),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_73),
.B(n_92),
.Y(n_137)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_75),
.Y(n_148)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_41),
.A2(n_1),
.B(n_2),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_101),
.C(n_51),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_35),
.B(n_2),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_82),
.Y(n_165)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_36),
.B(n_2),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_95),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_87),
.Y(n_158)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_42),
.B(n_3),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_36),
.B(n_3),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_44),
.B(n_3),
.C(n_4),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

INVx4_ASAP7_75t_SL g103 ( 
.A(n_22),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_76),
.A2(n_39),
.B1(n_48),
.B2(n_47),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_104),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_112),
.A2(n_50),
.B(n_29),
.Y(n_206)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_65),
.A2(n_30),
.B1(n_46),
.B2(n_44),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_130),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_39),
.B1(n_48),
.B2(n_47),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_152),
.B1(n_166),
.B2(n_21),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_68),
.A2(n_46),
.B1(n_31),
.B2(n_22),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_56),
.A2(n_46),
.B1(n_51),
.B2(n_34),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_74),
.A2(n_40),
.B1(n_38),
.B2(n_37),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_96),
.A2(n_40),
.B1(n_38),
.B2(n_37),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_144),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_228)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_98),
.A2(n_23),
.B1(n_27),
.B2(n_34),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_57),
.B(n_23),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_164),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_60),
.B(n_27),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_61),
.A2(n_62),
.B1(n_89),
.B2(n_72),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_168),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_124),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_169),
.B(n_179),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_170),
.B(n_177),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_158),
.A2(n_64),
.B1(n_59),
.B2(n_99),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_172),
.A2(n_178),
.B1(n_186),
.B2(n_191),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_173),
.Y(n_247)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_175),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_79),
.B1(n_85),
.B2(n_80),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_176),
.A2(n_157),
.B1(n_156),
.B2(n_146),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_117),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_158),
.A2(n_99),
.B1(n_87),
.B2(n_22),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_113),
.B(n_51),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_181),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_114),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_106),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_184),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_185),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_124),
.A2(n_31),
.B1(n_34),
.B2(n_32),
.Y(n_186)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_187),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_135),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_189),
.B(n_192),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_190),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_105),
.A2(n_31),
.B1(n_32),
.B2(n_50),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_137),
.Y(n_192)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_128),
.A2(n_31),
.B1(n_32),
.B2(n_50),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_194),
.A2(n_207),
.B1(n_217),
.B2(n_223),
.Y(n_273)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_114),
.Y(n_197)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_197),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_198),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_109),
.B(n_29),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_199),
.B(n_210),
.Y(n_232)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_115),
.Y(n_200)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_200),
.Y(n_268)
);

NOR2xp67_ASAP7_75t_L g202 ( 
.A(n_137),
.B(n_31),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_202),
.B(n_8),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_113),
.B(n_33),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_203),
.B(n_211),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_120),
.Y(n_204)
);

CKINVDCx12_ASAP7_75t_R g240 ( 
.A(n_204),
.Y(n_240)
);

AND2x2_ASAP7_75t_SL g266 ( 
.A(n_206),
.B(n_9),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_122),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_208),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_107),
.B(n_29),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_129),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_151),
.B(n_161),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_212),
.B(n_216),
.Y(n_258)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_108),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_213),
.Y(n_260)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_214),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_148),
.B(n_21),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_126),
.Y(n_217)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_121),
.B(n_3),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_218),
.Y(n_265)
);

AO22x2_ASAP7_75t_L g219 ( 
.A1(n_130),
.A2(n_21),
.B1(n_33),
.B2(n_6),
.Y(n_219)
);

AO22x1_ASAP7_75t_SL g236 ( 
.A1(n_219),
.A2(n_150),
.B1(n_138),
.B2(n_142),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_116),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_220),
.B(n_221),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_162),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_131),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_222),
.B(n_224),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_126),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_150),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_134),
.B(n_4),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_225),
.B(n_226),
.Y(n_274)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_121),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_148),
.B(n_4),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_227),
.B(n_229),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_228),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_231)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_133),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_231),
.A2(n_224),
.B1(n_223),
.B2(n_217),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_236),
.A2(n_13),
.B(n_17),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_215),
.A2(n_127),
.B1(n_160),
.B2(n_157),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_237),
.B(n_249),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_241),
.A2(n_233),
.B1(n_236),
.B2(n_230),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_171),
.B(n_156),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_242),
.B(n_245),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_209),
.A2(n_146),
.B1(n_125),
.B2(n_119),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_243),
.A2(n_279),
.B1(n_186),
.B2(n_191),
.Y(n_281)
);

AO22x1_ASAP7_75t_SL g245 ( 
.A1(n_219),
.A2(n_125),
.B1(n_119),
.B2(n_118),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_118),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_246),
.B(n_251),
.Y(n_292)
);

NAND2xp33_ASAP7_75t_SL g249 ( 
.A(n_177),
.B(n_162),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_250),
.B(n_12),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_18),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_SL g253 ( 
.A1(n_215),
.A2(n_9),
.B(n_11),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_253),
.Y(n_320)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_170),
.A2(n_18),
.B1(n_11),
.B2(n_12),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_256),
.A2(n_197),
.B1(n_182),
.B2(n_15),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_184),
.B(n_195),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_259),
.B(n_270),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_266),
.B(n_180),
.C(n_213),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_200),
.B(n_9),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_174),
.B(n_196),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_275),
.B(n_242),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_219),
.B(n_11),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_276),
.B(n_219),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_222),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_281),
.A2(n_285),
.B1(n_286),
.B2(n_291),
.Y(n_342)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_282),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_283),
.A2(n_269),
.B(n_277),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_263),
.A2(n_206),
.B(n_172),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_284),
.A2(n_307),
.B(n_322),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_276),
.A2(n_194),
.B1(n_178),
.B2(n_229),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_244),
.Y(n_287)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_287),
.Y(n_349)
);

OAI21x1_ASAP7_75t_R g288 ( 
.A1(n_245),
.A2(n_181),
.B(n_187),
.Y(n_288)
);

INVx11_ASAP7_75t_L g350 ( 
.A(n_288),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_258),
.B(n_232),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_289),
.B(n_293),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_276),
.A2(n_205),
.B1(n_188),
.B2(n_207),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_258),
.B(n_201),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_294),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_295),
.B(n_302),
.Y(n_330)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_268),
.Y(n_296)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_296),
.Y(n_365)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_297),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_299),
.B(n_317),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_300),
.A2(n_234),
.B1(n_271),
.B2(n_248),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_280),
.A2(n_198),
.B1(n_185),
.B2(n_183),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_255),
.B(n_175),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_168),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_303),
.B(n_306),
.Y(n_331)
);

BUFx24_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_304),
.Y(n_355)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_305),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_252),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_238),
.A2(n_193),
.B1(n_208),
.B2(n_190),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_240),
.Y(n_308)
);

NAND2x1_ASAP7_75t_SL g346 ( 
.A(n_308),
.B(n_257),
.Y(n_346)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_309),
.B(n_310),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_232),
.B(n_261),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_247),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_315),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_238),
.A2(n_204),
.B1(n_190),
.B2(n_15),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_312),
.A2(n_314),
.B1(n_233),
.B2(n_257),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_252),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_313),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_243),
.A2(n_204),
.B1(n_14),
.B2(n_16),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_254),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_316),
.A2(n_273),
.B1(n_231),
.B2(n_237),
.Y(n_341)
);

INVx8_ASAP7_75t_L g318 ( 
.A(n_234),
.Y(n_318)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_318),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_266),
.B(n_238),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_246),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_321),
.A2(n_236),
.B1(n_245),
.B2(n_230),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_265),
.A2(n_236),
.B1(n_245),
.B2(n_266),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_254),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_323),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_234),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_324),
.Y(n_353)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_254),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_325),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_283),
.A2(n_265),
.B(n_250),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_327),
.A2(n_366),
.B(n_339),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_333),
.A2(n_343),
.B1(n_311),
.B2(n_309),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_336),
.B(n_344),
.Y(n_368)
);

AOI32xp33_ASAP7_75t_L g338 ( 
.A1(n_284),
.A2(n_262),
.A3(n_249),
.B1(n_278),
.B2(n_272),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_310),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_341),
.A2(n_351),
.B1(n_354),
.B2(n_357),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_289),
.B(n_251),
.C(n_260),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_SL g395 ( 
.A(n_346),
.B(n_304),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_270),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_347),
.B(n_299),
.Y(n_374)
);

AND2x2_ASAP7_75t_SL g386 ( 
.A(n_348),
.B(n_292),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_290),
.A2(n_280),
.B1(n_235),
.B2(n_248),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_290),
.A2(n_280),
.B1(n_235),
.B2(n_271),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_316),
.A2(n_326),
.B(n_320),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_359),
.A2(n_326),
.B(n_307),
.Y(n_367)
);

OAI32xp33_ASAP7_75t_L g361 ( 
.A1(n_317),
.A2(n_264),
.A3(n_260),
.B1(n_277),
.B2(n_252),
.Y(n_361)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_361),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_324),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_363),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_322),
.A2(n_288),
.B1(n_282),
.B2(n_305),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_364),
.A2(n_312),
.B1(n_286),
.B2(n_293),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_326),
.A2(n_264),
.B(n_267),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_367),
.A2(n_375),
.B(n_395),
.Y(n_422)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_349),
.Y(n_370)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_370),
.Y(n_420)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_349),
.Y(n_371)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_371),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_373),
.B(n_377),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_338),
.Y(n_406)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_352),
.Y(n_376)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_376),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_341),
.A2(n_285),
.B1(n_281),
.B2(n_288),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_298),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_379),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_362),
.B(n_298),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_344),
.B(n_308),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_380),
.B(n_383),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_342),
.A2(n_300),
.B1(n_291),
.B2(n_314),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_381),
.A2(n_384),
.B1(n_389),
.B2(n_393),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_382),
.A2(n_385),
.B1(n_398),
.B2(n_343),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_331),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_342),
.A2(n_292),
.B1(n_313),
.B2(n_306),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_364),
.A2(n_297),
.B1(n_296),
.B2(n_287),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_386),
.A2(n_400),
.B(n_359),
.Y(n_412)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_352),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_387),
.B(n_388),
.Y(n_416)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_365),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_350),
.A2(n_294),
.B1(n_325),
.B2(n_323),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_365),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_392),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_330),
.B(n_304),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_391),
.B(n_355),
.Y(n_413)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_358),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_358),
.B(n_315),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_394),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_334),
.B(n_304),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_396),
.B(n_334),
.C(n_348),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_351),
.A2(n_324),
.B1(n_318),
.B2(n_267),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_360),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_399),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_339),
.A2(n_366),
.B(n_327),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_406),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_402),
.B(n_372),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_396),
.B(n_347),
.C(n_336),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_404),
.B(n_407),
.C(n_417),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_374),
.B(n_335),
.C(n_345),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_384),
.A2(n_357),
.B1(n_350),
.B2(n_345),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_409),
.A2(n_411),
.B1(n_421),
.B2(n_372),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_381),
.A2(n_354),
.B1(n_358),
.B2(n_337),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_412),
.A2(n_414),
.B(n_425),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_413),
.B(n_415),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_373),
.A2(n_337),
.B(n_346),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_394),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_368),
.B(n_386),
.C(n_400),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_369),
.A2(n_361),
.B1(n_329),
.B2(n_356),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_377),
.A2(n_335),
.B1(n_329),
.B2(n_340),
.Y(n_423)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_423),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_367),
.A2(n_369),
.B(n_395),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_368),
.B(n_346),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_427),
.B(n_382),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_386),
.A2(n_340),
.B(n_355),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_428),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_378),
.B(n_379),
.C(n_385),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_430),
.B(n_390),
.C(n_387),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_389),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_431),
.B(n_397),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_416),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_434),
.B(n_435),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_430),
.B(n_391),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_436),
.A2(n_454),
.B1(n_402),
.B2(n_423),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_416),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_439),
.B(n_442),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_448),
.Y(n_468)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_420),
.Y(n_441)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_441),
.Y(n_465)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_420),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_443),
.A2(n_446),
.B1(n_409),
.B2(n_411),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_410),
.A2(n_392),
.B1(n_399),
.B2(n_397),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_424),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_449),
.Y(n_472)
);

MAJx2_ASAP7_75t_L g448 ( 
.A(n_401),
.B(n_370),
.C(n_371),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_424),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_406),
.B(n_393),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_450),
.B(n_451),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_452),
.Y(n_464)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_418),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_453),
.Y(n_466)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_418),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_404),
.B(n_388),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_455),
.B(n_456),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_410),
.B(n_376),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_417),
.B(n_328),
.C(n_398),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_457),
.B(n_407),
.C(n_427),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_460),
.A2(n_453),
.B1(n_454),
.B2(n_449),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_461),
.A2(n_469),
.B1(n_471),
.B2(n_447),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_462),
.B(n_437),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_455),
.B(n_428),
.C(n_419),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_467),
.B(n_470),
.C(n_473),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_436),
.A2(n_432),
.B1(n_434),
.B2(n_439),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_419),
.C(n_412),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_432),
.A2(n_419),
.B1(n_403),
.B2(n_421),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_444),
.B(n_448),
.C(n_451),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_433),
.A2(n_425),
.B(n_414),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_474),
.A2(n_433),
.B(n_438),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_422),
.C(n_426),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_479),
.C(n_445),
.Y(n_489)
);

FAx1_ASAP7_75t_SL g477 ( 
.A(n_450),
.B(n_408),
.CI(n_422),
.CON(n_477),
.SN(n_477)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_477),
.B(n_440),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_443),
.A2(n_403),
.B1(n_408),
.B2(n_405),
.Y(n_478)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_478),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_437),
.B(n_429),
.C(n_356),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_484),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_472),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_481),
.B(n_483),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_463),
.Y(n_483)
);

FAx1_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_456),
.CI(n_445),
.CON(n_484),
.SN(n_484)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_485),
.B(n_468),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_458),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_486),
.B(n_488),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_489),
.B(n_479),
.C(n_473),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_465),
.Y(n_490)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_490),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_464),
.B(n_441),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_491),
.A2(n_477),
.B(n_318),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_492),
.A2(n_496),
.B1(n_471),
.B2(n_461),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_493),
.A2(n_495),
.B1(n_239),
.B2(n_487),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_466),
.B(n_442),
.Y(n_494)
);

OAI321xp33_ASAP7_75t_L g500 ( 
.A1(n_494),
.A2(n_474),
.A3(n_332),
.B1(n_477),
.B2(n_353),
.C(n_360),
.Y(n_500)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_478),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_460),
.A2(n_332),
.B1(n_353),
.B2(n_363),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_498),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_487),
.A2(n_470),
.B1(n_476),
.B2(n_467),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_499),
.A2(n_485),
.B1(n_480),
.B2(n_496),
.Y(n_519)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_500),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_475),
.C(n_462),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_504),
.B(n_506),
.C(n_508),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_482),
.B(n_475),
.C(n_459),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_507),
.B(n_510),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_489),
.B(n_459),
.C(n_468),
.Y(n_508)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_509),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_499),
.A2(n_495),
.B1(n_493),
.B2(n_483),
.Y(n_513)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_513),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_504),
.B(n_488),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_514),
.B(n_520),
.Y(n_524)
);

AND2x2_ASAP7_75t_SL g515 ( 
.A(n_505),
.B(n_484),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_515),
.B(n_502),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_498),
.B(n_492),
.C(n_484),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_517),
.B(n_519),
.C(n_521),
.Y(n_526)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_501),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_516),
.A2(n_503),
.B(n_506),
.Y(n_523)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_523),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_518),
.A2(n_510),
.B1(n_494),
.B2(n_508),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_525),
.B(n_526),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_527),
.B(n_528),
.Y(n_530)
);

OAI211xp5_ASAP7_75t_L g528 ( 
.A1(n_515),
.A2(n_502),
.B(n_511),
.C(n_513),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_524),
.B(n_512),
.C(n_517),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_531),
.B(n_512),
.Y(n_534)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_530),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_533),
.A2(n_534),
.B(n_529),
.Y(n_535)
);

A2O1A1O1Ixp25_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_532),
.B(n_522),
.C(n_528),
.D(n_515),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_536),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_537),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_538),
.A2(n_527),
.B(n_521),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_507),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_497),
.B(n_239),
.Y(n_541)
);


endmodule