module real_jpeg_17872_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_620;
wire n_328;
wire n_456;
wire n_578;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_634;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_594;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_572;
wire n_405;
wire n_412;
wire n_586;
wire n_548;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_636;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_597;
wire n_42;
wire n_268;
wire n_313;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_1),
.A2(n_246),
.B1(n_250),
.B2(n_251),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_1),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_1),
.A2(n_250),
.B1(n_266),
.B2(n_269),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_1),
.A2(n_250),
.B1(n_323),
.B2(n_326),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_1),
.A2(n_84),
.B1(n_250),
.B2(n_259),
.Y(n_400)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_2),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_2),
.Y(n_134)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_2),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g353 ( 
.A(n_2),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_3),
.A2(n_136),
.B1(n_141),
.B2(n_145),
.Y(n_135)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_3),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_3),
.A2(n_145),
.B1(n_208),
.B2(n_212),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_3),
.A2(n_145),
.B1(n_385),
.B2(n_387),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_SL g595 ( 
.A1(n_3),
.A2(n_145),
.B1(n_360),
.B2(n_596),
.Y(n_595)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_4),
.Y(n_90)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_4),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_4),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_5),
.A2(n_116),
.B1(n_123),
.B2(n_124),
.Y(n_115)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_5),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_5),
.A2(n_123),
.B1(n_231),
.B2(n_236),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_5),
.A2(n_123),
.B1(n_366),
.B2(n_369),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g575 ( 
.A1(n_5),
.A2(n_123),
.B1(n_576),
.B2(n_577),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_6),
.A2(n_181),
.B1(n_190),
.B2(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_6),
.Y(n_193)
);

OAI22x1_ASAP7_75t_L g392 ( 
.A1(n_6),
.A2(n_193),
.B1(n_212),
.B2(n_343),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_6),
.A2(n_193),
.B1(n_601),
.B2(n_604),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_6),
.A2(n_193),
.B1(n_634),
.B2(n_636),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_7),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_7),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_7),
.Y(n_226)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_8),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_8),
.B(n_174),
.Y(n_331)
);

OAI32xp33_ASAP7_75t_L g419 ( 
.A1(n_8),
.A2(n_54),
.A3(n_300),
.B1(n_420),
.B2(n_423),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g453 ( 
.A1(n_8),
.A2(n_83),
.B1(n_454),
.B2(n_459),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_8),
.B(n_79),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_8),
.A2(n_108),
.B1(n_542),
.B2(n_544),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_9),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_9),
.A2(n_39),
.B1(n_259),
.B2(n_262),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_9),
.A2(n_39),
.B1(n_251),
.B2(n_415),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_9),
.A2(n_39),
.B1(n_504),
.B2(n_507),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_10),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_10),
.Y(n_122)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_10),
.Y(n_140)
);

BUFx4f_ASAP7_75t_L g329 ( 
.A(n_10),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_11),
.A2(n_148),
.B1(n_149),
.B2(n_151),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_11),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_11),
.A2(n_148),
.B1(n_312),
.B2(n_316),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_11),
.A2(n_148),
.B1(n_496),
.B2(n_499),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_11),
.A2(n_148),
.B1(n_539),
.B2(n_543),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_12),
.A2(n_149),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_12),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_12),
.A2(n_173),
.B1(n_281),
.B2(n_284),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_12),
.A2(n_173),
.B1(n_447),
.B2(n_449),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_SL g527 ( 
.A1(n_12),
.A2(n_173),
.B1(n_487),
.B2(n_528),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_21),
.B(n_23),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_14),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_14),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_14),
.A2(n_182),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_14),
.A2(n_92),
.B1(n_182),
.B2(n_582),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_SL g621 ( 
.A1(n_14),
.A2(n_182),
.B1(n_361),
.B2(n_622),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_16),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_16),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_16),
.Y(n_301)
);

BUFx5_ASAP7_75t_L g348 ( 
.A(n_16),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_16),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_17),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_17),
.A2(n_75),
.B1(n_295),
.B2(n_299),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_17),
.A2(n_75),
.B1(n_359),
.B2(n_361),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_17),
.A2(n_75),
.B1(n_429),
.B2(n_432),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx8_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_19),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_19),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_19),
.Y(n_292)
);

BUFx12f_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_644),
.B(n_647),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_566),
.B(n_637),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_404),
.B(n_561),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_335),
.C(n_375),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_272),
.B(n_303),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_29),
.B(n_272),
.C(n_563),
.Y(n_562)
);

XNOR2x1_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_175),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_30),
.B(n_176),
.C(n_241),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_80),
.C(n_146),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_32),
.B(n_146),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_45),
.B1(n_72),
.B2(n_78),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22x1_ASAP7_75t_L g279 ( 
.A1(n_34),
.A2(n_79),
.B1(n_280),
.B2(n_287),
.Y(n_279)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_37),
.Y(n_271)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_37),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_38),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_38),
.Y(n_320)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_43),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_45),
.A2(n_72),
.B1(n_78),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_45),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_45),
.A2(n_78),
.B1(n_265),
.B2(n_365),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_45),
.A2(n_78),
.B1(n_311),
.B2(n_453),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_45),
.A2(n_78),
.B1(n_384),
.B2(n_581),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_45),
.A2(n_78),
.B1(n_581),
.B2(n_600),
.Y(n_599)
);

AO21x1_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_54),
.B(n_61),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_52),
.Y(n_286)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_52),
.Y(n_584)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_53),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_53),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_53),
.Y(n_268)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_53),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_59),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_59),
.Y(n_605)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_60),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_62),
.Y(n_425)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_64),
.Y(n_220)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_64),
.Y(n_235)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_71),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_71),
.Y(n_494)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_79),
.A2(n_280),
.B1(n_287),
.B2(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_79),
.A2(n_287),
.B1(n_382),
.B2(n_383),
.Y(n_381)
);

OAI21xp33_ASAP7_75t_R g617 ( 
.A1(n_79),
.A2(n_287),
.B(n_618),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_80),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_107),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_81),
.B(n_107),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_87),
.B1(n_96),
.B2(n_99),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_SL g289 ( 
.A1(n_82),
.A2(n_83),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_83),
.B(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_83),
.B(n_227),
.Y(n_480)
);

OAI21xp33_ASAP7_75t_SL g491 ( 
.A1(n_83),
.A2(n_480),
.B(n_492),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_83),
.B(n_253),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_83),
.B(n_197),
.Y(n_549)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g262 ( 
.A(n_86),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx8_ASAP7_75t_L g603 ( 
.A(n_95),
.Y(n_603)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OA21x2_ASAP7_75t_L g157 ( 
.A1(n_100),
.A2(n_158),
.B(n_163),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_101),
.Y(n_360)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_102),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_102),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_105),
.A2(n_164),
.B1(n_166),
.B2(n_168),
.Y(n_163)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_114),
.B1(n_128),
.B2(n_135),
.Y(n_107)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_108),
.A2(n_135),
.B1(n_180),
.B2(n_253),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_108),
.A2(n_189),
.B(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_108),
.A2(n_503),
.B1(n_512),
.B2(n_517),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_108),
.A2(n_527),
.B1(n_542),
.B2(n_548),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

INVx6_ASAP7_75t_L g548 ( 
.A(n_109),
.Y(n_548)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_113),
.Y(n_202)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_113),
.Y(n_431)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_113),
.Y(n_488)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_113),
.Y(n_511)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_115),
.A2(n_178),
.B1(n_322),
.B2(n_330),
.Y(n_321)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_127),
.Y(n_506)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_133),
.Y(n_254)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_134),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_138),
.Y(n_325)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_139),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_144),
.Y(n_434)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_144),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_157),
.B1(n_169),
.B2(n_174),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_147),
.A2(n_157),
.B1(n_174),
.B2(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_SL g257 ( 
.A(n_157),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_157),
.A2(n_594),
.B1(n_595),
.B2(n_597),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_SL g645 ( 
.A1(n_157),
.A2(n_597),
.B(n_646),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_162),
.Y(n_261)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_166),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_170),
.A2(n_257),
.B1(n_258),
.B2(n_263),
.Y(n_256)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_174),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_241),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_194),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_177),
.A2(n_195),
.B(n_216),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_185),
.B2(n_188),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_178),
.A2(n_322),
.B1(n_428),
.B2(n_435),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_178),
.A2(n_526),
.B1(n_530),
.B2(n_533),
.Y(n_525)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_187),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_216),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_206),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_196),
.A2(n_217),
.B1(n_294),
.B2(n_302),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_196),
.A2(n_217),
.B1(n_391),
.B2(n_392),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_196),
.A2(n_217),
.B1(n_414),
.B2(n_446),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_196),
.A2(n_217),
.B1(n_491),
.B2(n_495),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_196),
.A2(n_217),
.B1(n_446),
.B2(n_495),
.Y(n_521)
);

OA21x2_ASAP7_75t_L g585 ( 
.A1(n_196),
.A2(n_217),
.B(n_392),
.Y(n_585)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_197),
.A2(n_230),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_197),
.A2(n_207),
.B1(n_244),
.B2(n_342),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_197),
.A2(n_244),
.B1(n_413),
.B2(n_416),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g217 ( 
.A(n_198),
.B(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_200),
.Y(n_483)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_229),
.Y(n_216)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_221),
.B1(n_224),
.B2(n_227),
.Y(n_218)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_225),
.Y(n_479)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_232),
.Y(n_343)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_234),
.Y(n_470)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_235),
.Y(n_240)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_255),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_242),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_252),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_245),
.Y(n_302)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_248),
.Y(n_500)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g435 ( 
.A(n_253),
.Y(n_435)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_264),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_256),
.B(n_264),
.C(n_338),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_257),
.A2(n_258),
.B1(n_263),
.B2(n_358),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_257),
.A2(n_263),
.B1(n_358),
.B2(n_400),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_257),
.A2(n_263),
.B1(n_400),
.B2(n_575),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g619 ( 
.A1(n_257),
.A2(n_263),
.B1(n_620),
.B2(n_621),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_SL g632 ( 
.A1(n_257),
.A2(n_263),
.B1(n_621),
.B2(n_633),
.Y(n_632)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_262),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_263),
.Y(n_597)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_276),
.C(n_277),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_273),
.A2(n_274),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_276),
.B(n_278),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_288),
.C(n_293),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_293),
.Y(n_306)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx2_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_306),
.Y(n_305)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_290),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_292),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_294),
.Y(n_416)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_295),
.Y(n_415)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_298),
.Y(n_450)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_301),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_332),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_304),
.B(n_332),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.C(n_308),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_305),
.B(n_407),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_307),
.B(n_308),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_321),
.C(n_331),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_309),
.B(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_315),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_315),
.Y(n_422)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_320),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_321),
.B(n_331),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

A2O1A1O1Ixp25_ASAP7_75t_L g561 ( 
.A1(n_335),
.A2(n_375),
.B(n_562),
.C(n_564),
.D(n_565),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_374),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_336),
.B(n_374),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_339),
.Y(n_336)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_337),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_355),
.B1(n_372),
.B2(n_373),
.Y(n_339)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_340),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_340),
.B(n_373),
.C(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_349),
.B1(n_350),
.B2(n_354),
.Y(n_340)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_341),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_341),
.B(n_350),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_349),
.A2(n_350),
.B1(n_398),
.B2(n_399),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g588 ( 
.A1(n_349),
.A2(n_399),
.B(n_401),
.Y(n_588)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_355),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_371),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_364),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_371),
.C(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_363),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_364),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_365),
.Y(n_382)
);

INVx8_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_402),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_376),
.B(n_402),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_379),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_377),
.B(n_609),
.C(n_610),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_394),
.Y(n_379)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_380),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_381),
.A2(n_390),
.B(n_393),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_381),
.B(n_390),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_386),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_393),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_393),
.A2(n_572),
.B1(n_587),
.B2(n_613),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_394),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_395),
.A2(n_396),
.B1(n_397),
.B2(n_401),
.Y(n_394)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_395),
.Y(n_401)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

AOI21x1_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_436),
.B(n_560),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_408),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_406),
.B(n_408),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_412),
.C(n_417),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_409),
.A2(n_410),
.B1(n_439),
.B2(n_440),
.Y(n_438)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_412),
.A2(n_417),
.B1(n_418),
.B2(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_412),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_426),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_419),
.A2(n_426),
.B1(n_427),
.B2(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_419),
.Y(n_444)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_428),
.Y(n_517)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_464),
.B(n_559),
.Y(n_436)
);

NOR2x1_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_442),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_438),
.B(n_442),
.Y(n_559)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_445),
.C(n_451),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_443),
.B(n_556),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_445),
.A2(n_451),
.B1(n_452),
.B2(n_557),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_445),
.Y(n_557)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx6_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_465),
.A2(n_553),
.B(n_558),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_466),
.A2(n_523),
.B(n_552),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_501),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_467),
.B(n_501),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_489),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_468),
.A2(n_489),
.B1(n_490),
.B2(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_468),
.Y(n_535)
);

OAI32xp33_ASAP7_75t_L g468 ( 
.A1(n_469),
.A2(n_471),
.A3(n_476),
.B1(n_480),
.B2(n_481),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_484),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_518),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_502),
.B(n_520),
.C(n_522),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_503),
.Y(n_533)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_507),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_516),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_519),
.A2(n_520),
.B1(n_521),
.B2(n_522),
.Y(n_518)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_519),
.Y(n_522)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_524),
.A2(n_536),
.B(n_551),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_534),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_525),
.B(n_534),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_528),
.Y(n_543)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx4_ASAP7_75t_SL g531 ( 
.A(n_532),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_532),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_537),
.A2(n_546),
.B(n_550),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_541),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_540),
.Y(n_538)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_549),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_547),
.B(n_549),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_555),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_554),
.B(n_555),
.Y(n_558)
);

NOR3xp33_ASAP7_75t_L g566 ( 
.A(n_567),
.B(n_614),
.C(n_630),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_568),
.B(n_607),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_569),
.A2(n_640),
.B(n_641),
.Y(n_639)
);

NOR2xp67_ASAP7_75t_L g569 ( 
.A(n_570),
.B(n_589),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_570),
.B(n_589),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_571),
.B(n_587),
.C(n_588),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_572),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_573),
.A2(n_574),
.B1(n_579),
.B2(n_586),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_573),
.B(n_580),
.C(n_585),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_573),
.A2(n_574),
.B1(n_592),
.B2(n_606),
.Y(n_591)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_574),
.B(n_592),
.C(n_629),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_575),
.Y(n_594)
);

INVx3_ASAP7_75t_SL g577 ( 
.A(n_578),
.Y(n_577)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_578),
.Y(n_635)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_579),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_580),
.B(n_585),
.Y(n_579)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

XNOR2x1_ASAP7_75t_L g598 ( 
.A(n_585),
.B(n_599),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_585),
.B(n_593),
.C(n_627),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_588),
.B(n_612),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_590),
.B(n_591),
.Y(n_589)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_590),
.Y(n_629)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_592),
.Y(n_606)
);

XNOR2x1_ASAP7_75t_L g592 ( 
.A(n_593),
.B(n_598),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_595),
.Y(n_620)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_599),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_600),
.Y(n_618)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_608),
.B(n_611),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_608),
.B(n_611),
.Y(n_640)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_615),
.Y(n_614)
);

A2O1A1O1Ixp25_ASAP7_75t_L g638 ( 
.A1(n_615),
.A2(n_631),
.B(n_639),
.C(n_642),
.D(n_643),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_616),
.B(n_628),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_616),
.B(n_632),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_616),
.B(n_628),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_616),
.B(n_632),
.Y(n_643)
);

FAx1_ASAP7_75t_SL g616 ( 
.A(n_617),
.B(n_619),
.CI(n_626),
.CON(n_616),
.SN(n_616)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_623),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_624),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_632),
.B(n_645),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_632),
.B(n_645),
.Y(n_648)
);

CKINVDCx16_ASAP7_75t_R g646 ( 
.A(n_633),
.Y(n_646)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_635),
.Y(n_634)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_638),
.Y(n_637)
);

CKINVDCx16_ASAP7_75t_R g647 ( 
.A(n_648),
.Y(n_647)
);


endmodule