module fake_jpeg_28310_n_19 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_19);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_19;

wire n_13;
wire n_10;
wire n_14;
wire n_18;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_8),
.B(n_0),
.Y(n_10)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_10),
.A2(n_11),
.B(n_0),
.Y(n_13)
);

O2A1O1Ixp33_ASAP7_75t_L g11 ( 
.A1(n_8),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_11)
);

NAND3xp33_ASAP7_75t_L g12 ( 
.A(n_11),
.B(n_5),
.C(n_6),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_13),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_15),
.C(n_9),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_17),
.B(n_15),
.C(n_9),
.Y(n_18)
);

AOI322xp5_ASAP7_75t_L g19 ( 
.A1(n_18),
.A2(n_7),
.A3(n_2),
.B1(n_3),
.B2(n_6),
.C1(n_1),
.C2(n_0),
.Y(n_19)
);


endmodule