module fake_jpeg_22524_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_7),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_23),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_0),
.Y(n_53)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVxp67_ASAP7_75t_SL g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_43),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_32),
.B1(n_17),
.B2(n_28),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_24),
.B1(n_23),
.B2(n_21),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_32),
.B1(n_17),
.B2(n_26),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_26),
.B1(n_22),
.B2(n_24),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_32),
.B1(n_17),
.B2(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_56),
.B1(n_28),
.B2(n_27),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_49),
.B(n_53),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_51),
.Y(n_81)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_28),
.B1(n_31),
.B2(n_26),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_37),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_57),
.Y(n_64)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_58),
.B(n_62),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_68),
.Y(n_89)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_65),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_31),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_73),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_76),
.B1(n_80),
.B2(n_85),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_48),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_41),
.C(n_27),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_86),
.C(n_49),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_72),
.B(n_83),
.Y(n_110)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_75),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_77),
.A2(n_44),
.B1(n_52),
.B2(n_55),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_48),
.B(n_9),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_61),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_19),
.B1(n_18),
.B2(n_16),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_0),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_88),
.Y(n_121)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_94),
.Y(n_131)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_95),
.B(n_96),
.Y(n_117)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_97),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_70),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_62),
.C(n_59),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_100),
.C(n_98),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_61),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

OAI22x1_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_97),
.B1(n_105),
.B2(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_81),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_108),
.B(n_69),
.Y(n_112)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_106),
.B(n_109),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_76),
.B1(n_81),
.B2(n_70),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_81),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_86),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_112),
.A2(n_130),
.B(n_25),
.Y(n_162)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_113),
.B(n_120),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_63),
.C(n_66),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_118),
.C(n_135),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_126),
.B1(n_129),
.B2(n_84),
.Y(n_139)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_124),
.Y(n_141)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_133),
.B1(n_137),
.B2(n_103),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_91),
.A2(n_67),
.B1(n_64),
.B2(n_85),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_133),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_101),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_128),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_91),
.A2(n_64),
.B1(n_44),
.B2(n_60),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_92),
.A2(n_108),
.B(n_104),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_90),
.A2(n_44),
.B1(n_66),
.B2(n_60),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_68),
.B1(n_86),
.B2(n_52),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_90),
.C(n_93),
.Y(n_135)
);

XOR2x2_ASAP7_75t_SL g136 ( 
.A(n_100),
.B(n_68),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_SL g156 ( 
.A(n_136),
.B(n_25),
.C(n_18),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_60),
.B1(n_69),
.B2(n_58),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_86),
.Y(n_138)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_162),
.B1(n_120),
.B2(n_129),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_SL g171 ( 
.A1(n_140),
.A2(n_144),
.B(n_150),
.Y(n_171)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_143),
.B(n_156),
.Y(n_166)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_102),
.B(n_43),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_123),
.A2(n_134),
.B1(n_126),
.B2(n_118),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_152),
.B1(n_42),
.B2(n_16),
.Y(n_176)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_151),
.Y(n_170)
);

HB1xp67_ASAP7_75t_SL g150 ( 
.A(n_112),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_74),
.C(n_101),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_115),
.A2(n_94),
.B1(n_87),
.B2(n_42),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_42),
.Y(n_153)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_157),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_25),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_158),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_114),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_159),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_25),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_16),
.B(n_1),
.C(n_3),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_132),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_161),
.Y(n_177)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_119),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_19),
.Y(n_164)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_167),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_154),
.A2(n_124),
.B1(n_119),
.B2(n_114),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_169),
.A2(n_181),
.B(n_15),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_149),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_175),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_139),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_147),
.B1(n_152),
.B2(n_157),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_179),
.A2(n_186),
.B1(n_181),
.B2(n_173),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_146),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_182),
.Y(n_211)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_142),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_165),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_188),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_160),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_144),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_138),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_191),
.B(n_201),
.Y(n_218)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_197),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_145),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_162),
.B1(n_144),
.B2(n_164),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_143),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_145),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_153),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_203),
.A2(n_207),
.B1(n_209),
.B2(n_212),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_151),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_178),
.C(n_187),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_205),
.A2(n_208),
.B1(n_190),
.B2(n_183),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_1),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_206),
.Y(n_216)
);

AO21x1_ASAP7_75t_L g209 ( 
.A1(n_172),
.A2(n_4),
.B(n_5),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_176),
.B(n_4),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_210),
.B(n_186),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_220),
.Y(n_238)
);

FAx1_ASAP7_75t_SL g214 ( 
.A(n_198),
.B(n_172),
.CI(n_199),
.CON(n_214),
.SN(n_214)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_214),
.B(n_207),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_219),
.C(n_226),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_178),
.C(n_187),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_225),
.A2(n_210),
.B1(n_209),
.B2(n_10),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_180),
.C(n_184),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_180),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_228),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_184),
.Y(n_228)
);

INVx13_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_232),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_241),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_233),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_194),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_222),
.A2(n_198),
.B1(n_212),
.B2(n_208),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_237),
.A2(n_242),
.B1(n_213),
.B2(n_218),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_211),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_239),
.B(n_215),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_226),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_177),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_221),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_242)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_248),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_229),
.C(n_219),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_251),
.Y(n_260)
);

NAND4xp25_ASAP7_75t_SL g249 ( 
.A(n_231),
.B(n_8),
.C(n_9),
.D(n_11),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_249),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_236),
.B(n_237),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_229),
.C(n_12),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_238),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_262),
.C(n_246),
.Y(n_263)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_238),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_255),
.B(n_244),
.Y(n_267)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_257),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_15),
.B1(n_242),
.B2(n_252),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_261),
.B(n_243),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_15),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_267),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_244),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_265),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_262),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_271),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_263),
.A2(n_256),
.B(n_253),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_274),
.A2(n_270),
.B(n_269),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_275),
.Y(n_276)
);

A2O1A1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_273),
.B(n_266),
.C(n_264),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_249),
.B(n_260),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_254),
.Y(n_279)
);


endmodule