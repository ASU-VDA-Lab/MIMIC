module real_aes_6586_n_207 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_174, n_156, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_183, n_205, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_3, n_41, n_140, n_153, n_75, n_178, n_19, n_71, n_180, n_40, n_49, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_81, n_133, n_48, n_204, n_37, n_117, n_97, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_207);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_97;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_207;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_216;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_649;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_397;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_686;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_208;
wire n_215;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_0), .A2(n_52), .B1(n_255), .B2(n_423), .Y(n_535) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_1), .A2(n_76), .B1(n_244), .B2(n_354), .Y(n_534) );
AOI22xp33_ASAP7_75t_SL g660 ( .A1(n_2), .A2(n_19), .B1(n_354), .B2(n_582), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_3), .A2(n_90), .B1(n_378), .B2(n_379), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_4), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_5), .A2(n_157), .B1(n_457), .B2(n_460), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_6), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_7), .A2(n_21), .B1(n_492), .B2(n_493), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_8), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g414 ( .A(n_9), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_10), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_11), .A2(n_95), .B1(n_395), .B2(n_481), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_12), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_13), .A2(n_155), .B1(n_335), .B2(n_418), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_14), .A2(n_34), .B1(n_225), .B2(n_242), .Y(n_224) );
AO22x2_ASAP7_75t_L g239 ( .A1(n_15), .A2(n_65), .B1(n_231), .B2(n_236), .Y(n_239) );
INVx1_ASAP7_75t_L g678 ( .A(n_15), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_16), .A2(n_55), .B1(n_225), .B2(n_347), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_17), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_18), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_20), .A2(n_195), .B1(n_354), .B2(n_376), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_22), .A2(n_114), .B1(n_369), .B2(n_455), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_23), .A2(n_141), .B1(n_255), .B2(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_24), .A2(n_32), .B1(n_264), .B2(n_459), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_25), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_26), .A2(n_100), .B1(n_250), .B2(n_373), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_27), .Y(n_573) );
AOI22xp33_ASAP7_75t_SL g655 ( .A1(n_28), .A2(n_142), .B1(n_568), .B2(n_656), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_29), .A2(n_172), .B1(n_455), .B2(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_30), .A2(n_121), .B1(n_252), .B2(n_539), .Y(n_538) );
AO22x2_ASAP7_75t_L g241 ( .A1(n_31), .A2(n_68), .B1(n_231), .B2(n_232), .Y(n_241) );
INVx1_ASAP7_75t_L g679 ( .A(n_31), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g658 ( .A1(n_33), .A2(n_75), .B1(n_378), .B2(n_572), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_35), .A2(n_180), .B1(n_571), .B2(n_572), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_36), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_37), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_38), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_39), .A2(n_154), .B1(n_357), .B2(n_373), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_40), .A2(n_177), .B1(n_581), .B2(n_582), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_41), .A2(n_69), .B1(n_273), .B2(n_276), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_42), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_43), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_44), .A2(n_83), .B1(n_226), .B2(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_45), .A2(n_115), .B1(n_692), .B2(n_693), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_46), .A2(n_169), .B1(n_443), .B2(n_621), .Y(n_620) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_47), .A2(n_171), .B1(n_587), .B2(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_48), .A2(n_130), .B1(n_298), .B2(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_49), .A2(n_60), .B1(n_442), .B2(n_443), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_50), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_51), .A2(n_99), .B1(n_394), .B2(n_395), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_53), .B(n_603), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_54), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_56), .A2(n_72), .B1(n_587), .B2(n_588), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_57), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_58), .A2(n_62), .B1(n_347), .B2(n_418), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_59), .A2(n_110), .B1(n_261), .B2(n_266), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_61), .A2(n_111), .B1(n_385), .B2(n_387), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_63), .A2(n_113), .B1(n_252), .B2(n_254), .Y(n_349) );
AOI222xp33_ASAP7_75t_L g699 ( .A1(n_64), .A2(n_67), .B1(n_92), .B2(n_294), .C1(n_387), .C2(n_700), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_66), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_70), .Y(n_549) );
AOI22xp33_ASAP7_75t_SL g653 ( .A1(n_71), .A2(n_192), .B1(n_298), .B2(n_411), .Y(n_653) );
INVx1_ASAP7_75t_L g215 ( .A(n_73), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_74), .A2(n_188), .B1(n_356), .B2(n_568), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_77), .A2(n_205), .B1(n_250), .B2(n_539), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_78), .Y(n_663) );
INVx1_ASAP7_75t_L g213 ( .A(n_79), .Y(n_213) );
AOI211xp5_ASAP7_75t_L g207 ( .A1(n_80), .A2(n_208), .B(n_217), .C(n_680), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_81), .A2(n_97), .B1(n_307), .B2(n_411), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_82), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_84), .A2(n_173), .B1(n_369), .B2(n_371), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g594 ( .A(n_85), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_86), .B(n_306), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_87), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_88), .B(n_626), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_89), .Y(n_601) );
OA22x2_ASAP7_75t_L g400 ( .A1(n_91), .A2(n_401), .B1(n_402), .B2(n_426), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_91), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g296 ( .A(n_93), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_94), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_96), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_98), .A2(n_102), .B1(n_528), .B2(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_101), .A2(n_118), .B1(n_268), .B2(n_582), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_103), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_104), .B(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_105), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_106), .B(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g216 ( .A(n_107), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_108), .A2(n_128), .B1(n_358), .B2(n_591), .Y(n_590) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_109), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_112), .Y(n_314) );
AND2x6_ASAP7_75t_L g212 ( .A(n_116), .B(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_116), .Y(n_672) );
AO22x2_ASAP7_75t_L g230 ( .A1(n_117), .A2(n_166), .B1(n_231), .B2(n_232), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_119), .A2(n_140), .B1(n_347), .B2(n_463), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_120), .A2(n_146), .B1(n_352), .B2(n_353), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_122), .B(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_123), .A2(n_186), .B1(n_357), .B2(n_423), .Y(n_422) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_124), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_125), .A2(n_682), .B1(n_683), .B2(n_702), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_125), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_126), .A2(n_153), .B1(n_376), .B2(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g467 ( .A(n_127), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_129), .A2(n_176), .B1(n_356), .B2(n_358), .Y(n_355) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_131), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_132), .A2(n_139), .B1(n_338), .B2(n_385), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_133), .B(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_134), .A2(n_150), .B1(n_264), .B2(n_490), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_135), .A2(n_136), .B1(n_268), .B2(n_631), .Y(n_630) );
AO22x2_ASAP7_75t_L g235 ( .A1(n_137), .A2(n_178), .B1(n_231), .B2(n_236), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_138), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_143), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_144), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_145), .A2(n_152), .B1(n_591), .B2(n_686), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_147), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g661 ( .A1(n_148), .A2(n_175), .B1(n_454), .B2(n_662), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_149), .A2(n_165), .B1(n_395), .B2(n_481), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_151), .A2(n_577), .B1(n_608), .B2(n_609), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_151), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_156), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_158), .A2(n_185), .B1(n_454), .B2(n_455), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_159), .B(n_624), .Y(n_623) );
AOI22xp33_ASAP7_75t_SL g646 ( .A1(n_160), .A2(n_189), .B1(n_443), .B2(n_481), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_161), .B(n_651), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_162), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_163), .B(n_305), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_164), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_166), .B(n_677), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_167), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_168), .Y(n_605) );
INVx1_ASAP7_75t_L g365 ( .A(n_170), .Y(n_365) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_174), .Y(n_638) );
INVx1_ASAP7_75t_L g675 ( .A(n_178), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_179), .A2(n_196), .B1(n_376), .B2(n_418), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_181), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_182), .A2(n_187), .B1(n_378), .B2(n_425), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g282 ( .A(n_183), .Y(n_282) );
INVxp67_ASAP7_75t_L g712 ( .A(n_184), .Y(n_712) );
XNOR2x2_ASAP7_75t_L g713 ( .A(n_184), .B(n_683), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_190), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_191), .A2(n_221), .B1(n_320), .B2(n_321), .Y(n_220) );
INVx1_ASAP7_75t_L g320 ( .A(n_191), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_193), .Y(n_336) );
INVx1_ASAP7_75t_L g231 ( .A(n_194), .Y(n_231) );
INVx1_ASAP7_75t_L g233 ( .A(n_194), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_197), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_198), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_199), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_200), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g303 ( .A(n_201), .Y(n_303) );
OA22x2_ASAP7_75t_L g470 ( .A1(n_202), .A2(n_471), .B1(n_472), .B2(n_473), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_202), .Y(n_471) );
AOI22x1_ASAP7_75t_L g324 ( .A1(n_203), .A2(n_325), .B1(n_359), .B2(n_360), .Y(n_324) );
INVx1_ASAP7_75t_L g359 ( .A(n_203), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_204), .A2(n_206), .B1(n_250), .B2(n_254), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_209), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_210), .Y(n_209) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_212), .B(n_214), .Y(n_211) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_213), .Y(n_671) );
OAI21xp5_ASAP7_75t_L g710 ( .A1(n_214), .A2(n_670), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
AOI221xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_511), .B1(n_665), .B2(n_666), .C(n_667), .Y(n_217) );
INVx1_ASAP7_75t_L g665 ( .A(n_218), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_362), .B1(n_509), .B2(n_510), .Y(n_218) );
INVx1_ASAP7_75t_L g509 ( .A(n_219), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_322), .B1(n_323), .B2(n_361), .Y(n_219) );
INVx1_ASAP7_75t_L g361 ( .A(n_220), .Y(n_361) );
INVx2_ASAP7_75t_L g321 ( .A(n_221), .Y(n_321) );
AND2x2_ASAP7_75t_SL g221 ( .A(n_222), .B(n_280), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_259), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_249), .Y(n_223) );
BUFx3_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
BUFx3_ASAP7_75t_L g581 ( .A(n_226), .Y(n_581) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g370 ( .A(n_227), .Y(n_370) );
BUFx2_ASAP7_75t_SL g454 ( .A(n_227), .Y(n_454) );
BUFx2_ASAP7_75t_SL g698 ( .A(n_227), .Y(n_698) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_237), .Y(n_227) );
AND2x6_ASAP7_75t_L g246 ( .A(n_228), .B(n_247), .Y(n_246) );
AND2x4_ASAP7_75t_L g264 ( .A(n_228), .B(n_265), .Y(n_264) );
AND2x6_ASAP7_75t_L g294 ( .A(n_228), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_234), .Y(n_228) );
AND2x2_ASAP7_75t_L g253 ( .A(n_229), .B(n_235), .Y(n_253) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_230), .B(n_235), .Y(n_258) );
AND2x2_ASAP7_75t_L g270 ( .A(n_230), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g302 ( .A(n_230), .B(n_239), .Y(n_302) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g236 ( .A(n_233), .Y(n_236) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g271 ( .A(n_235), .Y(n_271) );
INVx1_ASAP7_75t_L g301 ( .A(n_235), .Y(n_301) );
AND2x4_ASAP7_75t_L g252 ( .A(n_237), .B(n_253), .Y(n_252) );
AND2x4_ASAP7_75t_L g256 ( .A(n_237), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g269 ( .A(n_237), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_237), .B(n_270), .Y(n_506) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_240), .Y(n_237) );
OR2x2_ASAP7_75t_L g248 ( .A(n_238), .B(n_241), .Y(n_248) );
AND2x2_ASAP7_75t_L g265 ( .A(n_238), .B(n_241), .Y(n_265) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g295 ( .A(n_239), .B(n_241), .Y(n_295) );
AND2x2_ASAP7_75t_L g300 ( .A(n_240), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g313 ( .A(n_240), .Y(n_313) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g279 ( .A(n_241), .Y(n_279) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx5_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g501 ( .A(n_245), .Y(n_501) );
INVx4_ASAP7_75t_L g631 ( .A(n_245), .Y(n_631) );
INVx11_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx11_ASAP7_75t_L g348 ( .A(n_246), .Y(n_348) );
AND2x4_ASAP7_75t_L g526 ( .A(n_247), .B(n_253), .Y(n_526) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g284 ( .A(n_248), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
BUFx3_ASAP7_75t_L g378 ( .A(n_252), .Y(n_378) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_252), .Y(n_465) );
BUFx3_ASAP7_75t_L g492 ( .A(n_252), .Y(n_492) );
BUFx3_ASAP7_75t_L g571 ( .A(n_252), .Y(n_571) );
INVx1_ASAP7_75t_L g285 ( .A(n_253), .Y(n_285) );
NAND2x1p5_ASAP7_75t_L g289 ( .A(n_253), .B(n_265), .Y(n_289) );
AND2x6_ASAP7_75t_L g529 ( .A(n_253), .B(n_265), .Y(n_529) );
BUFx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
BUFx2_ASAP7_75t_L g379 ( .A(n_256), .Y(n_379) );
BUFx3_ASAP7_75t_L g425 ( .A(n_256), .Y(n_425) );
BUFx2_ASAP7_75t_SL g455 ( .A(n_256), .Y(n_455) );
BUFx3_ASAP7_75t_L g633 ( .A(n_256), .Y(n_633) );
BUFx2_ASAP7_75t_SL g662 ( .A(n_256), .Y(n_662) );
AND2x2_ASAP7_75t_L g373 ( .A(n_257), .B(n_313), .Y(n_373) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x6_ASAP7_75t_L g278 ( .A(n_258), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_272), .Y(n_259) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
BUFx3_ASAP7_75t_L g352 ( .A(n_264), .Y(n_352) );
BUFx3_ASAP7_75t_L g376 ( .A(n_264), .Y(n_376) );
INVx6_ASAP7_75t_L g569 ( .A(n_264), .Y(n_569) );
AND2x2_ASAP7_75t_L g275 ( .A(n_265), .B(n_270), .Y(n_275) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx3_ASAP7_75t_L g354 ( .A(n_269), .Y(n_354) );
BUFx3_ASAP7_75t_L g418 ( .A(n_269), .Y(n_418) );
INVx1_ASAP7_75t_L g319 ( .A(n_271), .Y(n_319) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx5_ASAP7_75t_L g357 ( .A(n_274), .Y(n_357) );
INVx4_ASAP7_75t_L g459 ( .A(n_274), .Y(n_459) );
INVx1_ASAP7_75t_L g490 ( .A(n_274), .Y(n_490) );
INVx3_ASAP7_75t_L g636 ( .A(n_274), .Y(n_636) );
BUFx3_ASAP7_75t_L g657 ( .A(n_274), .Y(n_657) );
INVx8_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
BUFx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
BUFx4f_ASAP7_75t_SL g358 ( .A(n_277), .Y(n_358) );
BUFx2_ASAP7_75t_L g493 ( .A(n_277), .Y(n_493) );
BUFx2_ASAP7_75t_L g572 ( .A(n_277), .Y(n_572) );
INVx6_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_278), .A2(n_316), .B1(n_413), .B2(n_414), .Y(n_412) );
INVx1_ASAP7_75t_L g460 ( .A(n_278), .Y(n_460) );
INVx1_ASAP7_75t_SL g539 ( .A(n_278), .Y(n_539) );
INVx1_ASAP7_75t_L g386 ( .A(n_279), .Y(n_386) );
NOR3xp33_ASAP7_75t_L g280 ( .A(n_281), .B(n_290), .C(n_309), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B1(n_286), .B2(n_287), .Y(n_281) );
INVx1_ASAP7_75t_L g556 ( .A(n_283), .Y(n_556) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g330 ( .A(n_284), .Y(n_330) );
OAI221xp5_ASAP7_75t_L g380 ( .A1(n_284), .A2(n_381), .B1(n_382), .B2(n_383), .C(n_384), .Y(n_380) );
BUFx3_ASAP7_75t_L g406 ( .A(n_284), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_287), .A2(n_405), .B1(n_406), .B2(n_407), .Y(n_404) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g332 ( .A(n_288), .Y(n_332) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx3_ASAP7_75t_L g382 ( .A(n_289), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_296), .B1(n_297), .B2(n_303), .C(n_304), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx4_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
BUFx2_ASAP7_75t_L g440 ( .A(n_293), .Y(n_440) );
INVx4_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_294), .Y(n_335) );
BUFx3_ASAP7_75t_L g391 ( .A(n_294), .Y(n_391) );
INVx2_ASAP7_75t_L g519 ( .A(n_294), .Y(n_519) );
INVx2_ASAP7_75t_L g598 ( .A(n_294), .Y(n_598) );
INVx1_ASAP7_75t_L g317 ( .A(n_295), .Y(n_317) );
AND2x4_ASAP7_75t_L g388 ( .A(n_295), .B(n_319), .Y(n_388) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx2_ASAP7_75t_L g442 ( .A(n_298), .Y(n_442) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx4f_ASAP7_75t_SL g338 ( .A(n_299), .Y(n_338) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_299), .Y(n_394) );
BUFx2_ASAP7_75t_L g420 ( .A(n_299), .Y(n_420) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_299), .Y(n_485) );
AND2x4_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_L g308 ( .A(n_301), .Y(n_308) );
AND2x4_ASAP7_75t_L g307 ( .A(n_302), .B(n_308), .Y(n_307) );
NAND2x1p5_ASAP7_75t_L g312 ( .A(n_302), .B(n_313), .Y(n_312) );
AND2x4_ASAP7_75t_L g385 ( .A(n_302), .B(n_386), .Y(n_385) );
BUFx4f_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g548 ( .A(n_306), .Y(n_548) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx12f_ASAP7_75t_L g395 ( .A(n_307), .Y(n_395) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_307), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B1(n_314), .B2(n_315), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_311), .A2(n_315), .B1(n_342), .B2(n_343), .Y(n_341) );
OAI22xp33_ASAP7_75t_L g482 ( .A1(n_311), .A2(n_483), .B1(n_484), .B2(n_486), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_311), .A2(n_559), .B1(n_560), .B2(n_561), .Y(n_558) );
BUFx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx4_ASAP7_75t_L g447 ( .A(n_312), .Y(n_447) );
BUFx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_316), .Y(n_450) );
OR2x6_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_SL g360 ( .A(n_325), .Y(n_360) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_344), .Y(n_325) );
NOR3xp33_ASAP7_75t_L g326 ( .A(n_327), .B(n_333), .C(n_341), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_329), .B1(n_331), .B2(n_332), .Y(n_327) );
OAI22xp5_ASAP7_75t_SL g475 ( .A1(n_329), .A2(n_436), .B1(n_476), .B2(n_477), .Y(n_475) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g434 ( .A(n_330), .Y(n_434) );
OAI221xp5_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_336), .B1(n_337), .B2(n_339), .C(n_340), .Y(n_333) );
INVx2_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g546 ( .A(n_335), .Y(n_546) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_350), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_349), .Y(n_345) );
INVx2_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
INVx4_ASAP7_75t_L g371 ( .A(n_348), .Y(n_371) );
OAI21xp33_ASAP7_75t_SL g408 ( .A1(n_348), .A2(n_409), .B(n_410), .Y(n_408) );
INVx4_ASAP7_75t_L g582 ( .A(n_348), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_355), .Y(n_350) );
BUFx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g510 ( .A(n_362), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_396), .B2(n_508), .Y(n_362) );
INVx2_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
XNOR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
NOR4xp75_ASAP7_75t_L g366 ( .A(n_367), .B(n_374), .C(n_380), .D(n_389), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_368), .B(n_372), .Y(n_367) );
INVx3_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx3_ASAP7_75t_L g423 ( .A(n_370), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx2_ASAP7_75t_L g437 ( .A(n_382), .Y(n_437) );
BUFx3_ASAP7_75t_L g607 ( .A(n_382), .Y(n_607) );
BUFx2_ASAP7_75t_L g411 ( .A(n_385), .Y(n_411) );
BUFx3_ASAP7_75t_L g531 ( .A(n_385), .Y(n_531) );
INVx1_ASAP7_75t_L g694 ( .A(n_385), .Y(n_694) );
INVx1_ASAP7_75t_SL g552 ( .A(n_387), .Y(n_552) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx2_ASAP7_75t_SL g481 ( .A(n_388), .Y(n_481) );
BUFx2_ASAP7_75t_SL g621 ( .A(n_388), .Y(n_621) );
OAI21xp5_ASAP7_75t_SL g389 ( .A1(n_390), .A2(n_392), .B(n_393), .Y(n_389) );
OAI21xp33_ASAP7_75t_L g478 ( .A1(n_390), .A2(n_479), .B(n_480), .Y(n_478) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g560 ( .A(n_394), .Y(n_560) );
BUFx6f_ASAP7_75t_L g692 ( .A(n_394), .Y(n_692) );
INVx1_ASAP7_75t_L g508 ( .A(n_396), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B1(n_427), .B2(n_507), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g426 ( .A(n_402), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_415), .Y(n_402) );
NOR3xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_408), .C(n_412), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_421), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVx1_ASAP7_75t_L g589 ( .A(n_418), .Y(n_589) );
INVx1_ASAP7_75t_L g600 ( .A(n_420), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_424), .Y(n_421) );
INVx1_ASAP7_75t_L g507 ( .A(n_427), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B1(n_468), .B2(n_469), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
XOR2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_467), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_451), .Y(n_430) );
NOR3xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_438), .C(n_444), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B1(n_435), .B2(n_436), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_434), .A2(n_605), .B1(n_606), .B2(n_607), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_436), .A2(n_554), .B1(n_555), .B2(n_557), .Y(n_553) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI21xp33_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B(n_441), .Y(n_438) );
BUFx3_ASAP7_75t_L g603 ( .A(n_443), .Y(n_603) );
INVx2_ASAP7_75t_L g701 ( .A(n_443), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_448), .B2(n_449), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_446), .A2(n_594), .B1(n_595), .B2(n_596), .Y(n_593) );
INVx3_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g596 ( .A(n_450), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_461), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g496 ( .A(n_454), .Y(n_496) );
INVx1_ASAP7_75t_SL g498 ( .A(n_455), .Y(n_498) );
INVx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_459), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_466), .Y(n_461) );
INVx4_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx4_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_487), .Y(n_473) );
NOR3xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_478), .C(n_482), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_485), .Y(n_484) );
NOR3xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_494), .C(n_499), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
BUFx2_ASAP7_75t_L g584 ( .A(n_492), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B1(n_497), .B2(n_498), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_502), .B1(n_503), .B2(n_504), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g666 ( .A(n_511), .Y(n_666) );
AOI22xp5_ASAP7_75t_SL g511 ( .A1(n_512), .A2(n_513), .B1(n_612), .B2(n_664), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OAI22xp5_ASAP7_75t_SL g513 ( .A1(n_514), .A2(n_575), .B1(n_610), .B2(n_611), .Y(n_513) );
INVx2_ASAP7_75t_SL g610 ( .A(n_514), .Y(n_610) );
AO22x2_ASAP7_75t_SL g514 ( .A1(n_515), .A2(n_541), .B1(n_542), .B2(n_574), .Y(n_514) );
INVx3_ASAP7_75t_L g574 ( .A(n_515), .Y(n_574) );
XOR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_540), .Y(n_515) );
NAND2x1_ASAP7_75t_SL g516 ( .A(n_517), .B(n_532), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_522), .Y(n_517) );
OAI21xp5_ASAP7_75t_SL g518 ( .A1(n_519), .A2(n_520), .B(n_521), .Y(n_518) );
NAND3xp33_ASAP7_75t_L g522 ( .A(n_523), .B(n_527), .C(n_530), .Y(n_522) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g624 ( .A(n_525), .Y(n_624) );
INVx5_ASAP7_75t_L g652 ( .A(n_525), .Y(n_652) );
INVx2_ASAP7_75t_L g690 ( .A(n_525), .Y(n_690) );
INVx4_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx4f_ASAP7_75t_L g626 ( .A(n_529), .Y(n_626) );
BUFx2_ASAP7_75t_L g649 ( .A(n_529), .Y(n_649) );
NOR2x1_ASAP7_75t_L g532 ( .A(n_533), .B(n_536), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
XOR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_573), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_562), .Y(n_543) );
NOR3xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_553), .C(n_558), .Y(n_544) );
OAI221xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B1(n_548), .B2(n_549), .C(n_550), .Y(n_545) );
OAI21xp5_ASAP7_75t_L g618 ( .A1(n_546), .A2(n_619), .B(n_620), .Y(n_618) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_563), .B(n_566), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_570), .Y(n_566) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g587 ( .A(n_569), .Y(n_587) );
INVx2_ASAP7_75t_L g686 ( .A(n_569), .Y(n_686) );
INVx1_ASAP7_75t_L g611 ( .A(n_575), .Y(n_611) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_SL g609 ( .A(n_577), .Y(n_609) );
AND2x2_ASAP7_75t_SL g577 ( .A(n_578), .B(n_592), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_585), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_583), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_590), .Y(n_585) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR3xp33_ASAP7_75t_SL g592 ( .A(n_593), .B(n_597), .C(n_604), .Y(n_592) );
OAI221xp5_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_599), .B1(n_600), .B2(n_601), .C(n_602), .Y(n_597) );
OAI21xp5_ASAP7_75t_SL g644 ( .A1(n_598), .A2(n_645), .B(n_646), .Y(n_644) );
CKINVDCx16_ASAP7_75t_R g664 ( .A(n_612), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B1(n_639), .B2(n_640), .Y(n_612) );
INVx2_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
INVx3_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
XOR2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_638), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_617), .B(n_628), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_622), .Y(n_617) );
NAND3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .C(n_627), .Y(n_622) );
NOR2x1_ASAP7_75t_L g628 ( .A(n_629), .B(n_634), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
XOR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_663), .Y(n_641) );
NAND3x1_ASAP7_75t_L g642 ( .A(n_643), .B(n_654), .C(n_659), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_644), .B(n_647), .Y(n_643) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .C(n_653), .Y(n_647) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_658), .Y(n_654) );
INVx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
NOR2x1_ASAP7_75t_L g668 ( .A(n_669), .B(n_673), .Y(n_668) );
OR2x2_ASAP7_75t_SL g717 ( .A(n_669), .B(n_674), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_670), .Y(n_705) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_671), .B(n_708), .Y(n_711) );
CKINVDCx16_ASAP7_75t_R g708 ( .A(n_672), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
OAI322xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_703), .A3(n_706), .B1(n_709), .B2(n_712), .C1(n_713), .C2(n_714), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND4xp75_ASAP7_75t_L g683 ( .A(n_684), .B(n_688), .C(n_695), .D(n_699), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
AND2x2_ASAP7_75t_SL g688 ( .A(n_689), .B(n_691), .Y(n_688) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
CKINVDCx16_ASAP7_75t_R g709 ( .A(n_710), .Y(n_709) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_716), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_717), .Y(n_716) );
endmodule