module fake_ariane_232_n_891 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_891);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_891;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_779;
wire n_731;
wire n_754;
wire n_871;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_369;
wire n_240;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_889;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_88),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_150),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_145),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_36),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_21),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_49),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_89),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_82),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_181),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_157),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_33),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_130),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_16),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_168),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_105),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_99),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_171),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_55),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_131),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_115),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_53),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_134),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_126),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_166),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_12),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_151),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_15),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_10),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_45),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_197),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_65),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_29),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_47),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_73),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_14),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_137),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_48),
.B(n_125),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_7),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_7),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_179),
.B(n_43),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_159),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_94),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_160),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_66),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_70),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_67),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_5),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_75),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_84),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_26),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_169),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_71),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_44),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_80),
.B(n_193),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_19),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_91),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_54),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_146),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_18),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_135),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_92),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_50),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_72),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_64),
.B(n_127),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_136),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_68),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_40),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_58),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_30),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_6),
.Y(n_274)
);

OAI22x1_ASAP7_75t_R g275 ( 
.A1(n_228),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_231),
.B(n_239),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_206),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_215),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_251),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_230),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_243),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g284 ( 
.A(n_201),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_205),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_0),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_209),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_201),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_221),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_206),
.Y(n_294)
);

BUFx12f_ASAP7_75t_L g295 ( 
.A(n_221),
.Y(n_295)
);

OA21x2_ASAP7_75t_L g296 ( 
.A1(n_202),
.A2(n_1),
.B(n_2),
.Y(n_296)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_204),
.A2(n_3),
.B(n_4),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_205),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_217),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_199),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_206),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_254),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_217),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_206),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_203),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_247),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_220),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_262),
.Y(n_308)
);

AND2x4_ASAP7_75t_L g309 ( 
.A(n_203),
.B(n_6),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_223),
.B(n_8),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_200),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_221),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_225),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_224),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_227),
.B(n_8),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_235),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_224),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_238),
.Y(n_318)
);

OA21x2_ASAP7_75t_L g319 ( 
.A1(n_246),
.A2(n_9),
.B(n_10),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_232),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_232),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_260),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_208),
.B(n_9),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_261),
.B(n_11),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_240),
.B(n_11),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_264),
.B(n_12),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_294),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_276),
.B(n_249),
.Y(n_330)
);

AOI21x1_ASAP7_75t_L g331 ( 
.A1(n_310),
.A2(n_266),
.B(n_265),
.Y(n_331)
);

INVxp33_ASAP7_75t_SL g332 ( 
.A(n_306),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_267),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_294),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_270),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_301),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_300),
.B(n_311),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_306),
.B(n_207),
.Y(n_340)
);

AND3x2_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_253),
.C(n_273),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_301),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_279),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_298),
.B(n_210),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_301),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_301),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

NAND3xp33_ASAP7_75t_L g348 ( 
.A(n_309),
.B(n_268),
.C(n_244),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_282),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_291),
.B(n_211),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_304),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_298),
.B(n_212),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_288),
.B(n_213),
.Y(n_353)
);

AOI21x1_ASAP7_75t_L g354 ( 
.A1(n_315),
.A2(n_258),
.B(n_241),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_283),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_305),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_304),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_304),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_286),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_304),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_305),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_305),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_317),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_317),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_290),
.B(n_214),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_317),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_317),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_287),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_278),
.B(n_13),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_288),
.B(n_216),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_280),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_323),
.B(n_218),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_299),
.B(n_219),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_323),
.Y(n_375)
);

CKINVDCx6p67_ASAP7_75t_R g376 ( 
.A(n_295),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_299),
.B(n_222),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_303),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_325),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_327),
.B(n_325),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_343),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g382 ( 
.A(n_372),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_372),
.Y(n_384)
);

BUFx6f_ASAP7_75t_SL g385 ( 
.A(n_375),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_327),
.B(n_326),
.Y(n_386)
);

BUFx8_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_348),
.A2(n_326),
.B1(n_319),
.B2(n_296),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_337),
.B(n_289),
.Y(n_389)
);

NAND2xp33_ASAP7_75t_SL g390 ( 
.A(n_330),
.B(n_262),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_337),
.B(n_295),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_339),
.A2(n_302),
.B1(n_324),
.B2(n_285),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_337),
.B(n_303),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_349),
.Y(n_394)
);

NOR3xp33_ASAP7_75t_L g395 ( 
.A(n_373),
.B(n_281),
.C(n_316),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_355),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_314),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_375),
.B(n_284),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_347),
.Y(n_399)
);

NAND3xp33_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_281),
.C(n_322),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_376),
.B(n_284),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_376),
.B(n_292),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_370),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_353),
.B(n_322),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_352),
.B(n_314),
.Y(n_405)
);

OR2x6_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_292),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_375),
.B(n_307),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_341),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_371),
.B(n_374),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_344),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_347),
.Y(n_411)
);

NAND2xp33_ASAP7_75t_L g412 ( 
.A(n_333),
.B(n_335),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_363),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_377),
.B(n_307),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_354),
.B(n_322),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_360),
.B(n_369),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_332),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_356),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_356),
.B(n_313),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_363),
.Y(n_420)
);

NAND3xp33_ASAP7_75t_L g421 ( 
.A(n_340),
.B(n_318),
.C(n_313),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_357),
.B(n_318),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_357),
.B(n_320),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_364),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_364),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_362),
.B(n_320),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_362),
.B(n_320),
.Y(n_428)
);

A2O1A1Ixp33_ASAP7_75t_L g429 ( 
.A1(n_368),
.A2(n_241),
.B(n_321),
.C(n_320),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_354),
.B(n_226),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_368),
.B(n_321),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_350),
.B(n_321),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_367),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_331),
.B(n_229),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_367),
.B(n_321),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_365),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_331),
.B(n_365),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_365),
.B(n_233),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_365),
.Y(n_439)
);

AO221x1_ASAP7_75t_L g440 ( 
.A1(n_332),
.A2(n_275),
.B1(n_297),
.B2(n_296),
.C(n_319),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_328),
.B(n_234),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_328),
.A2(n_319),
.B1(n_297),
.B2(n_296),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_329),
.B(n_236),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_329),
.B(n_237),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_334),
.B(n_245),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_334),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_336),
.B(n_248),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_336),
.B(n_250),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_338),
.B(n_308),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_SL g450 ( 
.A(n_338),
.B(n_308),
.Y(n_450)
);

AND2x6_ASAP7_75t_L g451 ( 
.A(n_401),
.B(n_342),
.Y(n_451)
);

OAI21xp33_ASAP7_75t_L g452 ( 
.A1(n_392),
.A2(n_256),
.B(n_252),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_426),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_413),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_420),
.Y(n_455)
);

CKINVDCx10_ASAP7_75t_R g456 ( 
.A(n_385),
.Y(n_456)
);

OAI21xp33_ASAP7_75t_L g457 ( 
.A1(n_389),
.A2(n_269),
.B(n_257),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_409),
.A2(n_297),
.B(n_359),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_389),
.B(n_409),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_426),
.Y(n_460)
);

O2A1O1Ixp33_ASAP7_75t_L g461 ( 
.A1(n_416),
.A2(n_361),
.B(n_359),
.C(n_358),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_384),
.B(n_13),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_412),
.B(n_271),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_391),
.B(n_272),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_419),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_430),
.A2(n_361),
.B(n_358),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_382),
.B(n_342),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_391),
.B(n_345),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_415),
.A2(n_351),
.B(n_346),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_410),
.B(n_345),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_430),
.A2(n_351),
.B(n_346),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_405),
.B(n_414),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_407),
.B(n_14),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_379),
.A2(n_110),
.B(n_196),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_386),
.B(n_15),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_415),
.A2(n_111),
.B(n_195),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_449),
.B(n_16),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_424),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_380),
.A2(n_393),
.B(n_437),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_417),
.Y(n_480)
);

A2O1A1Ixp33_ASAP7_75t_L g481 ( 
.A1(n_404),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_425),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_404),
.A2(n_113),
.B(n_20),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_381),
.B(n_17),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_403),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_485)
);

A2O1A1Ixp33_ASAP7_75t_L g486 ( 
.A1(n_395),
.A2(n_25),
.B(n_27),
.C(n_28),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_433),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_394),
.B(n_31),
.Y(n_488)
);

AND2x4_ASAP7_75t_SL g489 ( 
.A(n_417),
.B(n_32),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_403),
.B(n_34),
.Y(n_490)
);

BUFx4f_ASAP7_75t_L g491 ( 
.A(n_402),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_434),
.A2(n_400),
.B(n_442),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_390),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_396),
.B(n_198),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_408),
.B(n_35),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_387),
.B(n_37),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_438),
.A2(n_38),
.B(n_39),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_397),
.B(n_41),
.Y(n_498)
);

NOR2x1p5_ASAP7_75t_L g499 ( 
.A(n_385),
.B(n_194),
.Y(n_499)
);

AOI22x1_ASAP7_75t_SL g500 ( 
.A1(n_387),
.A2(n_440),
.B1(n_406),
.B2(n_418),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_406),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_434),
.A2(n_42),
.B(n_46),
.Y(n_502)
);

AO21x1_ASAP7_75t_L g503 ( 
.A1(n_423),
.A2(n_51),
.B(n_52),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_383),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_395),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_432),
.B(n_192),
.Y(n_506)
);

INVx11_ASAP7_75t_L g507 ( 
.A(n_398),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_399),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_422),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_427),
.Y(n_510)
);

O2A1O1Ixp33_ASAP7_75t_L g511 ( 
.A1(n_429),
.A2(n_411),
.B(n_445),
.C(n_444),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_450),
.Y(n_512)
);

CKINVDCx10_ASAP7_75t_R g513 ( 
.A(n_406),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_432),
.B(n_60),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_428),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_421),
.A2(n_61),
.B(n_62),
.Y(n_516)
);

OAI21xp33_ASAP7_75t_L g517 ( 
.A1(n_388),
.A2(n_63),
.B(n_69),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_441),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_441),
.B(n_74),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_447),
.A2(n_76),
.B(n_77),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_443),
.B(n_448),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_388),
.B(n_443),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_431),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_480),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_459),
.A2(n_439),
.B1(n_436),
.B2(n_446),
.Y(n_525)
);

A2O1A1Ixp33_ASAP7_75t_L g526 ( 
.A1(n_518),
.A2(n_522),
.B(n_517),
.C(n_472),
.Y(n_526)
);

INVx3_ASAP7_75t_SL g527 ( 
.A(n_489),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_521),
.A2(n_435),
.B(n_79),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_465),
.B(n_78),
.Y(n_529)
);

AND2x2_ASAP7_75t_SL g530 ( 
.A(n_496),
.B(n_81),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_510),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_456),
.Y(n_532)
);

AOI21xp33_ASAP7_75t_L g533 ( 
.A1(n_452),
.A2(n_83),
.B(n_85),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_460),
.Y(n_534)
);

AOI21x1_ASAP7_75t_L g535 ( 
.A1(n_458),
.A2(n_86),
.B(n_87),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_479),
.A2(n_90),
.B(n_93),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_492),
.A2(n_95),
.B(n_96),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_515),
.Y(n_538)
);

NOR2x1_ASAP7_75t_L g539 ( 
.A(n_499),
.B(n_97),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_463),
.A2(n_98),
.B(n_100),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_454),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_501),
.Y(n_542)
);

NAND2x1p5_ASAP7_75t_L g543 ( 
.A(n_491),
.B(n_101),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_491),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_477),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_509),
.B(n_106),
.Y(n_546)
);

OAI21x1_ASAP7_75t_L g547 ( 
.A1(n_469),
.A2(n_107),
.B(n_108),
.Y(n_547)
);

AO31x2_ASAP7_75t_L g548 ( 
.A1(n_503),
.A2(n_109),
.A3(n_114),
.B(n_116),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_462),
.B(n_117),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_455),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_490),
.B(n_118),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_464),
.A2(n_119),
.B(n_120),
.Y(n_552)
);

AO21x1_ASAP7_75t_L g553 ( 
.A1(n_476),
.A2(n_121),
.B(n_122),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_477),
.B(n_123),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_513),
.Y(n_555)
);

A2O1A1Ixp33_ASAP7_75t_L g556 ( 
.A1(n_475),
.A2(n_124),
.B(n_128),
.C(n_129),
.Y(n_556)
);

AO31x2_ASAP7_75t_L g557 ( 
.A1(n_466),
.A2(n_132),
.A3(n_133),
.B(n_138),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_495),
.B(n_139),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_523),
.Y(n_559)
);

AOI21x1_ASAP7_75t_L g560 ( 
.A1(n_488),
.A2(n_140),
.B(n_141),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_495),
.B(n_142),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_493),
.B(n_143),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_451),
.B(n_144),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_451),
.B(n_147),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_460),
.Y(n_565)
);

OR2x6_ASAP7_75t_L g566 ( 
.A(n_513),
.B(n_148),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_451),
.B(n_149),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_451),
.B(n_152),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_506),
.A2(n_153),
.B(n_154),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_468),
.A2(n_155),
.B(n_158),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_478),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_473),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_460),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_482),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_498),
.A2(n_165),
.B(n_167),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_487),
.Y(n_576)
);

A2O1A1Ixp33_ASAP7_75t_L g577 ( 
.A1(n_457),
.A2(n_170),
.B(n_172),
.C(n_173),
.Y(n_577)
);

AND3x2_ASAP7_75t_L g578 ( 
.A(n_456),
.B(n_500),
.C(n_507),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_512),
.B(n_470),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_484),
.B(n_174),
.Y(n_580)
);

OAI21x1_ASAP7_75t_L g581 ( 
.A1(n_471),
.A2(n_176),
.B(n_177),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_504),
.B(n_180),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_494),
.A2(n_182),
.B(n_183),
.Y(n_583)
);

BUFx4f_ASAP7_75t_L g584 ( 
.A(n_530),
.Y(n_584)
);

OAI21x1_ASAP7_75t_L g585 ( 
.A1(n_547),
.A2(n_502),
.B(n_497),
.Y(n_585)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_535),
.A2(n_483),
.B(n_519),
.Y(n_586)
);

AO21x1_ASAP7_75t_L g587 ( 
.A1(n_537),
.A2(n_516),
.B(n_485),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_541),
.Y(n_588)
);

BUFx8_ASAP7_75t_SL g589 ( 
.A(n_532),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_531),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_524),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_538),
.B(n_504),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_526),
.A2(n_511),
.B(n_461),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_542),
.B(n_467),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_579),
.Y(n_595)
);

OA21x2_ASAP7_75t_L g596 ( 
.A1(n_536),
.A2(n_583),
.B(n_581),
.Y(n_596)
);

AO21x2_ASAP7_75t_L g597 ( 
.A1(n_580),
.A2(n_514),
.B(n_486),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_551),
.A2(n_474),
.B(n_520),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_555),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_544),
.A2(n_508),
.B1(n_505),
.B2(n_453),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_534),
.Y(n_601)
);

OA21x2_ASAP7_75t_L g602 ( 
.A1(n_553),
.A2(n_481),
.B(n_508),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_566),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_559),
.B(n_453),
.Y(n_604)
);

OAI21x1_ASAP7_75t_L g605 ( 
.A1(n_528),
.A2(n_560),
.B(n_552),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_554),
.B(n_184),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_538),
.B(n_185),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_563),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_554),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_563),
.Y(n_610)
);

OAI21x1_ASAP7_75t_L g611 ( 
.A1(n_575),
.A2(n_190),
.B(n_191),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_550),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_534),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_527),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_571),
.Y(n_615)
);

AOI21xp33_ASAP7_75t_L g616 ( 
.A1(n_561),
.A2(n_558),
.B(n_549),
.Y(n_616)
);

OA21x2_ASAP7_75t_L g617 ( 
.A1(n_577),
.A2(n_533),
.B(n_540),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_576),
.Y(n_618)
);

OA21x2_ASAP7_75t_L g619 ( 
.A1(n_529),
.A2(n_546),
.B(n_570),
.Y(n_619)
);

OA21x2_ASAP7_75t_L g620 ( 
.A1(n_582),
.A2(n_556),
.B(n_525),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_574),
.B(n_566),
.Y(n_621)
);

OAI21x1_ASAP7_75t_L g622 ( 
.A1(n_564),
.A2(n_568),
.B(n_567),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_534),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_572),
.A2(n_569),
.B(n_543),
.Y(n_624)
);

OAI21x1_ASAP7_75t_L g625 ( 
.A1(n_562),
.A2(n_573),
.B(n_545),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_557),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_573),
.B(n_539),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_565),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_557),
.Y(n_629)
);

AO21x2_ASAP7_75t_L g630 ( 
.A1(n_557),
.A2(n_548),
.B(n_565),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g631 ( 
.A1(n_548),
.A2(n_565),
.B(n_578),
.Y(n_631)
);

OAI21x1_ASAP7_75t_L g632 ( 
.A1(n_548),
.A2(n_547),
.B(n_535),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_534),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_595),
.B(n_590),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_618),
.Y(n_635)
);

CKINVDCx6p67_ASAP7_75t_R g636 ( 
.A(n_599),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_588),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_614),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g639 ( 
.A(n_591),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_584),
.B(n_606),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_633),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_584),
.A2(n_606),
.B1(n_608),
.B2(n_610),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_633),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_588),
.Y(n_644)
);

AOI21x1_ASAP7_75t_L g645 ( 
.A1(n_632),
.A2(n_598),
.B(n_617),
.Y(n_645)
);

AOI22x1_ASAP7_75t_L g646 ( 
.A1(n_593),
.A2(n_587),
.B1(n_627),
.B2(n_610),
.Y(n_646)
);

BUFx2_ASAP7_75t_SL g647 ( 
.A(n_613),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_612),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_633),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_612),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_615),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_608),
.B(n_610),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_SL g653 ( 
.A1(n_584),
.A2(n_606),
.B1(n_603),
.B2(n_621),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_613),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_589),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_615),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_592),
.Y(n_657)
);

AOI21x1_ASAP7_75t_L g658 ( 
.A1(n_632),
.A2(n_617),
.B(n_629),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_594),
.Y(n_659)
);

OAI21x1_ASAP7_75t_L g660 ( 
.A1(n_605),
.A2(n_585),
.B(n_586),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_604),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_626),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_633),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_608),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_589),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_621),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_623),
.Y(n_667)
);

AO21x2_ASAP7_75t_L g668 ( 
.A1(n_629),
.A2(n_630),
.B(n_605),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_602),
.Y(n_669)
);

NAND2x1p5_ASAP7_75t_L g670 ( 
.A(n_627),
.B(n_624),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_623),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_602),
.Y(n_672)
);

BUFx4f_ASAP7_75t_SL g673 ( 
.A(n_599),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_628),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_601),
.B(n_630),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_603),
.B(n_606),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_661),
.B(n_601),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_666),
.Y(n_678)
);

INVxp67_ASAP7_75t_R g679 ( 
.A(n_640),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_662),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_640),
.B(n_631),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_662),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_635),
.B(n_630),
.Y(n_683)
);

NAND3xp33_ASAP7_75t_L g684 ( 
.A(n_646),
.B(n_616),
.C(n_609),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_669),
.B(n_631),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_669),
.B(n_602),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_659),
.B(n_600),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_663),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_663),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_657),
.B(n_607),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_670),
.B(n_625),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_639),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_670),
.B(n_625),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_634),
.B(n_624),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_654),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_670),
.B(n_597),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_653),
.A2(n_597),
.B1(n_617),
.B2(n_620),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_675),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_637),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_637),
.Y(n_700)
);

AND2x4_ASAP7_75t_SL g701 ( 
.A(n_636),
.B(n_611),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_675),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_672),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_672),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_664),
.B(n_620),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_648),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_664),
.B(n_620),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_648),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_638),
.B(n_611),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_668),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_668),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_664),
.B(n_622),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_668),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_658),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_636),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_652),
.B(n_622),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_663),
.Y(n_717)
);

AO31x2_ASAP7_75t_L g718 ( 
.A1(n_650),
.A2(n_596),
.A3(n_619),
.B(n_586),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_667),
.B(n_596),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_638),
.B(n_654),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_674),
.B(n_619),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_663),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_676),
.B(n_619),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_663),
.Y(n_724)
);

OAI222xp33_ASAP7_75t_L g725 ( 
.A1(n_642),
.A2(n_585),
.B1(n_596),
.B2(n_644),
.C1(n_646),
.C2(n_651),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_667),
.B(n_671),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_678),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_706),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_692),
.B(n_671),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_677),
.B(n_671),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_720),
.B(n_695),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_706),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_698),
.B(n_652),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_695),
.B(n_667),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_686),
.B(n_658),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_686),
.B(n_645),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_681),
.B(n_683),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_SL g738 ( 
.A1(n_684),
.A2(n_673),
.B1(n_647),
.B2(n_656),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_698),
.B(n_702),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_683),
.B(n_645),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_708),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_687),
.B(n_641),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_708),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_681),
.B(n_641),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_690),
.B(n_643),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_702),
.B(n_660),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_705),
.B(n_660),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_705),
.B(n_643),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_724),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_681),
.B(n_649),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_707),
.B(n_649),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_680),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_699),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_699),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_726),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_717),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_707),
.B(n_656),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_719),
.B(n_647),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_724),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_700),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_681),
.A2(n_655),
.B1(n_665),
.B2(n_685),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_700),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_694),
.B(n_655),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_682),
.Y(n_764)
);

INVxp67_ASAP7_75t_SL g765 ( 
.A(n_721),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_727),
.B(n_723),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_755),
.B(n_717),
.Y(n_767)
);

OR2x6_ASAP7_75t_L g768 ( 
.A(n_744),
.B(n_750),
.Y(n_768)
);

NAND2x1p5_ASAP7_75t_L g769 ( 
.A(n_749),
.B(n_688),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_733),
.B(n_716),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_735),
.B(n_758),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_746),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_728),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_745),
.B(n_716),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_748),
.B(n_751),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_735),
.B(n_719),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_739),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_739),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_SL g779 ( 
.A1(n_738),
.A2(n_701),
.B(n_725),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_728),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_732),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_733),
.B(n_716),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_741),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_759),
.Y(n_784)
);

NOR2x1_ASAP7_75t_L g785 ( 
.A(n_763),
.B(n_709),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_743),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_748),
.B(n_679),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_744),
.B(n_693),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_730),
.B(n_712),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_751),
.B(n_679),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_758),
.B(n_736),
.Y(n_791)
);

INVxp67_ASAP7_75t_SL g792 ( 
.A(n_765),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_736),
.B(n_685),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_740),
.B(n_737),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_729),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_773),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_795),
.Y(n_797)
);

INVxp67_ASAP7_75t_SL g798 ( 
.A(n_792),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_794),
.B(n_740),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_794),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_773),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_791),
.B(n_771),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_768),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_781),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_772),
.B(n_746),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_783),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_780),
.Y(n_807)
);

NOR4xp25_ASAP7_75t_L g808 ( 
.A(n_779),
.B(n_731),
.C(n_761),
.D(n_742),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_786),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_791),
.B(n_747),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_SL g811 ( 
.A(n_784),
.B(n_715),
.Y(n_811)
);

OAI32xp33_ASAP7_75t_L g812 ( 
.A1(n_808),
.A2(n_772),
.A3(n_774),
.B1(n_778),
.B2(n_777),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_798),
.A2(n_792),
.B(n_785),
.C(n_766),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_802),
.B(n_810),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_807),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_800),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_800),
.A2(n_788),
.B1(n_768),
.B2(n_770),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_802),
.B(n_771),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_797),
.B(n_793),
.Y(n_819)
);

INVx1_ASAP7_75t_SL g820 ( 
.A(n_811),
.Y(n_820)
);

NAND2xp33_ASAP7_75t_R g821 ( 
.A(n_805),
.B(n_788),
.Y(n_821)
);

OAI22xp33_ASAP7_75t_L g822 ( 
.A1(n_821),
.A2(n_788),
.B1(n_768),
.B2(n_803),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_815),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_812),
.A2(n_803),
.B(n_715),
.C(n_805),
.Y(n_824)
);

INVx1_ASAP7_75t_SL g825 ( 
.A(n_820),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_819),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_813),
.B(n_806),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_827),
.B(n_813),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_826),
.Y(n_829)
);

AOI32xp33_ASAP7_75t_L g830 ( 
.A1(n_825),
.A2(n_817),
.A3(n_814),
.B1(n_818),
.B2(n_809),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_823),
.Y(n_831)
);

OAI32xp33_ASAP7_75t_L g832 ( 
.A1(n_824),
.A2(n_821),
.A3(n_816),
.B1(n_804),
.B2(n_767),
.Y(n_832)
);

AOI221xp5_ASAP7_75t_L g833 ( 
.A1(n_822),
.A2(n_807),
.B1(n_697),
.B2(n_801),
.C(n_793),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_824),
.B(n_799),
.Y(n_834)
);

OAI321xp33_ASAP7_75t_L g835 ( 
.A1(n_828),
.A2(n_789),
.A3(n_734),
.B1(n_801),
.B2(n_790),
.C(n_787),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_829),
.B(n_665),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_834),
.B(n_832),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_831),
.B(n_799),
.Y(n_838)
);

AOI22x1_ASAP7_75t_L g839 ( 
.A1(n_837),
.A2(n_830),
.B1(n_769),
.B2(n_810),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_836),
.A2(n_833),
.B1(n_796),
.B2(n_744),
.Y(n_840)
);

AND2x2_ASAP7_75t_SL g841 ( 
.A(n_840),
.B(n_838),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_839),
.Y(n_842)
);

NOR2x1_ASAP7_75t_L g843 ( 
.A(n_839),
.B(n_835),
.Y(n_843)
);

NOR2x1_ASAP7_75t_L g844 ( 
.A(n_842),
.B(n_784),
.Y(n_844)
);

NAND4xp75_ASAP7_75t_L g845 ( 
.A(n_843),
.B(n_776),
.C(n_696),
.D(n_691),
.Y(n_845)
);

OAI322xp33_ASAP7_75t_L g846 ( 
.A1(n_841),
.A2(n_782),
.A3(n_714),
.B1(n_776),
.B2(n_775),
.C1(n_769),
.C2(n_749),
.Y(n_846)
);

AO22x2_ASAP7_75t_L g847 ( 
.A1(n_842),
.A2(n_796),
.B1(n_749),
.B2(n_689),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_841),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_841),
.B(n_747),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_848),
.B(n_756),
.Y(n_850)
);

NOR2x1_ASAP7_75t_L g851 ( 
.A(n_844),
.B(n_722),
.Y(n_851)
);

OR3x2_ASAP7_75t_L g852 ( 
.A(n_845),
.B(n_714),
.C(n_701),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_847),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_SL g854 ( 
.A1(n_846),
.A2(n_759),
.B1(n_689),
.B2(n_688),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_849),
.B(n_759),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_853),
.A2(n_722),
.B(n_688),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_850),
.A2(n_759),
.B(n_722),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_852),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_854),
.A2(n_750),
.B1(n_712),
.B2(n_691),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_855),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_851),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_856),
.A2(n_750),
.B(n_693),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_860),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_861),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_858),
.A2(n_857),
.B(n_859),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_861),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_861),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_858),
.A2(n_696),
.B1(n_757),
.B2(n_737),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_861),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_860),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_860),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_866),
.B(n_737),
.Y(n_872)
);

AOI21xp33_ASAP7_75t_L g873 ( 
.A1(n_869),
.A2(n_762),
.B(n_754),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_863),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_871),
.Y(n_875)
);

AO21x2_ASAP7_75t_L g876 ( 
.A1(n_864),
.A2(n_867),
.B(n_870),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_865),
.A2(n_713),
.B1(n_711),
.B2(n_710),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_868),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_862),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_866),
.B(n_718),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_874),
.A2(n_713),
.B1(n_711),
.B2(n_710),
.Y(n_881)
);

OA21x2_ASAP7_75t_L g882 ( 
.A1(n_875),
.A2(n_760),
.B(n_753),
.Y(n_882)
);

INVxp33_ASAP7_75t_SL g883 ( 
.A(n_872),
.Y(n_883)
);

OAI222xp33_ASAP7_75t_L g884 ( 
.A1(n_879),
.A2(n_877),
.B1(n_878),
.B2(n_880),
.C1(n_876),
.C2(n_873),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_874),
.A2(n_757),
.B(n_703),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_876),
.A2(n_703),
.B(n_704),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_883),
.B(n_718),
.Y(n_887)
);

AO21x2_ASAP7_75t_L g888 ( 
.A1(n_884),
.A2(n_704),
.B(n_764),
.Y(n_888)
);

INVxp67_ASAP7_75t_L g889 ( 
.A(n_888),
.Y(n_889)
);

AOI221xp5_ASAP7_75t_L g890 ( 
.A1(n_889),
.A2(n_887),
.B1(n_886),
.B2(n_881),
.C(n_885),
.Y(n_890)
);

AOI21xp33_ASAP7_75t_SL g891 ( 
.A1(n_890),
.A2(n_882),
.B(n_752),
.Y(n_891)
);


endmodule