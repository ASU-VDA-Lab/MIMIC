module fake_netlist_6_4648_n_10 (n_1, n_0, n_10);

input n_1;
input n_0;

output n_10;

wire n_7;
wire n_6;
wire n_4;
wire n_2;
wire n_5;
wire n_3;
wire n_9;
wire n_8;

INVx4_ASAP7_75t_L g2 ( 
.A(n_1),
.Y(n_2)
);

BUFx3_ASAP7_75t_L g3 ( 
.A(n_1),
.Y(n_3)
);

OAI21x1_ASAP7_75t_L g4 ( 
.A1(n_2),
.A2(n_3),
.B(n_0),
.Y(n_4)
);

BUFx2_ASAP7_75t_L g5 ( 
.A(n_3),
.Y(n_5)
);

AOI33xp33_ASAP7_75t_L g6 ( 
.A1(n_5),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_4),
.B3(n_3),
.Y(n_6)
);

AO22x2_ASAP7_75t_L g7 ( 
.A1(n_6),
.A2(n_2),
.B1(n_4),
.B2(n_1),
.Y(n_7)
);

AOI21xp33_ASAP7_75t_L g8 ( 
.A1(n_7),
.A2(n_2),
.B(n_5),
.Y(n_8)
);

AOI22x1_ASAP7_75t_L g9 ( 
.A1(n_8),
.A2(n_7),
.B1(n_4),
.B2(n_0),
.Y(n_9)
);

OAI221xp5_ASAP7_75t_R g10 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_8),
.C(n_7),
.Y(n_10)
);


endmodule