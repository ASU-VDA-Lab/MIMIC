module fake_ariane_1162_n_2959 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_598, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_620, n_228, n_325, n_276, n_93, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_588, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_2959);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_588;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_2959;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_2484;
wire n_2866;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_2879;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_2663;
wire n_2914;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_2950;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_2885;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_2867;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1654;
wire n_1560;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2326;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2926;
wire n_2620;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2549;
wire n_2499;
wire n_762;
wire n_1253;
wire n_1661;
wire n_1468;
wire n_2791;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2952;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_2922;
wire n_2871;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_2628;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_2294;
wire n_2274;
wire n_2895;
wire n_2903;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_2924;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_2811;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_2937;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2783;
wire n_2599;
wire n_699;
wire n_727;
wire n_2075;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_2496;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_2853;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_957;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_845;
wire n_2894;
wire n_2300;
wire n_2949;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_2946;
wire n_1734;
wire n_1860;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_704;
wire n_2958;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_1191;
wire n_2492;
wire n_2939;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_2928;
wire n_943;
wire n_1118;
wire n_678;
wire n_2905;
wire n_2884;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_2936;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_858;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_2947;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2820;
wire n_2613;
wire n_1165;
wire n_2934;
wire n_1641;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_2935;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_2920;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_683;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_1193;
wire n_1345;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_2938;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_2931;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_2828;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_2927;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_2951;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_2858;
wire n_972;
wire n_2251;
wire n_2923;
wire n_2843;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2872;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_1024;
wire n_830;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_2868;
wire n_2723;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_2012;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_2948;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_2897;
wire n_1322;
wire n_2583;
wire n_2918;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_701;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_1459;
wire n_840;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_2206;
wire n_997;
wire n_635;
wire n_1902;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2933;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_709;
wire n_2917;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_2957;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_1043;
wire n_2869;
wire n_1923;
wire n_2955;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2275;
wire n_2205;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2940;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2915;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_1308;
wire n_796;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g623 ( 
.A(n_130),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_557),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_69),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_222),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_30),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_34),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_597),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_132),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_289),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_525),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_387),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_603),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_587),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_605),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_500),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_592),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_6),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_83),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_494),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_499),
.Y(n_642)
);

BUFx8_ASAP7_75t_SL g643 ( 
.A(n_369),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_363),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_164),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_64),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_420),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_111),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_361),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_596),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_307),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_243),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_137),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_52),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_61),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_595),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_283),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_563),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_543),
.Y(n_659)
);

CKINVDCx16_ASAP7_75t_R g660 ( 
.A(n_550),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_273),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_386),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_27),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_433),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_604),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_401),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_211),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_160),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_400),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_582),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_109),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_438),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_505),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_350),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_316),
.Y(n_675)
);

BUFx5_ASAP7_75t_L g676 ( 
.A(n_591),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_587),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_102),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_519),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_81),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_149),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_77),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_267),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_254),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_256),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_586),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_122),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_614),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_534),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_256),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_74),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_82),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_478),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_222),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_385),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_588),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_535),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_593),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_543),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_1),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_601),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_589),
.Y(n_702)
);

CKINVDCx16_ASAP7_75t_R g703 ( 
.A(n_602),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_426),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_608),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_172),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_586),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_412),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_591),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_585),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_9),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_606),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_488),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_119),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_553),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_583),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_365),
.Y(n_717)
);

BUFx8_ASAP7_75t_SL g718 ( 
.A(n_366),
.Y(n_718)
);

CKINVDCx16_ASAP7_75t_R g719 ( 
.A(n_310),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_266),
.Y(n_720)
);

BUFx5_ASAP7_75t_L g721 ( 
.A(n_351),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_129),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_555),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_23),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_300),
.Y(n_725)
);

BUFx10_ASAP7_75t_L g726 ( 
.A(n_57),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_307),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_171),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_472),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_140),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_494),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_1),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_269),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_313),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_379),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_147),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_392),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_295),
.Y(n_738)
);

CKINVDCx12_ASAP7_75t_R g739 ( 
.A(n_5),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_532),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_250),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_215),
.Y(n_742)
);

CKINVDCx20_ASAP7_75t_R g743 ( 
.A(n_76),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_544),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_584),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_171),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_523),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_346),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_210),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_190),
.Y(n_750)
);

BUFx8_ASAP7_75t_SL g751 ( 
.A(n_375),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_212),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_46),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_89),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_193),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_126),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_599),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_46),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_387),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_531),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_363),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_197),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_278),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_389),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_275),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_583),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_485),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_376),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_170),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_507),
.Y(n_770)
);

BUFx5_ASAP7_75t_L g771 ( 
.A(n_335),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_347),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_490),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_49),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_38),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_240),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_362),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_172),
.Y(n_778)
);

INVxp67_ASAP7_75t_SL g779 ( 
.A(n_73),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_544),
.Y(n_780)
);

BUFx10_ASAP7_75t_L g781 ( 
.A(n_537),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_469),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_556),
.Y(n_783)
);

HB1xp67_ASAP7_75t_SL g784 ( 
.A(n_138),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_566),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_335),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_216),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_313),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_370),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_552),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_589),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_506),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_579),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_284),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_393),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_3),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_85),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_321),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_489),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_353),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_194),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_205),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_411),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_155),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_430),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_522),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_290),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_179),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_365),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_421),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_571),
.Y(n_811)
);

BUFx8_ASAP7_75t_SL g812 ( 
.A(n_362),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_259),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_234),
.Y(n_814)
);

BUFx10_ASAP7_75t_L g815 ( 
.A(n_496),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_478),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_348),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_476),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_78),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_22),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_441),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_262),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_170),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_355),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_578),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_579),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_461),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_483),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_147),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_272),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_447),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_594),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_413),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_107),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_319),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_108),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_194),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_265),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_598),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_484),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_468),
.Y(n_841)
);

BUFx10_ASAP7_75t_L g842 ( 
.A(n_260),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_546),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_434),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_160),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_345),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_212),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_411),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_388),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_611),
.Y(n_850)
);

BUFx10_ASAP7_75t_L g851 ( 
.A(n_20),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_402),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_607),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_553),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_117),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_436),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_36),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_462),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_620),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_567),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_590),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_622),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_600),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_354),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_9),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_534),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_161),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_235),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_657),
.B(n_2),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_692),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_628),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_628),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_707),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_635),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_688),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_635),
.Y(n_876)
);

NOR2xp67_ASAP7_75t_L g877 ( 
.A(n_624),
.B(n_0),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_643),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_646),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_794),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_646),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_750),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_750),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_658),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_676),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_718),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_776),
.Y(n_887)
);

INVx1_ASAP7_75t_SL g888 ( 
.A(n_784),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_751),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_641),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_776),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_641),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_676),
.Y(n_893)
);

BUFx10_ASAP7_75t_L g894 ( 
.A(n_658),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_812),
.Y(n_895)
);

INVxp67_ASAP7_75t_SL g896 ( 
.A(n_658),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_862),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_726),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_862),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_676),
.Y(n_900)
);

BUFx2_ASAP7_75t_SL g901 ( 
.A(n_859),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_676),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_676),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_676),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_843),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_676),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_721),
.Y(n_907)
);

NOR2xp67_ASAP7_75t_L g908 ( 
.A(n_624),
.B(n_0),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_658),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_664),
.Y(n_910)
);

CKINVDCx16_ASAP7_75t_R g911 ( 
.A(n_660),
.Y(n_911)
);

BUFx10_ASAP7_75t_L g912 ( 
.A(n_658),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_664),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_703),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_728),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_721),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_721),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_721),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_721),
.Y(n_919)
);

CKINVDCx16_ASAP7_75t_R g920 ( 
.A(n_719),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_868),
.Y(n_921)
);

NOR2xp67_ASAP7_75t_L g922 ( 
.A(n_630),
.B(n_2),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_728),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_625),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_721),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_721),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_771),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_771),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_771),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_771),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_771),
.Y(n_931)
);

INVx1_ASAP7_75t_SL g932 ( 
.A(n_735),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_626),
.Y(n_933)
);

INVxp33_ASAP7_75t_SL g934 ( 
.A(n_637),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_726),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_627),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_630),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_636),
.B(n_3),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_771),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_771),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_637),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_798),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_623),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_631),
.Y(n_944)
);

CKINVDCx16_ASAP7_75t_R g945 ( 
.A(n_726),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_798),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_798),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_629),
.Y(n_948)
);

CKINVDCx16_ASAP7_75t_R g949 ( 
.A(n_781),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_633),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_735),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_632),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_661),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_634),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_665),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_666),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_638),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_640),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_645),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_743),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_743),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_651),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_859),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_745),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_639),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_798),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_659),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_669),
.Y(n_968)
);

CKINVDCx16_ASAP7_75t_R g969 ( 
.A(n_781),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_662),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_674),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_639),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_888),
.Y(n_973)
);

NOR2xp67_ASAP7_75t_L g974 ( 
.A(n_897),
.B(n_647),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_897),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_896),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_899),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_893),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_899),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_900),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_902),
.Y(n_981)
);

INVxp67_ASAP7_75t_SL g982 ( 
.A(n_963),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_903),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_914),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_904),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_906),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_878),
.Y(n_987)
);

CKINVDCx16_ASAP7_75t_R g988 ( 
.A(n_945),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_916),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_878),
.Y(n_990)
);

CKINVDCx20_ASAP7_75t_R g991 ( 
.A(n_890),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_921),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_886),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_886),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_917),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_889),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_918),
.Y(n_997)
);

INVxp33_ASAP7_75t_SL g998 ( 
.A(n_889),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_919),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_925),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_926),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_895),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_929),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_930),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_895),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_931),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_901),
.B(n_647),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_939),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_940),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_890),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_892),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_943),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_944),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_952),
.Y(n_1014)
);

CKINVDCx16_ASAP7_75t_R g1015 ( 
.A(n_949),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_892),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_924),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_941),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_965),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_909),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_954),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_972),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_957),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_910),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_924),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_933),
.Y(n_1026)
);

INVxp33_ASAP7_75t_SL g1027 ( 
.A(n_914),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_933),
.Y(n_1028)
);

INVxp67_ASAP7_75t_SL g1029 ( 
.A(n_963),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_958),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_936),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_936),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_948),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_884),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_948),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_959),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_950),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_932),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1034),
.Y(n_1039)
);

BUFx12f_ASAP7_75t_L g1040 ( 
.A(n_987),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_1038),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_976),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_978),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_980),
.Y(n_1044)
);

INVx4_ASAP7_75t_L g1045 ( 
.A(n_1020),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_1034),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_1020),
.Y(n_1047)
);

INVx6_ASAP7_75t_L g1048 ( 
.A(n_982),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_SL g1049 ( 
.A1(n_991),
.A2(n_913),
.B1(n_915),
.B2(n_910),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_975),
.A2(n_869),
.B1(n_758),
.B2(n_773),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_981),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1029),
.B(n_898),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_975),
.B(n_950),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_983),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_985),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_974),
.B(n_898),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_986),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_989),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_987),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_995),
.Y(n_1060)
);

NAND2xp33_ASAP7_75t_L g1061 ( 
.A(n_977),
.B(n_798),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_997),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_999),
.Y(n_1063)
);

OA21x2_ASAP7_75t_L g1064 ( 
.A1(n_1000),
.A2(n_907),
.B(n_885),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1001),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1003),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1004),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1006),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1012),
.B(n_875),
.Y(n_1069)
);

OA21x2_ASAP7_75t_L g1070 ( 
.A1(n_1008),
.A2(n_907),
.B(n_885),
.Y(n_1070)
);

INVx5_ASAP7_75t_L g1071 ( 
.A(n_1009),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1013),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1014),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1021),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1023),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_1030),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_977),
.B(n_953),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_979),
.A2(n_758),
.B1(n_773),
.B2(n_745),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1007),
.B(n_973),
.Y(n_1079)
);

OA21x2_ASAP7_75t_L g1080 ( 
.A1(n_1036),
.A2(n_928),
.B(n_927),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_992),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_979),
.B(n_935),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1018),
.B(n_935),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_1019),
.B(n_934),
.Y(n_1084)
);

CKINVDCx14_ASAP7_75t_R g1085 ( 
.A(n_990),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1022),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_1017),
.Y(n_1087)
);

OA21x2_ASAP7_75t_L g1088 ( 
.A1(n_1017),
.A2(n_928),
.B(n_927),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1025),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_1025),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_1026),
.Y(n_1091)
);

OA21x2_ASAP7_75t_L g1092 ( 
.A1(n_1026),
.A2(n_942),
.B(n_962),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1028),
.A2(n_807),
.B1(n_808),
.B2(n_793),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1028),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_1031),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_1031),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1032),
.B(n_875),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1032),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1033),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_1033),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_1035),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1035),
.B(n_871),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_990),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_1037),
.Y(n_1104)
);

BUFx8_ASAP7_75t_SL g1105 ( 
.A(n_1010),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1037),
.A2(n_934),
.B1(n_908),
.B2(n_922),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_SL g1107 ( 
.A(n_1027),
.B(n_969),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_993),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_993),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_984),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_994),
.B(n_938),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_988),
.B(n_953),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_1015),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_994),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_996),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_SL g1116 ( 
.A1(n_1011),
.A2(n_915),
.B1(n_923),
.B2(n_913),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_998),
.A2(n_884),
.B(n_942),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_996),
.B(n_872),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1002),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1002),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1005),
.B(n_874),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1005),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_1016),
.B(n_938),
.Y(n_1123)
);

NOR2x1_ASAP7_75t_L g1124 ( 
.A(n_1024),
.B(n_877),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1012),
.B(n_876),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1034),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_982),
.B(n_955),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1079),
.B(n_955),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1076),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1076),
.Y(n_1130)
);

OAI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1050),
.A2(n_807),
.B1(n_808),
.B2(n_793),
.Y(n_1131)
);

OAI22xp33_ASAP7_75t_R g1132 ( 
.A1(n_1084),
.A2(n_779),
.B1(n_960),
.B2(n_951),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1065),
.A2(n_656),
.B1(n_642),
.B2(n_648),
.Y(n_1133)
);

OAI22xp33_ASAP7_75t_SL g1134 ( 
.A1(n_1050),
.A2(n_961),
.B1(n_880),
.B2(n_937),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1102),
.A2(n_968),
.B1(n_971),
.B2(n_956),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_1041),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1041),
.B(n_911),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1076),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1076),
.Y(n_1139)
);

OAI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1087),
.A2(n_861),
.B1(n_828),
.B2(n_968),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1076),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1042),
.B(n_956),
.Y(n_1142)
);

OAI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1087),
.A2(n_861),
.B1(n_828),
.B2(n_971),
.Y(n_1143)
);

AO22x2_ASAP7_75t_L g1144 ( 
.A1(n_1123),
.A2(n_964),
.B1(n_923),
.B2(n_671),
.Y(n_1144)
);

OAI22xp33_ASAP7_75t_SL g1145 ( 
.A1(n_1078),
.A2(n_920),
.B1(n_705),
.B2(n_724),
.Y(n_1145)
);

OAI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1087),
.A2(n_681),
.B1(n_863),
.B2(n_822),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1102),
.A2(n_684),
.B1(n_833),
.B2(n_761),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1056),
.A2(n_681),
.B1(n_678),
.B2(n_680),
.Y(n_1148)
);

OAI22xp33_ASAP7_75t_SL g1149 ( 
.A1(n_1078),
.A2(n_870),
.B1(n_873),
.B2(n_905),
.Y(n_1149)
);

OAI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1087),
.A2(n_642),
.B1(n_648),
.B2(n_644),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1042),
.B(n_636),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1048),
.B(n_685),
.Y(n_1152)
);

OAI22xp33_ASAP7_75t_SL g1153 ( 
.A1(n_1093),
.A2(n_649),
.B1(n_650),
.B2(n_644),
.Y(n_1153)
);

OA22x2_ASAP7_75t_L g1154 ( 
.A1(n_1093),
.A2(n_964),
.B1(n_970),
.B2(n_967),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_SL g1155 ( 
.A(n_1123),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1080),
.Y(n_1156)
);

OAI22xp33_ASAP7_75t_R g1157 ( 
.A1(n_1089),
.A2(n_667),
.B1(n_668),
.B2(n_663),
.Y(n_1157)
);

OR2x6_ASAP7_75t_L g1158 ( 
.A(n_1040),
.B(n_879),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1080),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1056),
.A2(n_683),
.B1(n_686),
.B2(n_675),
.Y(n_1160)
);

INVx8_ASAP7_75t_L g1161 ( 
.A(n_1040),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1090),
.B(n_881),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1056),
.A2(n_689),
.B1(n_690),
.B2(n_687),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1039),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1080),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1090),
.B(n_882),
.Y(n_1166)
);

AO22x2_ASAP7_75t_L g1167 ( 
.A1(n_1123),
.A2(n_694),
.B1(n_699),
.B2(n_685),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1056),
.A2(n_693),
.B1(n_695),
.B2(n_691),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1039),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_1100),
.B(n_883),
.Y(n_1170)
);

AO22x2_ASAP7_75t_L g1171 ( 
.A1(n_1123),
.A2(n_699),
.B1(n_765),
.B2(n_694),
.Y(n_1171)
);

AO22x2_ASAP7_75t_L g1172 ( 
.A1(n_1049),
.A2(n_767),
.B1(n_820),
.B2(n_765),
.Y(n_1172)
);

OAI22xp33_ASAP7_75t_SL g1173 ( 
.A1(n_1089),
.A2(n_653),
.B1(n_654),
.B2(n_652),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1068),
.A2(n_654),
.B1(n_655),
.B2(n_653),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_1113),
.Y(n_1175)
);

OAI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1087),
.A2(n_748),
.B1(n_860),
.B2(n_655),
.Y(n_1176)
);

OR2x6_ASAP7_75t_L g1177 ( 
.A(n_1113),
.B(n_887),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1100),
.B(n_891),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1080),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1126),
.Y(n_1180)
);

OAI22xp33_ASAP7_75t_SL g1181 ( 
.A1(n_1098),
.A2(n_860),
.B1(n_864),
.B2(n_748),
.Y(n_1181)
);

AND2x2_ASAP7_75t_SL g1182 ( 
.A(n_1107),
.B(n_831),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_SL g1183 ( 
.A1(n_1049),
.A2(n_739),
.B1(n_865),
.B2(n_864),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1126),
.Y(n_1184)
);

NAND2xp33_ASAP7_75t_SL g1185 ( 
.A(n_1091),
.B(n_865),
.Y(n_1185)
);

OR2x6_ASAP7_75t_L g1186 ( 
.A(n_1113),
.B(n_767),
.Y(n_1186)
);

OA22x2_ASAP7_75t_L g1187 ( 
.A1(n_1081),
.A2(n_868),
.B1(n_866),
.B2(n_697),
.Y(n_1187)
);

OAI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1091),
.A2(n_866),
.B1(n_821),
.B2(n_831),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1091),
.B(n_670),
.Y(n_1189)
);

AO22x2_ASAP7_75t_L g1190 ( 
.A1(n_1116),
.A2(n_821),
.B1(n_834),
.B2(n_820),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1072),
.Y(n_1191)
);

AO22x2_ASAP7_75t_L g1192 ( 
.A1(n_1116),
.A2(n_852),
.B1(n_834),
.B2(n_673),
.Y(n_1192)
);

OAI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1091),
.A2(n_852),
.B1(n_698),
.B2(n_700),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1072),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1081),
.B(n_781),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1086),
.B(n_815),
.Y(n_1196)
);

OAI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1091),
.A2(n_701),
.B1(n_702),
.B2(n_696),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1068),
.A2(n_706),
.B1(n_708),
.B2(n_704),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1086),
.B(n_711),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1083),
.A2(n_710),
.B1(n_712),
.B2(n_709),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1083),
.B(n_1111),
.Y(n_1201)
);

AO22x2_ASAP7_75t_L g1202 ( 
.A1(n_1111),
.A2(n_677),
.B1(n_679),
.B2(n_672),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1083),
.B(n_815),
.Y(n_1203)
);

OAI22xp33_ASAP7_75t_SL g1204 ( 
.A1(n_1098),
.A2(n_1099),
.B1(n_1094),
.B2(n_1104),
.Y(n_1204)
);

OR2x6_ASAP7_75t_L g1205 ( 
.A(n_1113),
.B(n_766),
.Y(n_1205)
);

OAI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1095),
.A2(n_1101),
.B1(n_1099),
.B2(n_1094),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1046),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1083),
.A2(n_713),
.B1(n_717),
.B2(n_715),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_SL g1209 ( 
.A1(n_1059),
.A2(n_736),
.B1(n_747),
.B2(n_725),
.Y(n_1209)
);

OAI22xp33_ASAP7_75t_R g1210 ( 
.A1(n_1114),
.A2(n_714),
.B1(n_716),
.B2(n_682),
.Y(n_1210)
);

OAI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1095),
.A2(n_722),
.B1(n_729),
.B2(n_720),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1118),
.A2(n_732),
.B1(n_733),
.B2(n_731),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1118),
.A2(n_738),
.B1(n_740),
.B2(n_737),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1082),
.B(n_741),
.Y(n_1214)
);

OAI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1095),
.A2(n_1101),
.B1(n_1104),
.B2(n_1108),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1046),
.Y(n_1216)
);

OR2x6_ASAP7_75t_L g1217 ( 
.A(n_1108),
.B(n_1109),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1074),
.Y(n_1218)
);

AO22x2_ASAP7_75t_L g1219 ( 
.A1(n_1111),
.A2(n_727),
.B1(n_730),
.B2(n_723),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_1105),
.Y(n_1220)
);

OAI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1095),
.A2(n_742),
.B1(n_753),
.B2(n_746),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1095),
.B(n_1101),
.Y(n_1222)
);

AO22x2_ASAP7_75t_L g1223 ( 
.A1(n_1111),
.A2(n_744),
.B1(n_749),
.B2(n_734),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1046),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1075),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1096),
.B(n_815),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1104),
.B(n_842),
.Y(n_1227)
);

XOR2xp5_ASAP7_75t_L g1228 ( 
.A(n_1059),
.B(n_754),
.Y(n_1228)
);

OAI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1101),
.A2(n_755),
.B1(n_757),
.B2(n_756),
.Y(n_1229)
);

XNOR2xp5_ASAP7_75t_L g1230 ( 
.A(n_1103),
.B(n_759),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1101),
.B(n_762),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1104),
.B(n_842),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_SL g1233 ( 
.A1(n_1103),
.A2(n_783),
.B1(n_792),
.B2(n_770),
.Y(n_1233)
);

AO22x2_ASAP7_75t_L g1234 ( 
.A1(n_1106),
.A2(n_1110),
.B1(n_1122),
.B2(n_1114),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1075),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1127),
.B(n_763),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1121),
.A2(n_769),
.B1(n_775),
.B2(n_764),
.Y(n_1237)
);

AO22x2_ASAP7_75t_L g1238 ( 
.A1(n_1110),
.A2(n_760),
.B1(n_768),
.B2(n_752),
.Y(n_1238)
);

OR2x6_ASAP7_75t_L g1239 ( 
.A(n_1108),
.B(n_785),
.Y(n_1239)
);

AO22x2_ASAP7_75t_L g1240 ( 
.A1(n_1122),
.A2(n_774),
.B1(n_778),
.B2(n_772),
.Y(n_1240)
);

INVxp33_ASAP7_75t_L g1241 ( 
.A(n_1112),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_SL g1242 ( 
.A1(n_1085),
.A2(n_801),
.B1(n_811),
.B2(n_789),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1108),
.A2(n_782),
.B1(n_786),
.B2(n_777),
.Y(n_1243)
);

INVx5_ASAP7_75t_L g1244 ( 
.A(n_1048),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1121),
.A2(n_787),
.B1(n_790),
.B2(n_788),
.Y(n_1245)
);

XNOR2xp5_ASAP7_75t_L g1246 ( 
.A(n_1119),
.B(n_791),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1108),
.A2(n_795),
.B1(n_797),
.B2(n_796),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1097),
.A2(n_803),
.B1(n_804),
.B2(n_800),
.Y(n_1248)
);

AND2x2_ASAP7_75t_SL g1249 ( 
.A(n_1109),
.B(n_780),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1115),
.B(n_842),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1109),
.Y(n_1251)
);

AOI22x1_ASAP7_75t_SL g1252 ( 
.A1(n_1115),
.A2(n_806),
.B1(n_809),
.B2(n_805),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1115),
.B(n_851),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1115),
.B(n_851),
.Y(n_1254)
);

AO22x2_ASAP7_75t_L g1255 ( 
.A1(n_1120),
.A2(n_802),
.B1(n_813),
.B2(n_799),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1109),
.B(n_817),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_R g1257 ( 
.A1(n_1120),
.A2(n_824),
.B1(n_841),
.B2(n_819),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1073),
.Y(n_1258)
);

AO22x2_ASAP7_75t_L g1259 ( 
.A1(n_1053),
.A2(n_845),
.B1(n_847),
.B2(n_844),
.Y(n_1259)
);

OR2x6_ASAP7_75t_L g1260 ( 
.A(n_1109),
.B(n_853),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1073),
.Y(n_1261)
);

OAI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1077),
.A2(n_814),
.B1(n_816),
.B2(n_810),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1052),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_1161),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1180),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1244),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1244),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1249),
.B(n_1054),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1136),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1137),
.B(n_1069),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1164),
.B(n_1063),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1169),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1244),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1184),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1201),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1222),
.B(n_1054),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1191),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1175),
.B(n_1069),
.Y(n_1278)
);

AND2x6_ASAP7_75t_L g1279 ( 
.A(n_1222),
.B(n_1156),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1194),
.Y(n_1280)
);

AND3x2_ASAP7_75t_L g1281 ( 
.A(n_1203),
.B(n_1131),
.C(n_1195),
.Y(n_1281)
);

BUFx10_ASAP7_75t_L g1282 ( 
.A(n_1189),
.Y(n_1282)
);

INVx6_ASAP7_75t_L g1283 ( 
.A(n_1161),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1258),
.B(n_1063),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1217),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1218),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1261),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1158),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1263),
.B(n_1043),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1225),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1207),
.B(n_1216),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1239),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_L g1293 ( 
.A(n_1135),
.B(n_1061),
.C(n_1044),
.Y(n_1293)
);

INVx4_ASAP7_75t_L g1294 ( 
.A(n_1217),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1128),
.B(n_1048),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1235),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1129),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1224),
.B(n_1063),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1130),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1152),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1151),
.Y(n_1301)
);

INVxp33_ASAP7_75t_L g1302 ( 
.A(n_1246),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1138),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1241),
.B(n_1048),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1139),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1141),
.Y(n_1306)
);

NAND2xp33_ASAP7_75t_L g1307 ( 
.A(n_1251),
.B(n_1227),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1189),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1157),
.A2(n_1092),
.B1(n_1088),
.B2(n_1055),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1158),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1239),
.Y(n_1311)
);

INVxp67_ASAP7_75t_L g1312 ( 
.A(n_1162),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1260),
.Y(n_1313)
);

INVxp33_ASAP7_75t_L g1314 ( 
.A(n_1246),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1256),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1232),
.Y(n_1316)
);

INVx5_ASAP7_75t_L g1317 ( 
.A(n_1260),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1170),
.B(n_1125),
.Y(n_1318)
);

OR2x6_ASAP7_75t_L g1319 ( 
.A(n_1177),
.B(n_1124),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1250),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1253),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1177),
.B(n_1125),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1159),
.Y(n_1323)
);

INVx4_ASAP7_75t_L g1324 ( 
.A(n_1186),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1210),
.A2(n_1092),
.B1(n_1088),
.B2(n_1055),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1166),
.B(n_1051),
.Y(n_1326)
);

NAND2xp33_ASAP7_75t_L g1327 ( 
.A(n_1254),
.B(n_1142),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1178),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1165),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1182),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1204),
.B(n_1063),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1236),
.B(n_1066),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_SL g1333 ( 
.A1(n_1259),
.A2(n_851),
.B1(n_867),
.B2(n_856),
.Y(n_1333)
);

INVx2_ASAP7_75t_SL g1334 ( 
.A(n_1196),
.Y(n_1334)
);

INVx6_ASAP7_75t_L g1335 ( 
.A(n_1186),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1179),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1199),
.Y(n_1337)
);

OR2x2_ASAP7_75t_L g1338 ( 
.A(n_1205),
.B(n_1051),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1205),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1255),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1226),
.B(n_1124),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1255),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1215),
.B(n_1043),
.Y(n_1343)
);

BUFx10_ASAP7_75t_L g1344 ( 
.A(n_1214),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1140),
.B(n_1057),
.Y(n_1345)
);

INVx5_ASAP7_75t_L g1346 ( 
.A(n_1206),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1143),
.B(n_1160),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1234),
.B(n_1057),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1234),
.Y(n_1349)
);

INVx5_ASAP7_75t_L g1350 ( 
.A(n_1185),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1231),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1240),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1187),
.Y(n_1353)
);

AND2x6_ASAP7_75t_L g1354 ( 
.A(n_1220),
.B(n_1043),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1257),
.A2(n_1092),
.B1(n_1088),
.B2(n_1067),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1155),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1167),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1197),
.B(n_1043),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1230),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1230),
.B(n_1092),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1167),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1240),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1171),
.Y(n_1363)
);

NAND3xp33_ASAP7_75t_L g1364 ( 
.A(n_1248),
.B(n_1044),
.C(n_1043),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1171),
.Y(n_1365)
);

BUFx8_ASAP7_75t_SL g1366 ( 
.A(n_1228),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1228),
.B(n_1066),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1163),
.B(n_1067),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1188),
.B(n_1088),
.Y(n_1369)
);

AO22x2_ASAP7_75t_L g1370 ( 
.A1(n_1144),
.A2(n_1132),
.B1(n_1219),
.B2(n_1202),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1242),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1262),
.Y(n_1372)
);

INVxp67_ASAP7_75t_L g1373 ( 
.A(n_1202),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1168),
.B(n_1044),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1193),
.B(n_1044),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1219),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1212),
.B(n_1058),
.C(n_1044),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1150),
.B(n_1058),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1223),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1183),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1238),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1147),
.B(n_1058),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1154),
.Y(n_1383)
);

NOR3xp33_ASAP7_75t_L g1384 ( 
.A(n_1176),
.B(n_823),
.C(n_818),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1238),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1172),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1172),
.Y(n_1387)
);

NAND2xp33_ASAP7_75t_L g1388 ( 
.A(n_1200),
.B(n_1058),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1190),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1146),
.B(n_1058),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1190),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1192),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1198),
.Y(n_1393)
);

BUFx4f_ASAP7_75t_L g1394 ( 
.A(n_1252),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1148),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_1144),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1133),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1211),
.Y(n_1398)
);

BUFx2_ASAP7_75t_L g1399 ( 
.A(n_1209),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1208),
.B(n_1060),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1213),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1221),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1237),
.B(n_1117),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1229),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1245),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1243),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1247),
.B(n_1060),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1174),
.B(n_825),
.Y(n_1408)
);

BUFx4f_ASAP7_75t_L g1409 ( 
.A(n_1134),
.Y(n_1409)
);

INVxp67_ASAP7_75t_L g1410 ( 
.A(n_1233),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1173),
.B(n_1060),
.Y(n_1411)
);

AND2x6_ASAP7_75t_L g1412 ( 
.A(n_1181),
.B(n_1060),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1153),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1145),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1149),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1180),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1249),
.A2(n_1060),
.B1(n_1062),
.B2(n_1045),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_SL g1418 ( 
.A(n_1249),
.B(n_1045),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1131),
.A2(n_1062),
.B1(n_1070),
.B2(n_1064),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1201),
.B(n_1117),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1164),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1244),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1136),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1136),
.B(n_826),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1249),
.B(n_1062),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1249),
.B(n_1062),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1164),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1136),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1164),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1164),
.B(n_1062),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1164),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1244),
.Y(n_1432)
);

INVx5_ASAP7_75t_L g1433 ( 
.A(n_1217),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1128),
.B(n_1045),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1180),
.Y(n_1435)
);

INVxp33_ASAP7_75t_L g1436 ( 
.A(n_1137),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1164),
.Y(n_1437)
);

OR2x6_ASAP7_75t_L g1438 ( 
.A(n_1161),
.B(n_1045),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1180),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1180),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1136),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1164),
.B(n_1064),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1164),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1249),
.B(n_1071),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1249),
.B(n_1071),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1164),
.Y(n_1446)
);

BUFx10_ASAP7_75t_L g1447 ( 
.A(n_1136),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1164),
.Y(n_1448)
);

CKINVDCx16_ASAP7_75t_R g1449 ( 
.A(n_1137),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1249),
.A2(n_1047),
.B1(n_1071),
.B2(n_1070),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1164),
.B(n_1064),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1131),
.A2(n_1064),
.B1(n_1070),
.B2(n_1071),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1244),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1164),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1164),
.B(n_1070),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1249),
.A2(n_1047),
.B1(n_1071),
.B2(n_829),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1136),
.B(n_827),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1180),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1180),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1180),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1164),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1367),
.B(n_830),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1265),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1449),
.B(n_832),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1287),
.Y(n_1465)
);

OA22x2_ASAP7_75t_L g1466 ( 
.A1(n_1281),
.A2(n_836),
.B1(n_837),
.B2(n_835),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1347),
.A2(n_1410),
.B1(n_1397),
.B2(n_1384),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1433),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1416),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1272),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1435),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1274),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1439),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1421),
.Y(n_1474)
);

AND2x6_ASAP7_75t_L g1475 ( 
.A(n_1285),
.B(n_884),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1427),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1433),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1429),
.Y(n_1478)
);

INVx8_ASAP7_75t_L g1479 ( 
.A(n_1433),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1431),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1318),
.B(n_1047),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1347),
.B(n_1047),
.Y(n_1482)
);

BUFx10_ASAP7_75t_L g1483 ( 
.A(n_1283),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1440),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1458),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1366),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1283),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1264),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1433),
.Y(n_1489)
);

NAND2x1p5_ASAP7_75t_L g1490 ( 
.A(n_1317),
.B(n_1071),
.Y(n_1490)
);

INVxp33_ASAP7_75t_L g1491 ( 
.A(n_1269),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1332),
.B(n_1295),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1437),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1285),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1443),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1436),
.B(n_1304),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1283),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1459),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1446),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1460),
.Y(n_1500)
);

BUFx4f_ASAP7_75t_L g1501 ( 
.A(n_1354),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1337),
.B(n_1312),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1448),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1277),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1280),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1312),
.B(n_838),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1286),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1317),
.B(n_966),
.Y(n_1508)
);

NAND2x1p5_ASAP7_75t_L g1509 ( 
.A(n_1317),
.B(n_966),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1454),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1304),
.B(n_839),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1290),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1332),
.B(n_840),
.Y(n_1513)
);

OAI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1418),
.A2(n_848),
.B1(n_849),
.B2(n_846),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1317),
.B(n_1322),
.Y(n_1515)
);

INVx8_ASAP7_75t_L g1516 ( 
.A(n_1354),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1461),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1326),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1410),
.A2(n_1384),
.B1(n_1418),
.B2(n_1399),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1322),
.B(n_850),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1339),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1296),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1348),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1359),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1295),
.B(n_1301),
.Y(n_1525)
);

AND2x6_ASAP7_75t_L g1526 ( 
.A(n_1285),
.B(n_909),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1423),
.B(n_854),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1348),
.Y(n_1528)
);

AND2x6_ASAP7_75t_L g1529 ( 
.A(n_1349),
.B(n_909),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1328),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1422),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1294),
.B(n_4),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1434),
.B(n_855),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1346),
.A2(n_858),
.B1(n_857),
.B2(n_6),
.Y(n_1534)
);

INVxp67_ASAP7_75t_L g1535 ( 
.A(n_1269),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1323),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1428),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1428),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1291),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1270),
.Y(n_1540)
);

INVxp67_ASAP7_75t_SL g1541 ( 
.A(n_1430),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1291),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1338),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1447),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1308),
.Y(n_1545)
);

INVx4_ASAP7_75t_L g1546 ( 
.A(n_1294),
.Y(n_1546)
);

INVx4_ASAP7_75t_L g1547 ( 
.A(n_1422),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1333),
.A2(n_912),
.B1(n_894),
.B2(n_946),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1356),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1360),
.B(n_894),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1284),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1434),
.B(n_894),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_1275),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1311),
.B(n_912),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1356),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1284),
.Y(n_1556)
);

INVx4_ASAP7_75t_L g1557 ( 
.A(n_1422),
.Y(n_1557)
);

AND2x6_ASAP7_75t_L g1558 ( 
.A(n_1453),
.B(n_909),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1278),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_1453),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1329),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1453),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1313),
.B(n_912),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1441),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1278),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1336),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1297),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1299),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1303),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1292),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1279),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1305),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1300),
.B(n_4),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1447),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1306),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1292),
.B(n_5),
.Y(n_1576)
);

AND2x6_ASAP7_75t_L g1577 ( 
.A(n_1420),
.B(n_1266),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1424),
.B(n_7),
.Y(n_1578)
);

BUFx4f_ASAP7_75t_L g1579 ( 
.A(n_1354),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1271),
.B(n_7),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1279),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1430),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1344),
.B(n_8),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1279),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1279),
.Y(n_1585)
);

AND2x6_ASAP7_75t_L g1586 ( 
.A(n_1420),
.B(n_909),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1271),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1438),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1279),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1344),
.B(n_1302),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1438),
.Y(n_1591)
);

AND2x6_ASAP7_75t_L g1592 ( 
.A(n_1266),
.B(n_946),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1340),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1356),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1342),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1331),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1371),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1314),
.B(n_8),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1442),
.Y(n_1599)
);

CKINVDCx20_ASAP7_75t_R g1600 ( 
.A(n_1288),
.Y(n_1600)
);

OR2x6_ASAP7_75t_L g1601 ( 
.A(n_1310),
.B(n_946),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1401),
.B(n_10),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1335),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_1438),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1457),
.B(n_612),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1442),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1345),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1315),
.Y(n_1608)
);

INVx8_ASAP7_75t_L g1609 ( 
.A(n_1354),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1298),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1335),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1298),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1268),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1267),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1354),
.Y(n_1615)
);

INVx5_ASAP7_75t_L g1616 ( 
.A(n_1335),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1324),
.B(n_10),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1357),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1316),
.B(n_1320),
.Y(n_1619)
);

AO22x2_ASAP7_75t_L g1620 ( 
.A1(n_1396),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1451),
.Y(n_1621)
);

NAND2x1p5_ASAP7_75t_L g1622 ( 
.A(n_1267),
.B(n_946),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1455),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1321),
.B(n_11),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1282),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1324),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1455),
.Y(n_1627)
);

BUFx6f_ASAP7_75t_L g1628 ( 
.A(n_1273),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1330),
.B(n_12),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1393),
.B(n_13),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1273),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1405),
.B(n_1309),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1282),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1380),
.B(n_14),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1309),
.B(n_15),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1373),
.B(n_15),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1361),
.Y(n_1637)
);

INVx4_ASAP7_75t_L g1638 ( 
.A(n_1432),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1334),
.B(n_16),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_SL g1640 ( 
.A1(n_1333),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1276),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1365),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1373),
.B(n_17),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1346),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1325),
.B(n_19),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1383),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1368),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1386),
.B(n_1376),
.Y(n_1648)
);

OAI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1346),
.A2(n_1395),
.B1(n_1402),
.B2(n_1398),
.Y(n_1649)
);

AND2x6_ASAP7_75t_L g1650 ( 
.A(n_1432),
.B(n_947),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1368),
.Y(n_1651)
);

INVxp67_ASAP7_75t_L g1652 ( 
.A(n_1425),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1319),
.B(n_21),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1319),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1386),
.B(n_22),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1319),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1350),
.Y(n_1657)
);

CKINVDCx8_ASAP7_75t_R g1658 ( 
.A(n_1412),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1382),
.Y(n_1659)
);

AOI22x1_ASAP7_75t_L g1660 ( 
.A1(n_1351),
.A2(n_947),
.B1(n_26),
.B2(n_24),
.Y(n_1660)
);

AO22x2_ASAP7_75t_L g1661 ( 
.A1(n_1396),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1661)
);

INVx4_ASAP7_75t_L g1662 ( 
.A(n_1350),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1325),
.B(n_25),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1512),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1467),
.A2(n_1378),
.B1(n_1406),
.B2(n_1404),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1607),
.B(n_1281),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1492),
.A2(n_1307),
.B(n_1327),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1519),
.B(n_1372),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1466),
.A2(n_1370),
.B1(n_1415),
.B2(n_1409),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1518),
.B(n_1381),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1467),
.B(n_1385),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1492),
.B(n_1355),
.Y(n_1672)
);

INVx8_ASAP7_75t_L g1673 ( 
.A(n_1479),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1519),
.B(n_1341),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1514),
.B(n_1372),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1539),
.B(n_1355),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1542),
.B(n_1374),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1530),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1463),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1597),
.B(n_1372),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1465),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1462),
.A2(n_1408),
.B1(n_1412),
.B2(n_1370),
.Y(n_1682)
);

INVx5_ASAP7_75t_L g1683 ( 
.A(n_1516),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1469),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1553),
.B(n_1524),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1471),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1470),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1516),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1502),
.B(n_1352),
.Y(n_1689)
);

INVx4_ASAP7_75t_L g1690 ( 
.A(n_1483),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1472),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1540),
.B(n_1362),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1540),
.B(n_1379),
.Y(n_1693)
);

NAND2x1p5_ASAP7_75t_L g1694 ( 
.A(n_1501),
.B(n_1350),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1474),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1553),
.B(n_1363),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_SL g1697 ( 
.A1(n_1640),
.A2(n_1413),
.B1(n_1415),
.B2(n_1392),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1496),
.B(n_1363),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1491),
.B(n_1413),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1476),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1514),
.B(n_1374),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1482),
.B(n_1350),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1473),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1538),
.B(n_1391),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1464),
.B(n_1370),
.Y(n_1705)
);

INVx3_ASAP7_75t_L g1706 ( 
.A(n_1516),
.Y(n_1706)
);

NOR3xp33_ASAP7_75t_L g1707 ( 
.A(n_1534),
.B(n_1411),
.C(n_1293),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1478),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1484),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1543),
.B(n_1391),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1480),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1466),
.A2(n_1409),
.B1(n_1412),
.B2(n_1414),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_1486),
.Y(n_1713)
);

A2O1A1Ixp33_ASAP7_75t_SL g1714 ( 
.A1(n_1583),
.A2(n_1411),
.B(n_1378),
.C(n_1353),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1535),
.B(n_1389),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1535),
.B(n_1289),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1537),
.B(n_1387),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1534),
.A2(n_1412),
.B1(n_1388),
.B2(n_1426),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1551),
.B(n_1556),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1537),
.B(n_1412),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1513),
.B(n_1382),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1493),
.Y(n_1722)
);

AND2x6_ASAP7_75t_L g1723 ( 
.A(n_1615),
.B(n_1417),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1579),
.B(n_1400),
.Y(n_1724)
);

NAND3xp33_ASAP7_75t_L g1725 ( 
.A(n_1644),
.B(n_1602),
.C(n_1513),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1590),
.B(n_1444),
.Y(n_1726)
);

NAND2xp33_ASAP7_75t_L g1727 ( 
.A(n_1615),
.B(n_1407),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1485),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1564),
.B(n_1445),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1653),
.B(n_1394),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1521),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1495),
.Y(n_1732)
);

INVxp67_ASAP7_75t_L g1733 ( 
.A(n_1570),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1498),
.Y(n_1734)
);

INVx2_ASAP7_75t_SL g1735 ( 
.A(n_1616),
.Y(n_1735)
);

OAI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1635),
.A2(n_1390),
.B1(n_1456),
.B2(n_1407),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_L g1737 ( 
.A(n_1479),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1579),
.B(n_1390),
.Y(n_1738)
);

AND2x4_ASAP7_75t_SL g1739 ( 
.A(n_1483),
.B(n_1515),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1549),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1488),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1663),
.A2(n_1452),
.B1(n_1419),
.B2(n_1375),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1615),
.B(n_1375),
.Y(n_1743)
);

INVx3_ASAP7_75t_L g1744 ( 
.A(n_1609),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1499),
.Y(n_1745)
);

INVx4_ASAP7_75t_L g1746 ( 
.A(n_1479),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1500),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1503),
.Y(n_1748)
);

NAND2xp33_ASAP7_75t_L g1749 ( 
.A(n_1609),
.B(n_1657),
.Y(n_1749)
);

BUFx3_ASAP7_75t_L g1750 ( 
.A(n_1555),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1616),
.B(n_1403),
.Y(n_1751)
);

A2O1A1Ixp33_ASAP7_75t_SL g1752 ( 
.A1(n_1533),
.A2(n_1450),
.B(n_1369),
.C(n_1394),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_L g1753 ( 
.A(n_1644),
.B(n_1645),
.C(n_1635),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1510),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1517),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1663),
.A2(n_1369),
.B1(n_1377),
.B2(n_1364),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1609),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1616),
.B(n_1358),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1653),
.A2(n_1343),
.B1(n_947),
.B2(n_29),
.Y(n_1759)
);

AND2x6_ASAP7_75t_L g1760 ( 
.A(n_1571),
.B(n_947),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1587),
.B(n_27),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1525),
.B(n_28),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1645),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1525),
.B(n_31),
.Y(n_1764)
);

A2O1A1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1630),
.A2(n_33),
.B(n_34),
.C(n_32),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1649),
.B(n_31),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1599),
.B(n_32),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1596),
.B(n_1515),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1520),
.B(n_1651),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1603),
.B(n_613),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1522),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1566),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1619),
.Y(n_1773)
);

BUFx2_ASAP7_75t_L g1774 ( 
.A(n_1600),
.Y(n_1774)
);

A2O1A1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1630),
.A2(n_37),
.B(n_38),
.C(n_36),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1619),
.B(n_35),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1545),
.Y(n_1777)
);

OR2x6_ASAP7_75t_L g1778 ( 
.A(n_1477),
.B(n_35),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1647),
.B(n_37),
.Y(n_1779)
);

INVx5_ASAP7_75t_L g1780 ( 
.A(n_1477),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1574),
.B(n_1477),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1548),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1625),
.B(n_39),
.Y(n_1783)
);

AND2x6_ASAP7_75t_SL g1784 ( 
.A(n_1598),
.B(n_40),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1634),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1648),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1618),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1625),
.B(n_42),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1633),
.B(n_43),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1504),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1506),
.B(n_44),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_SL g1792 ( 
.A(n_1658),
.B(n_1662),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1574),
.B(n_44),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1548),
.A2(n_48),
.B1(n_45),
.B2(n_47),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1505),
.Y(n_1795)
);

AO221x1_ASAP7_75t_L g1796 ( 
.A1(n_1620),
.A2(n_48),
.B1(n_45),
.B2(n_47),
.C(n_49),
.Y(n_1796)
);

INVx2_ASAP7_75t_SL g1797 ( 
.A(n_1487),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1613),
.B(n_50),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1613),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1633),
.B(n_1582),
.Y(n_1800)
);

HB1xp67_ASAP7_75t_L g1801 ( 
.A(n_1559),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1481),
.B(n_1646),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1637),
.Y(n_1803)
);

AOI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1629),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1620),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1523),
.B(n_55),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1642),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1528),
.B(n_1611),
.Y(n_1808)
);

OAI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1655),
.A2(n_64),
.B1(n_72),
.B2(n_56),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1565),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1511),
.B(n_610),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1576),
.B(n_56),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1629),
.B(n_611),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1507),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1593),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1639),
.A2(n_1578),
.B1(n_1605),
.B2(n_1577),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1532),
.B(n_612),
.Y(n_1817)
);

BUFx3_ASAP7_75t_L g1818 ( 
.A(n_1497),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1554),
.B(n_57),
.Y(n_1819)
);

BUFx2_ASAP7_75t_L g1820 ( 
.A(n_1626),
.Y(n_1820)
);

INVx4_ASAP7_75t_L g1821 ( 
.A(n_1657),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1661),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1822)
);

INVx5_ASAP7_75t_L g1823 ( 
.A(n_1489),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1532),
.B(n_1546),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1536),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1561),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1595),
.Y(n_1827)
);

NOR3xp33_ASAP7_75t_L g1828 ( 
.A(n_1533),
.B(n_1527),
.C(n_1624),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1568),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1608),
.B(n_58),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1552),
.A2(n_616),
.B(n_615),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1569),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1662),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1489),
.B(n_1562),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1575),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1567),
.Y(n_1836)
);

INVxp67_ASAP7_75t_L g1837 ( 
.A(n_1563),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1577),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1572),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1546),
.B(n_62),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1641),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1541),
.B(n_63),
.Y(n_1842)
);

INVx4_ASAP7_75t_L g1843 ( 
.A(n_1657),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1541),
.B(n_63),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1544),
.B(n_65),
.Y(n_1845)
);

NAND3xp33_ASAP7_75t_L g1846 ( 
.A(n_1660),
.B(n_65),
.C(n_66),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1661),
.A2(n_1643),
.B1(n_1636),
.B2(n_1573),
.C(n_1580),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1659),
.Y(n_1848)
);

XNOR2xp5_ASAP7_75t_L g1849 ( 
.A(n_1656),
.B(n_66),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1606),
.B(n_67),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1617),
.B(n_67),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1550),
.B(n_68),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1681),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1687),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1664),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1677),
.B(n_1621),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1691),
.Y(n_1857)
);

AND2x4_ASAP7_75t_L g1858 ( 
.A(n_1683),
.B(n_1780),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1695),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1673),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1772),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1700),
.Y(n_1862)
);

AO22x1_ASAP7_75t_L g1863 ( 
.A1(n_1680),
.A2(n_1617),
.B1(n_1475),
.B2(n_1654),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1708),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1839),
.Y(n_1865)
);

INVx2_ASAP7_75t_SL g1866 ( 
.A(n_1740),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1677),
.B(n_1623),
.Y(n_1867)
);

CKINVDCx6p67_ASAP7_75t_R g1868 ( 
.A(n_1818),
.Y(n_1868)
);

INVx4_ASAP7_75t_L g1869 ( 
.A(n_1673),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1786),
.B(n_1632),
.Y(n_1870)
);

AND2x6_ASAP7_75t_SL g1871 ( 
.A(n_1730),
.B(n_1601),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1711),
.Y(n_1872)
);

INVx5_ASAP7_75t_L g1873 ( 
.A(n_1723),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1665),
.B(n_1627),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1722),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1732),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1673),
.Y(n_1877)
);

BUFx6f_ASAP7_75t_L g1878 ( 
.A(n_1737),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1746),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1683),
.B(n_1588),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1665),
.B(n_1632),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1679),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1745),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1791),
.B(n_1494),
.Y(n_1884)
);

BUFx3_ASAP7_75t_L g1885 ( 
.A(n_1750),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1683),
.B(n_1780),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1672),
.B(n_1610),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1672),
.B(n_1612),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1684),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1748),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1754),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1755),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1678),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1686),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1771),
.Y(n_1895)
);

BUFx3_ASAP7_75t_L g1896 ( 
.A(n_1774),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1671),
.B(n_1577),
.Y(n_1897)
);

INVx3_ASAP7_75t_L g1898 ( 
.A(n_1746),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1725),
.A2(n_1580),
.B1(n_1552),
.B2(n_1652),
.Y(n_1899)
);

INVx4_ASAP7_75t_L g1900 ( 
.A(n_1741),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1851),
.B(n_1494),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_1737),
.Y(n_1902)
);

INVx2_ASAP7_75t_SL g1903 ( 
.A(n_1739),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1689),
.B(n_1494),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1685),
.B(n_1547),
.Y(n_1905)
);

INVx2_ASAP7_75t_SL g1906 ( 
.A(n_1797),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1703),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1713),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1773),
.B(n_1719),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1777),
.Y(n_1910)
);

INVx4_ASAP7_75t_L g1911 ( 
.A(n_1690),
.Y(n_1911)
);

BUFx2_ASAP7_75t_L g1912 ( 
.A(n_1731),
.Y(n_1912)
);

NOR2xp33_ASAP7_75t_L g1913 ( 
.A(n_1726),
.B(n_1547),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1709),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1812),
.B(n_1594),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1836),
.Y(n_1916)
);

BUFx3_ASAP7_75t_L g1917 ( 
.A(n_1820),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1719),
.B(n_1529),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1670),
.Y(n_1919)
);

NOR2xp67_ASAP7_75t_L g1920 ( 
.A(n_1690),
.B(n_1557),
.Y(n_1920)
);

BUFx4f_ASAP7_75t_L g1921 ( 
.A(n_1737),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1676),
.B(n_1529),
.Y(n_1922)
);

HAxp5_ASAP7_75t_L g1923 ( 
.A(n_1784),
.B(n_68),
.CON(n_1923),
.SN(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1787),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1803),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1728),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1717),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1676),
.B(n_1529),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1734),
.Y(n_1929)
);

INVx3_ASAP7_75t_L g1930 ( 
.A(n_1821),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1747),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1790),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1807),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1692),
.B(n_1601),
.Y(n_1934)
);

BUFx12f_ASAP7_75t_SL g1935 ( 
.A(n_1778),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1733),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1795),
.Y(n_1937)
);

INVx1_ASAP7_75t_SL g1938 ( 
.A(n_1696),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1814),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1825),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1826),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_1751),
.Y(n_1942)
);

NOR2xp67_ASAP7_75t_L g1943 ( 
.A(n_1735),
.B(n_1557),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1705),
.B(n_1508),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1815),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1837),
.B(n_1628),
.Y(n_1946)
);

OR2x6_ASAP7_75t_SL g1947 ( 
.A(n_1763),
.B(n_1475),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1829),
.Y(n_1948)
);

AOI22xp33_ASAP7_75t_L g1949 ( 
.A1(n_1796),
.A2(n_1529),
.B1(n_1475),
.B2(n_1588),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1827),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1780),
.Y(n_1951)
);

INVx5_ASAP7_75t_L g1952 ( 
.A(n_1723),
.Y(n_1952)
);

INVx2_ASAP7_75t_SL g1953 ( 
.A(n_1823),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_SL g1954 ( 
.A(n_1816),
.B(n_1591),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1725),
.B(n_1591),
.Y(n_1955)
);

AOI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1697),
.A2(n_1591),
.B1(n_1604),
.B2(n_1508),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1721),
.B(n_1468),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_R g1958 ( 
.A(n_1824),
.B(n_1531),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1674),
.B(n_1531),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1832),
.Y(n_1960)
);

HB1xp67_ASAP7_75t_L g1961 ( 
.A(n_1704),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1848),
.B(n_1468),
.Y(n_1962)
);

INVxp67_ASAP7_75t_L g1963 ( 
.A(n_1720),
.Y(n_1963)
);

HB1xp67_ASAP7_75t_L g1964 ( 
.A(n_1753),
.Y(n_1964)
);

CKINVDCx5p33_ASAP7_75t_R g1965 ( 
.A(n_1849),
.Y(n_1965)
);

OAI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1785),
.A2(n_1604),
.B1(n_1601),
.B2(n_1581),
.Y(n_1966)
);

NAND2x1p5_ASAP7_75t_L g1967 ( 
.A(n_1823),
.B(n_1571),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1693),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1715),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1710),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_1699),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1682),
.A2(n_1581),
.B1(n_1585),
.B2(n_1584),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1847),
.B(n_1792),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1835),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1753),
.B(n_1604),
.Y(n_1975)
);

BUFx6f_ASAP7_75t_L g1976 ( 
.A(n_1823),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1688),
.B(n_1584),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1841),
.Y(n_1978)
);

AOI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1701),
.A2(n_1585),
.B1(n_1589),
.B2(n_1586),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1768),
.Y(n_1980)
);

INVx2_ASAP7_75t_SL g1981 ( 
.A(n_1770),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1800),
.Y(n_1982)
);

BUFx2_ASAP7_75t_L g1983 ( 
.A(n_1802),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_SL g1984 ( 
.A(n_1778),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1767),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1694),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1668),
.B(n_1614),
.Y(n_1987)
);

BUFx6f_ASAP7_75t_L g1988 ( 
.A(n_1694),
.Y(n_1988)
);

CKINVDCx5p33_ASAP7_75t_R g1989 ( 
.A(n_1845),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1792),
.B(n_1589),
.Y(n_1990)
);

INVx3_ASAP7_75t_L g1991 ( 
.A(n_1821),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1817),
.B(n_1531),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1801),
.Y(n_1993)
);

INVxp33_ASAP7_75t_L g1994 ( 
.A(n_1729),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1707),
.B(n_1614),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1698),
.B(n_1560),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1810),
.Y(n_1997)
);

BUFx3_ASAP7_75t_L g1998 ( 
.A(n_1770),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1666),
.B(n_1586),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1842),
.B(n_1844),
.Y(n_2000)
);

BUFx2_ASAP7_75t_L g2001 ( 
.A(n_1843),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1762),
.B(n_1586),
.Y(n_2002)
);

BUFx6f_ASAP7_75t_L g2003 ( 
.A(n_1843),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1813),
.B(n_1560),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1762),
.B(n_1586),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1808),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1767),
.Y(n_2007)
);

AOI22xp33_ASAP7_75t_L g2008 ( 
.A1(n_1805),
.A2(n_1526),
.B1(n_1509),
.B2(n_1628),
.Y(n_2008)
);

INVx2_ASAP7_75t_SL g2009 ( 
.A(n_1778),
.Y(n_2009)
);

INVxp67_ASAP7_75t_L g2010 ( 
.A(n_1716),
.Y(n_2010)
);

NAND3xp33_ASAP7_75t_SL g2011 ( 
.A(n_1822),
.B(n_1490),
.C(n_1509),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1850),
.Y(n_2012)
);

HB1xp67_ASAP7_75t_L g2013 ( 
.A(n_1756),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_1756),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1850),
.Y(n_2015)
);

AND2x4_ASAP7_75t_L g2016 ( 
.A(n_1688),
.B(n_1560),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1761),
.Y(n_2017)
);

NAND2xp33_ASAP7_75t_L g2018 ( 
.A(n_1828),
.B(n_1628),
.Y(n_2018)
);

CKINVDCx20_ASAP7_75t_R g2019 ( 
.A(n_1769),
.Y(n_2019)
);

AOI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1811),
.A2(n_1526),
.B1(n_1631),
.B2(n_1562),
.Y(n_2020)
);

INVx4_ASAP7_75t_L g2021 ( 
.A(n_1706),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1702),
.B(n_1638),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1913),
.B(n_1667),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1853),
.Y(n_2024)
);

AOI21xp5_ASAP7_75t_L g2025 ( 
.A1(n_2013),
.A2(n_1766),
.B(n_1727),
.Y(n_2025)
);

NOR2x1_ASAP7_75t_L g2026 ( 
.A(n_2000),
.B(n_1781),
.Y(n_2026)
);

A2O1A1Ixp33_ASAP7_75t_L g2027 ( 
.A1(n_1973),
.A2(n_2000),
.B(n_1675),
.C(n_1804),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1961),
.B(n_1830),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_1989),
.B(n_1783),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_2010),
.B(n_1718),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1961),
.B(n_1764),
.Y(n_2031)
);

BUFx6f_ASAP7_75t_L g2032 ( 
.A(n_1951),
.Y(n_2032)
);

OR2x6_ASAP7_75t_L g2033 ( 
.A(n_1863),
.B(n_1758),
.Y(n_2033)
);

A2O1A1Ixp33_ASAP7_75t_L g2034 ( 
.A1(n_2013),
.A2(n_1759),
.B(n_1798),
.C(n_1840),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1959),
.B(n_1819),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_2010),
.B(n_1788),
.Y(n_2036)
);

NAND2x1p5_ASAP7_75t_L g2037 ( 
.A(n_1921),
.B(n_1562),
.Y(n_2037)
);

NOR2xp33_ASAP7_75t_L g2038 ( 
.A(n_1905),
.B(n_1789),
.Y(n_2038)
);

AOI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_2014),
.A2(n_1736),
.B(n_1742),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1884),
.B(n_1669),
.Y(n_2040)
);

AOI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_2014),
.A2(n_1742),
.B(n_1831),
.Y(n_2041)
);

AOI21xp5_ASAP7_75t_L g2042 ( 
.A1(n_1899),
.A2(n_1752),
.B(n_1846),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1854),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1865),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1855),
.Y(n_2045)
);

OAI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_1899),
.A2(n_1846),
.B(n_1794),
.Y(n_2046)
);

AOI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_1964),
.A2(n_1738),
.B(n_1724),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1971),
.B(n_1873),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1901),
.B(n_1712),
.Y(n_2049)
);

NOR2xp33_ASAP7_75t_SL g2050 ( 
.A(n_1935),
.B(n_1706),
.Y(n_2050)
);

BUFx8_ASAP7_75t_L g2051 ( 
.A(n_1984),
.Y(n_2051)
);

O2A1O1Ixp5_ASAP7_75t_L g2052 ( 
.A1(n_1955),
.A2(n_1794),
.B(n_1763),
.C(n_1775),
.Y(n_2052)
);

INVx3_ASAP7_75t_L g2053 ( 
.A(n_1885),
.Y(n_2053)
);

A2O1A1Ixp33_ASAP7_75t_L g2054 ( 
.A1(n_1949),
.A2(n_1765),
.B(n_1799),
.C(n_1838),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1857),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1881),
.A2(n_1714),
.B(n_1761),
.Y(n_2056)
);

INVx3_ASAP7_75t_L g2057 ( 
.A(n_1868),
.Y(n_2057)
);

OAI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_1947),
.A2(n_1782),
.B1(n_1809),
.B2(n_1776),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1951),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1859),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1881),
.A2(n_1749),
.B(n_1743),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1992),
.B(n_1852),
.Y(n_2062)
);

AOI21xp5_ASAP7_75t_L g2063 ( 
.A1(n_2002),
.A2(n_1806),
.B(n_1833),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1873),
.B(n_1833),
.Y(n_2064)
);

BUFx3_ASAP7_75t_L g2065 ( 
.A(n_1866),
.Y(n_2065)
);

NOR2xp33_ASAP7_75t_L g2066 ( 
.A(n_1900),
.B(n_1793),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_1900),
.B(n_1631),
.Y(n_2067)
);

AOI21xp5_ASAP7_75t_L g2068 ( 
.A1(n_2002),
.A2(n_2005),
.B(n_1995),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1861),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_2005),
.A2(n_1834),
.B(n_1779),
.Y(n_2070)
);

AOI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_1995),
.A2(n_1757),
.B(n_1744),
.Y(n_2071)
);

AOI22xp5_ASAP7_75t_L g2072 ( 
.A1(n_1984),
.A2(n_1723),
.B1(n_1757),
.B2(n_1744),
.Y(n_2072)
);

BUFx8_ASAP7_75t_L g2073 ( 
.A(n_1912),
.Y(n_2073)
);

O2A1O1Ixp33_ASAP7_75t_L g2074 ( 
.A1(n_1923),
.A2(n_2018),
.B(n_1966),
.C(n_2017),
.Y(n_2074)
);

O2A1O1Ixp33_ASAP7_75t_L g2075 ( 
.A1(n_1966),
.A2(n_1622),
.B(n_1490),
.C(n_71),
.Y(n_2075)
);

AOI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1874),
.A2(n_1638),
.B(n_1622),
.Y(n_2076)
);

AND2x2_ASAP7_75t_SL g2077 ( 
.A(n_1858),
.B(n_1526),
.Y(n_2077)
);

AOI21xp5_ASAP7_75t_L g2078 ( 
.A1(n_1874),
.A2(n_1760),
.B(n_1558),
.Y(n_2078)
);

AOI22xp5_ASAP7_75t_L g2079 ( 
.A1(n_1954),
.A2(n_1760),
.B1(n_1592),
.B2(n_1650),
.Y(n_2079)
);

BUFx5_ASAP7_75t_L g2080 ( 
.A(n_1858),
.Y(n_2080)
);

NOR2x1_ASAP7_75t_L g2081 ( 
.A(n_1998),
.B(n_1558),
.Y(n_2081)
);

OAI21x1_ASAP7_75t_L g2082 ( 
.A1(n_1999),
.A2(n_1975),
.B(n_1918),
.Y(n_2082)
);

CKINVDCx10_ASAP7_75t_R g2083 ( 
.A(n_1965),
.Y(n_2083)
);

BUFx2_ASAP7_75t_L g2084 ( 
.A(n_1917),
.Y(n_2084)
);

AOI21xp5_ASAP7_75t_L g2085 ( 
.A1(n_2022),
.A2(n_1558),
.B(n_1592),
.Y(n_2085)
);

AOI21xp5_ASAP7_75t_L g2086 ( 
.A1(n_2022),
.A2(n_1650),
.B(n_1592),
.Y(n_2086)
);

AOI21xp5_ASAP7_75t_L g2087 ( 
.A1(n_1990),
.A2(n_1650),
.B(n_71),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1978),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_1873),
.B(n_617),
.Y(n_2089)
);

AO21x1_ASAP7_75t_L g2090 ( 
.A1(n_1975),
.A2(n_69),
.B(n_70),
.Y(n_2090)
);

AOI21xp5_ASAP7_75t_L g2091 ( 
.A1(n_1909),
.A2(n_73),
.B(n_72),
.Y(n_2091)
);

OAI22xp5_ASAP7_75t_L g2092 ( 
.A1(n_1963),
.A2(n_1936),
.B1(n_1981),
.B2(n_2008),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1983),
.B(n_70),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_SL g2094 ( 
.A(n_1873),
.B(n_618),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_2006),
.B(n_74),
.Y(n_2095)
);

BUFx6f_ASAP7_75t_L g2096 ( 
.A(n_1951),
.Y(n_2096)
);

INVx2_ASAP7_75t_SL g2097 ( 
.A(n_1906),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1952),
.B(n_619),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1909),
.B(n_75),
.Y(n_2099)
);

OAI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_2012),
.A2(n_75),
.B(n_76),
.Y(n_2100)
);

NAND3xp33_ASAP7_75t_L g2101 ( 
.A(n_2015),
.B(n_77),
.C(n_78),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2004),
.B(n_79),
.Y(n_2102)
);

O2A1O1Ixp5_ASAP7_75t_L g2103 ( 
.A1(n_1922),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1938),
.B(n_80),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1882),
.Y(n_2105)
);

OAI22xp5_ASAP7_75t_L g2106 ( 
.A1(n_1963),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_SL g2107 ( 
.A(n_1952),
.B(n_621),
.Y(n_2107)
);

AOI21xp5_ASAP7_75t_L g2108 ( 
.A1(n_1952),
.A2(n_86),
.B(n_85),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_1908),
.B(n_608),
.Y(n_2109)
);

NOR2xp33_ASAP7_75t_L g2110 ( 
.A(n_1896),
.B(n_609),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1862),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1889),
.Y(n_2112)
);

AOI22xp5_ASAP7_75t_L g2113 ( 
.A1(n_2019),
.A2(n_2009),
.B1(n_1956),
.B2(n_2011),
.Y(n_2113)
);

NOR2xp33_ASAP7_75t_L g2114 ( 
.A(n_1994),
.B(n_609),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1938),
.B(n_84),
.Y(n_2115)
);

BUFx6f_ASAP7_75t_L g2116 ( 
.A(n_1976),
.Y(n_2116)
);

INVx6_ASAP7_75t_L g2117 ( 
.A(n_1869),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1864),
.Y(n_2118)
);

OAI22xp5_ASAP7_75t_L g2119 ( 
.A1(n_2008),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_1944),
.B(n_87),
.Y(n_2120)
);

BUFx8_ASAP7_75t_L g2121 ( 
.A(n_1915),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1894),
.Y(n_2122)
);

NAND2xp33_ASAP7_75t_L g2123 ( 
.A(n_1879),
.B(n_88),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1872),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1982),
.B(n_89),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1927),
.B(n_90),
.Y(n_2126)
);

AOI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_1952),
.A2(n_92),
.B(n_91),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_1993),
.B(n_90),
.Y(n_2128)
);

AOI21xp5_ASAP7_75t_L g2129 ( 
.A1(n_1887),
.A2(n_93),
.B(n_92),
.Y(n_2129)
);

HB1xp67_ASAP7_75t_L g2130 ( 
.A(n_1997),
.Y(n_2130)
);

AOI21xp5_ASAP7_75t_L g2131 ( 
.A1(n_1887),
.A2(n_94),
.B(n_93),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1907),
.Y(n_2132)
);

AOI21xp5_ASAP7_75t_L g2133 ( 
.A1(n_1888),
.A2(n_95),
.B(n_94),
.Y(n_2133)
);

INVx3_ASAP7_75t_L g2134 ( 
.A(n_1976),
.Y(n_2134)
);

INVx6_ASAP7_75t_L g2135 ( 
.A(n_1869),
.Y(n_2135)
);

O2A1O1Ixp33_ASAP7_75t_L g2136 ( 
.A1(n_1946),
.A2(n_96),
.B(n_91),
.C(n_95),
.Y(n_2136)
);

AO31x2_ASAP7_75t_L g2137 ( 
.A1(n_2041),
.A2(n_1922),
.A3(n_1928),
.B(n_1888),
.Y(n_2137)
);

OAI21x1_ASAP7_75t_L g2138 ( 
.A1(n_2085),
.A2(n_1999),
.B(n_1928),
.Y(n_2138)
);

AOI21xp5_ASAP7_75t_L g2139 ( 
.A1(n_2046),
.A2(n_2042),
.B(n_2039),
.Y(n_2139)
);

OAI21xp5_ASAP7_75t_L g2140 ( 
.A1(n_2034),
.A2(n_2011),
.B(n_1957),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2084),
.B(n_1875),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2044),
.Y(n_2142)
);

OAI21xp5_ASAP7_75t_L g2143 ( 
.A1(n_2052),
.A2(n_1957),
.B(n_1979),
.Y(n_2143)
);

BUFx3_ASAP7_75t_L g2144 ( 
.A(n_2065),
.Y(n_2144)
);

OAI21x1_ASAP7_75t_SL g2145 ( 
.A1(n_2100),
.A2(n_1911),
.B(n_1962),
.Y(n_2145)
);

NOR2xp33_ASAP7_75t_L g2146 ( 
.A(n_2053),
.B(n_1903),
.Y(n_2146)
);

NOR2x1_ASAP7_75t_SL g2147 ( 
.A(n_2033),
.B(n_1897),
.Y(n_2147)
);

AOI21xp5_ASAP7_75t_L g2148 ( 
.A1(n_2123),
.A2(n_1897),
.B(n_1962),
.Y(n_2148)
);

NOR2xp33_ASAP7_75t_L g2149 ( 
.A(n_2038),
.B(n_1911),
.Y(n_2149)
);

AOI21x1_ASAP7_75t_L g2150 ( 
.A1(n_2023),
.A2(n_2001),
.B(n_1985),
.Y(n_2150)
);

BUFx2_ASAP7_75t_L g2151 ( 
.A(n_2073),
.Y(n_2151)
);

AO31x2_ASAP7_75t_L g2152 ( 
.A1(n_2056),
.A2(n_2007),
.A3(n_1968),
.B(n_1924),
.Y(n_2152)
);

OAI21x1_ASAP7_75t_L g2153 ( 
.A1(n_2078),
.A2(n_1987),
.B(n_1972),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2130),
.Y(n_2154)
);

NAND3xp33_ASAP7_75t_L g2155 ( 
.A(n_2129),
.B(n_1970),
.C(n_1987),
.Y(n_2155)
);

O2A1O1Ixp5_ASAP7_75t_L g2156 ( 
.A1(n_2090),
.A2(n_2021),
.B(n_1930),
.C(n_1991),
.Y(n_2156)
);

A2O1A1Ixp33_ASAP7_75t_L g2157 ( 
.A1(n_2027),
.A2(n_2020),
.B(n_1919),
.C(n_1942),
.Y(n_2157)
);

OAI21xp5_ASAP7_75t_L g2158 ( 
.A1(n_2054),
.A2(n_1942),
.B(n_1934),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2024),
.Y(n_2159)
);

AO21x1_ASAP7_75t_L g2160 ( 
.A1(n_2030),
.A2(n_1883),
.B(n_1876),
.Y(n_2160)
);

OAI21xp5_ASAP7_75t_L g2161 ( 
.A1(n_2025),
.A2(n_1867),
.B(n_1856),
.Y(n_2161)
);

AOI21x1_ASAP7_75t_L g2162 ( 
.A1(n_2104),
.A2(n_1920),
.B(n_1916),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2068),
.B(n_1890),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2045),
.Y(n_2164)
);

BUFx3_ASAP7_75t_L g2165 ( 
.A(n_2073),
.Y(n_2165)
);

OAI21x1_ASAP7_75t_L g2166 ( 
.A1(n_2086),
.A2(n_1867),
.B(n_1856),
.Y(n_2166)
);

OAI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_2058),
.A2(n_1892),
.B1(n_1893),
.B2(n_1891),
.Y(n_2167)
);

OAI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_2101),
.A2(n_1996),
.B(n_1969),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2069),
.Y(n_2169)
);

OA21x2_ASAP7_75t_L g2170 ( 
.A1(n_2082),
.A2(n_1925),
.B(n_1910),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2031),
.B(n_1895),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2043),
.B(n_1933),
.Y(n_2172)
);

AND2x4_ASAP7_75t_L g2173 ( 
.A(n_2055),
.B(n_1945),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2088),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2062),
.B(n_1950),
.Y(n_2175)
);

AOI21xp33_ASAP7_75t_L g2176 ( 
.A1(n_2074),
.A2(n_1904),
.B(n_1870),
.Y(n_2176)
);

OAI21x1_ASAP7_75t_L g2177 ( 
.A1(n_2076),
.A2(n_1930),
.B(n_1991),
.Y(n_2177)
);

BUFx3_ASAP7_75t_L g2178 ( 
.A(n_2057),
.Y(n_2178)
);

OAI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_2103),
.A2(n_1921),
.B(n_1967),
.Y(n_2179)
);

A2O1A1Ixp33_ASAP7_75t_L g2180 ( 
.A1(n_2136),
.A2(n_1943),
.B(n_1980),
.C(n_1880),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2060),
.Y(n_2181)
);

OAI21xp5_ASAP7_75t_L g2182 ( 
.A1(n_2131),
.A2(n_1967),
.B(n_1953),
.Y(n_2182)
);

OAI22xp5_ASAP7_75t_L g2183 ( 
.A1(n_2099),
.A2(n_2021),
.B1(n_1898),
.B2(n_1879),
.Y(n_2183)
);

OAI21x1_ASAP7_75t_L g2184 ( 
.A1(n_2063),
.A2(n_1898),
.B(n_1877),
.Y(n_2184)
);

OAI21xp33_ASAP7_75t_L g2185 ( 
.A1(n_2114),
.A2(n_2003),
.B(n_1958),
.Y(n_2185)
);

OAI21xp5_ASAP7_75t_L g2186 ( 
.A1(n_2133),
.A2(n_2091),
.B(n_2075),
.Y(n_2186)
);

OAI21xp33_ASAP7_75t_L g2187 ( 
.A1(n_2106),
.A2(n_2003),
.B(n_2016),
.Y(n_2187)
);

OAI21x1_ASAP7_75t_L g2188 ( 
.A1(n_2071),
.A2(n_1877),
.B(n_1860),
.Y(n_2188)
);

OAI21x1_ASAP7_75t_L g2189 ( 
.A1(n_2070),
.A2(n_1860),
.B(n_1914),
.Y(n_2189)
);

OAI21xp5_ASAP7_75t_L g2190 ( 
.A1(n_2119),
.A2(n_2127),
.B(n_2108),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2111),
.B(n_1926),
.Y(n_2191)
);

OAI21x1_ASAP7_75t_L g2192 ( 
.A1(n_2061),
.A2(n_1931),
.B(n_1929),
.Y(n_2192)
);

AOI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_2064),
.A2(n_1886),
.B(n_1977),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2028),
.B(n_2003),
.Y(n_2194)
);

AND2x4_ASAP7_75t_L g2195 ( 
.A(n_2118),
.B(n_1886),
.Y(n_2195)
);

OAI21x1_ASAP7_75t_L g2196 ( 
.A1(n_2047),
.A2(n_1937),
.B(n_1932),
.Y(n_2196)
);

OAI21x1_ASAP7_75t_L g2197 ( 
.A1(n_2026),
.A2(n_1940),
.B(n_1939),
.Y(n_2197)
);

AOI21xp5_ASAP7_75t_L g2198 ( 
.A1(n_2089),
.A2(n_1977),
.B(n_2016),
.Y(n_2198)
);

AOI21xp5_ASAP7_75t_L g2199 ( 
.A1(n_2094),
.A2(n_1976),
.B(n_1880),
.Y(n_2199)
);

NAND3x1_ASAP7_75t_L g2200 ( 
.A(n_2036),
.B(n_1871),
.C(n_1878),
.Y(n_2200)
);

OA21x2_ASAP7_75t_L g2201 ( 
.A1(n_2113),
.A2(n_1960),
.B(n_1948),
.Y(n_2201)
);

AOI21xp5_ASAP7_75t_L g2202 ( 
.A1(n_2098),
.A2(n_1988),
.B(n_1986),
.Y(n_2202)
);

AOI21xp5_ASAP7_75t_L g2203 ( 
.A1(n_2107),
.A2(n_1988),
.B(n_1986),
.Y(n_2203)
);

CKINVDCx20_ASAP7_75t_R g2204 ( 
.A(n_2165),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2142),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_2149),
.B(n_2029),
.Y(n_2206)
);

OAI21x1_ASAP7_75t_L g2207 ( 
.A1(n_2150),
.A2(n_2092),
.B(n_2048),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2141),
.B(n_2035),
.Y(n_2208)
);

CKINVDCx11_ASAP7_75t_R g2209 ( 
.A(n_2151),
.Y(n_2209)
);

BUFx6f_ASAP7_75t_L g2210 ( 
.A(n_2178),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2172),
.Y(n_2211)
);

AO32x2_ASAP7_75t_L g2212 ( 
.A1(n_2167),
.A2(n_2097),
.A3(n_2124),
.B1(n_2112),
.B2(n_2122),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2164),
.Y(n_2213)
);

OAI21x1_ASAP7_75t_L g2214 ( 
.A1(n_2162),
.A2(n_2072),
.B(n_2081),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2172),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2169),
.Y(n_2216)
);

AOI21xp5_ASAP7_75t_L g2217 ( 
.A1(n_2139),
.A2(n_2077),
.B(n_2115),
.Y(n_2217)
);

OAI21x1_ASAP7_75t_SL g2218 ( 
.A1(n_2160),
.A2(n_2126),
.B(n_2095),
.Y(n_2218)
);

AOI21xp5_ASAP7_75t_L g2219 ( 
.A1(n_2140),
.A2(n_2087),
.B(n_2125),
.Y(n_2219)
);

O2A1O1Ixp33_ASAP7_75t_L g2220 ( 
.A1(n_2186),
.A2(n_2093),
.B(n_2110),
.C(n_2109),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2154),
.B(n_2102),
.Y(n_2221)
);

AOI21xp5_ASAP7_75t_L g2222 ( 
.A1(n_2140),
.A2(n_2033),
.B(n_2079),
.Y(n_2222)
);

OR2x2_ASAP7_75t_L g2223 ( 
.A(n_2171),
.B(n_2128),
.Y(n_2223)
);

HB1xp67_ASAP7_75t_L g2224 ( 
.A(n_2163),
.Y(n_2224)
);

AOI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_2167),
.A2(n_2050),
.B1(n_2049),
.B2(n_2066),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2159),
.Y(n_2226)
);

OAI21x1_ASAP7_75t_L g2227 ( 
.A1(n_2177),
.A2(n_2134),
.B(n_2132),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2174),
.Y(n_2228)
);

NOR2xp33_ASAP7_75t_SL g2229 ( 
.A(n_2185),
.B(n_2080),
.Y(n_2229)
);

INVx6_ASAP7_75t_L g2230 ( 
.A(n_2144),
.Y(n_2230)
);

AO31x2_ASAP7_75t_L g2231 ( 
.A1(n_2147),
.A2(n_2105),
.A3(n_1974),
.B(n_1941),
.Y(n_2231)
);

A2O1A1Ixp33_ASAP7_75t_L g2232 ( 
.A1(n_2186),
.A2(n_2040),
.B(n_2120),
.C(n_2067),
.Y(n_2232)
);

AOI21xp33_ASAP7_75t_L g2233 ( 
.A1(n_2155),
.A2(n_2121),
.B(n_2134),
.Y(n_2233)
);

AO21x1_ASAP7_75t_L g2234 ( 
.A1(n_2163),
.A2(n_2037),
.B(n_2121),
.Y(n_2234)
);

INVx3_ASAP7_75t_L g2235 ( 
.A(n_2195),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2181),
.Y(n_2236)
);

AOI21x1_ASAP7_75t_L g2237 ( 
.A1(n_2183),
.A2(n_2203),
.B(n_2202),
.Y(n_2237)
);

A2O1A1Ixp33_ASAP7_75t_L g2238 ( 
.A1(n_2158),
.A2(n_2059),
.B(n_2096),
.C(n_2032),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2137),
.B(n_2080),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2173),
.Y(n_2240)
);

NOR2xp67_ASAP7_75t_SL g2241 ( 
.A(n_2199),
.B(n_2117),
.Y(n_2241)
);

A2O1A1Ixp33_ASAP7_75t_L g2242 ( 
.A1(n_2158),
.A2(n_2059),
.B(n_2096),
.C(n_2032),
.Y(n_2242)
);

OR2x2_ASAP7_75t_L g2243 ( 
.A(n_2171),
.B(n_2032),
.Y(n_2243)
);

OAI21xp5_ASAP7_75t_L g2244 ( 
.A1(n_2168),
.A2(n_96),
.B(n_97),
.Y(n_2244)
);

NAND3xp33_ASAP7_75t_L g2245 ( 
.A(n_2168),
.B(n_2051),
.C(n_2059),
.Y(n_2245)
);

AO31x2_ASAP7_75t_L g2246 ( 
.A1(n_2148),
.A2(n_2080),
.A3(n_2116),
.B(n_2096),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2173),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2137),
.B(n_2080),
.Y(n_2248)
);

OAI21x1_ASAP7_75t_L g2249 ( 
.A1(n_2237),
.A2(n_2138),
.B(n_2166),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_2212),
.Y(n_2250)
);

BUFx12f_ASAP7_75t_L g2251 ( 
.A(n_2209),
.Y(n_2251)
);

NOR2xp33_ASAP7_75t_L g2252 ( 
.A(n_2206),
.B(n_2146),
.Y(n_2252)
);

OAI21x1_ASAP7_75t_L g2253 ( 
.A1(n_2207),
.A2(n_2248),
.B(n_2239),
.Y(n_2253)
);

OA21x2_ASAP7_75t_L g2254 ( 
.A1(n_2239),
.A2(n_2184),
.B(n_2161),
.Y(n_2254)
);

INVx2_ASAP7_75t_SL g2255 ( 
.A(n_2230),
.Y(n_2255)
);

INVx4_ASAP7_75t_L g2256 ( 
.A(n_2210),
.Y(n_2256)
);

OAI221xp5_ASAP7_75t_SL g2257 ( 
.A1(n_2219),
.A2(n_2157),
.B1(n_2187),
.B2(n_2180),
.C(n_2194),
.Y(n_2257)
);

CKINVDCx11_ASAP7_75t_R g2258 ( 
.A(n_2204),
.Y(n_2258)
);

OAI21xp5_ASAP7_75t_L g2259 ( 
.A1(n_2244),
.A2(n_2200),
.B(n_2190),
.Y(n_2259)
);

NOR2x1_ASAP7_75t_SL g2260 ( 
.A(n_2245),
.B(n_2183),
.Y(n_2260)
);

OAI21xp5_ASAP7_75t_L g2261 ( 
.A1(n_2244),
.A2(n_2190),
.B(n_2143),
.Y(n_2261)
);

OA21x2_ASAP7_75t_L g2262 ( 
.A1(n_2248),
.A2(n_2161),
.B(n_2189),
.Y(n_2262)
);

NOR2xp67_ASAP7_75t_R g2263 ( 
.A(n_2230),
.B(n_2117),
.Y(n_2263)
);

OAI21x1_ASAP7_75t_L g2264 ( 
.A1(n_2222),
.A2(n_2153),
.B(n_2192),
.Y(n_2264)
);

NOR2xp33_ASAP7_75t_L g2265 ( 
.A(n_2210),
.B(n_2135),
.Y(n_2265)
);

OAI21x1_ASAP7_75t_L g2266 ( 
.A1(n_2222),
.A2(n_2188),
.B(n_2196),
.Y(n_2266)
);

OA21x2_ASAP7_75t_L g2267 ( 
.A1(n_2227),
.A2(n_2197),
.B(n_2176),
.Y(n_2267)
);

OAI22xp5_ASAP7_75t_L g2268 ( 
.A1(n_2225),
.A2(n_2143),
.B1(n_2182),
.B2(n_2175),
.Y(n_2268)
);

HB1xp67_ASAP7_75t_L g2269 ( 
.A(n_2224),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2226),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2236),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2211),
.B(n_2152),
.Y(n_2272)
);

AOI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_2219),
.A2(n_2182),
.B(n_2198),
.Y(n_2273)
);

INVx3_ASAP7_75t_L g2274 ( 
.A(n_2246),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2269),
.B(n_2215),
.Y(n_2275)
);

NAND2x1p5_ASAP7_75t_L g2276 ( 
.A(n_2256),
.B(n_2241),
.Y(n_2276)
);

OAI21x1_ASAP7_75t_L g2277 ( 
.A1(n_2274),
.A2(n_2253),
.B(n_2249),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2250),
.Y(n_2278)
);

INVx4_ASAP7_75t_L g2279 ( 
.A(n_2251),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2270),
.B(n_2223),
.Y(n_2280)
);

AO21x2_ASAP7_75t_L g2281 ( 
.A1(n_2250),
.A2(n_2218),
.B(n_2217),
.Y(n_2281)
);

OAI21x1_ASAP7_75t_L g2282 ( 
.A1(n_2274),
.A2(n_2214),
.B(n_2235),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2270),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2273),
.B(n_2208),
.Y(n_2284)
);

OAI21xp5_ASAP7_75t_SL g2285 ( 
.A1(n_2276),
.A2(n_2261),
.B(n_2259),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2280),
.Y(n_2286)
);

OAI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_2284),
.A2(n_2261),
.B1(n_2259),
.B2(n_2268),
.Y(n_2287)
);

CKINVDCx20_ASAP7_75t_R g2288 ( 
.A(n_2279),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2278),
.Y(n_2289)
);

AOI22xp33_ASAP7_75t_L g2290 ( 
.A1(n_2281),
.A2(n_2268),
.B1(n_2250),
.B2(n_2245),
.Y(n_2290)
);

BUFx2_ASAP7_75t_L g2291 ( 
.A(n_2279),
.Y(n_2291)
);

OAI22x1_ASAP7_75t_L g2292 ( 
.A1(n_2279),
.A2(n_2255),
.B1(n_2252),
.B2(n_2256),
.Y(n_2292)
);

OA21x2_ASAP7_75t_L g2293 ( 
.A1(n_2285),
.A2(n_2277),
.B(n_2282),
.Y(n_2293)
);

OA21x2_ASAP7_75t_L g2294 ( 
.A1(n_2290),
.A2(n_2277),
.B(n_2282),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2289),
.Y(n_2295)
);

BUFx2_ASAP7_75t_L g2296 ( 
.A(n_2288),
.Y(n_2296)
);

HB1xp67_ASAP7_75t_L g2297 ( 
.A(n_2287),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2289),
.Y(n_2298)
);

INVxp67_ASAP7_75t_R g2299 ( 
.A(n_2292),
.Y(n_2299)
);

INVxp33_ASAP7_75t_L g2300 ( 
.A(n_2291),
.Y(n_2300)
);

AO21x2_ASAP7_75t_L g2301 ( 
.A1(n_2286),
.A2(n_2278),
.B(n_2281),
.Y(n_2301)
);

AOI22xp33_ASAP7_75t_L g2302 ( 
.A1(n_2290),
.A2(n_2281),
.B1(n_2262),
.B2(n_2254),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2297),
.B(n_2283),
.Y(n_2303)
);

OR2x2_ASAP7_75t_L g2304 ( 
.A(n_2297),
.B(n_2280),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2299),
.B(n_2251),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2295),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_2299),
.B(n_2251),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2295),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2299),
.B(n_2296),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2296),
.B(n_2258),
.Y(n_2310)
);

INVx4_ASAP7_75t_SL g2311 ( 
.A(n_2300),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2298),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2301),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2310),
.B(n_2300),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_2305),
.B(n_2256),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2305),
.B(n_2256),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2306),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2311),
.Y(n_2318)
);

HB1xp67_ASAP7_75t_L g2319 ( 
.A(n_2311),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2307),
.B(n_2255),
.Y(n_2320)
);

INVx3_ASAP7_75t_L g2321 ( 
.A(n_2309),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_L g2322 ( 
.A(n_2307),
.B(n_2083),
.Y(n_2322)
);

INVx2_ASAP7_75t_SL g2323 ( 
.A(n_2314),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2321),
.B(n_2309),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2322),
.B(n_2311),
.Y(n_2325)
);

HB1xp67_ASAP7_75t_L g2326 ( 
.A(n_2321),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2326),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2326),
.Y(n_2328)
);

AOI22xp33_ASAP7_75t_L g2329 ( 
.A1(n_2324),
.A2(n_2321),
.B1(n_2313),
.B2(n_2302),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2325),
.B(n_2322),
.Y(n_2330)
);

NOR2x1p5_ASAP7_75t_L g2331 ( 
.A(n_2330),
.B(n_2318),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2329),
.B(n_2323),
.Y(n_2332)
);

OR2x2_ASAP7_75t_L g2333 ( 
.A(n_2327),
.B(n_2304),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2329),
.B(n_2319),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2328),
.B(n_2320),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2327),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2333),
.Y(n_2337)
);

NAND4xp25_ASAP7_75t_L g2338 ( 
.A(n_2332),
.B(n_2318),
.C(n_2317),
.D(n_2315),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_2335),
.B(n_2319),
.Y(n_2339)
);

OAI21xp5_ASAP7_75t_L g2340 ( 
.A1(n_2334),
.A2(n_2303),
.B(n_2302),
.Y(n_2340)
);

AND2x4_ASAP7_75t_L g2341 ( 
.A(n_2331),
.B(n_2336),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2331),
.B(n_2316),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2331),
.B(n_2308),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2331),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2333),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2331),
.Y(n_2346)
);

OR2x2_ASAP7_75t_L g2347 ( 
.A(n_2337),
.B(n_2345),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2341),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2342),
.B(n_2312),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2341),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2343),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2339),
.B(n_2301),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2344),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2346),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2338),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2340),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2341),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2342),
.B(n_2293),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2341),
.Y(n_2359)
);

OR2x2_ASAP7_75t_L g2360 ( 
.A(n_2347),
.B(n_2301),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2356),
.B(n_2301),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_2348),
.B(n_2293),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_2350),
.B(n_2293),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2349),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2357),
.Y(n_2365)
);

INVx3_ASAP7_75t_L g2366 ( 
.A(n_2359),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2356),
.Y(n_2367)
);

NOR2xp33_ASAP7_75t_L g2368 ( 
.A(n_2353),
.B(n_2354),
.Y(n_2368)
);

OR2x2_ASAP7_75t_L g2369 ( 
.A(n_2355),
.B(n_2301),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2352),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2358),
.B(n_2294),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2351),
.B(n_2294),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2352),
.B(n_2294),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2348),
.B(n_2293),
.Y(n_2374)
);

AOI22xp5_ASAP7_75t_L g2375 ( 
.A1(n_2362),
.A2(n_2313),
.B1(n_2294),
.B2(n_2293),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2366),
.Y(n_2376)
);

INVx2_ASAP7_75t_SL g2377 ( 
.A(n_2366),
.Y(n_2377)
);

OAI221xp5_ASAP7_75t_L g2378 ( 
.A1(n_2371),
.A2(n_2294),
.B1(n_2298),
.B2(n_2220),
.C(n_2276),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2368),
.B(n_2283),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2364),
.B(n_2210),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2365),
.B(n_2253),
.Y(n_2381)
);

AND2x4_ASAP7_75t_SL g2382 ( 
.A(n_2374),
.B(n_2265),
.Y(n_2382)
);

OAI21xp33_ASAP7_75t_L g2383 ( 
.A1(n_2363),
.A2(n_2276),
.B(n_2275),
.Y(n_2383)
);

INVx2_ASAP7_75t_SL g2384 ( 
.A(n_2360),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2367),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2367),
.Y(n_2386)
);

AOI21xp33_ASAP7_75t_L g2387 ( 
.A1(n_2372),
.A2(n_2051),
.B(n_2274),
.Y(n_2387)
);

AOI22xp5_ASAP7_75t_L g2388 ( 
.A1(n_2373),
.A2(n_2234),
.B1(n_2221),
.B2(n_2233),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2386),
.Y(n_2389)
);

NAND2x1_ASAP7_75t_L g2390 ( 
.A(n_2376),
.B(n_2369),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_2377),
.B(n_2370),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2385),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2379),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_L g2394 ( 
.A(n_2382),
.B(n_2361),
.Y(n_2394)
);

AOI221xp5_ASAP7_75t_L g2395 ( 
.A1(n_2387),
.A2(n_2233),
.B1(n_2257),
.B2(n_2274),
.C(n_2271),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2380),
.B(n_2249),
.Y(n_2396)
);

O2A1O1Ixp33_ASAP7_75t_L g2397 ( 
.A1(n_2384),
.A2(n_2232),
.B(n_99),
.C(n_97),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2383),
.B(n_2381),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2378),
.Y(n_2399)
);

O2A1O1Ixp5_ASAP7_75t_L g2400 ( 
.A1(n_2375),
.A2(n_2388),
.B(n_2271),
.C(n_2156),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2376),
.B(n_2260),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2386),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2386),
.Y(n_2403)
);

AOI221xp5_ASAP7_75t_L g2404 ( 
.A1(n_2387),
.A2(n_2272),
.B1(n_2179),
.B2(n_2145),
.C(n_2176),
.Y(n_2404)
);

OAI21xp5_ASAP7_75t_L g2405 ( 
.A1(n_2377),
.A2(n_2179),
.B(n_2266),
.Y(n_2405)
);

AOI22xp33_ASAP7_75t_L g2406 ( 
.A1(n_2386),
.A2(n_2267),
.B1(n_2262),
.B2(n_2254),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2386),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2376),
.B(n_2260),
.Y(n_2408)
);

OAI21xp5_ASAP7_75t_L g2409 ( 
.A1(n_2377),
.A2(n_2266),
.B(n_2264),
.Y(n_2409)
);

AOI22xp33_ASAP7_75t_L g2410 ( 
.A1(n_2386),
.A2(n_2267),
.B1(n_2262),
.B2(n_2254),
.Y(n_2410)
);

OR2x2_ASAP7_75t_L g2411 ( 
.A(n_2389),
.B(n_2254),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2402),
.B(n_2262),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2403),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2407),
.Y(n_2414)
);

NOR2xp33_ASAP7_75t_L g2415 ( 
.A(n_2392),
.B(n_98),
.Y(n_2415)
);

OAI21xp33_ASAP7_75t_L g2416 ( 
.A1(n_2401),
.A2(n_2247),
.B(n_2240),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2391),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2408),
.B(n_2267),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2390),
.Y(n_2419)
);

AOI211xp5_ASAP7_75t_L g2420 ( 
.A1(n_2398),
.A2(n_100),
.B(n_101),
.C(n_99),
.Y(n_2420)
);

INVxp67_ASAP7_75t_L g2421 ( 
.A(n_2394),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_2393),
.Y(n_2422)
);

AOI322xp5_ASAP7_75t_L g2423 ( 
.A1(n_2399),
.A2(n_2238),
.A3(n_2242),
.B1(n_2229),
.B2(n_2272),
.C1(n_2263),
.C2(n_2212),
.Y(n_2423)
);

OR2x2_ASAP7_75t_L g2424 ( 
.A(n_2396),
.B(n_98),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2400),
.Y(n_2425)
);

CKINVDCx20_ASAP7_75t_R g2426 ( 
.A(n_2409),
.Y(n_2426)
);

INVx1_ASAP7_75t_SL g2427 ( 
.A(n_2405),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2397),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_SL g2429 ( 
.A(n_2395),
.B(n_1878),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2404),
.B(n_2410),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2406),
.B(n_2267),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2405),
.Y(n_2432)
);

OAI21xp5_ASAP7_75t_L g2433 ( 
.A1(n_2389),
.A2(n_2264),
.B(n_2229),
.Y(n_2433)
);

AO32x1_ASAP7_75t_L g2434 ( 
.A1(n_2389),
.A2(n_2263),
.A3(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_2434)
);

AOI21xp33_ASAP7_75t_L g2435 ( 
.A1(n_2394),
.A2(n_103),
.B(n_104),
.Y(n_2435)
);

NAND3xp33_ASAP7_75t_L g2436 ( 
.A(n_2394),
.B(n_1902),
.C(n_1878),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2389),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2389),
.Y(n_2438)
);

OAI22xp5_ASAP7_75t_L g2439 ( 
.A1(n_2392),
.A2(n_2135),
.B1(n_1902),
.B2(n_2243),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_2401),
.B(n_2235),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2389),
.Y(n_2441)
);

XNOR2x1_ASAP7_75t_L g2442 ( 
.A(n_2391),
.B(n_103),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_2389),
.B(n_104),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2401),
.B(n_2246),
.Y(n_2444)
);

NOR2x1_ASAP7_75t_L g2445 ( 
.A(n_2389),
.B(n_105),
.Y(n_2445)
);

INVxp67_ASAP7_75t_L g2446 ( 
.A(n_2389),
.Y(n_2446)
);

OR2x2_ASAP7_75t_L g2447 ( 
.A(n_2389),
.B(n_105),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2445),
.B(n_2419),
.Y(n_2448)
);

AOI22xp5_ASAP7_75t_L g2449 ( 
.A1(n_2426),
.A2(n_1902),
.B1(n_2201),
.B2(n_2116),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2417),
.B(n_106),
.Y(n_2450)
);

AO21x1_ASAP7_75t_L g2451 ( 
.A1(n_2413),
.A2(n_114),
.B(n_106),
.Y(n_2451)
);

AOI221xp5_ASAP7_75t_L g2452 ( 
.A1(n_2446),
.A2(n_2427),
.B1(n_2432),
.B2(n_2437),
.C(n_2414),
.Y(n_2452)
);

AOI22xp5_ASAP7_75t_L g2453 ( 
.A1(n_2425),
.A2(n_2201),
.B1(n_2116),
.B2(n_2195),
.Y(n_2453)
);

AOI22xp5_ASAP7_75t_L g2454 ( 
.A1(n_2438),
.A2(n_2170),
.B1(n_2191),
.B2(n_2205),
.Y(n_2454)
);

OAI21xp33_ASAP7_75t_L g2455 ( 
.A1(n_2442),
.A2(n_2193),
.B(n_107),
.Y(n_2455)
);

OAI21xp5_ASAP7_75t_L g2456 ( 
.A1(n_2441),
.A2(n_2191),
.B(n_108),
.Y(n_2456)
);

NOR2xp33_ASAP7_75t_L g2457 ( 
.A(n_2447),
.B(n_109),
.Y(n_2457)
);

AND2x2_ASAP7_75t_L g2458 ( 
.A(n_2422),
.B(n_2246),
.Y(n_2458)
);

AOI22xp5_ASAP7_75t_L g2459 ( 
.A1(n_2428),
.A2(n_2170),
.B1(n_2216),
.B2(n_2213),
.Y(n_2459)
);

XOR2x2_ASAP7_75t_L g2460 ( 
.A(n_2420),
.B(n_110),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2440),
.B(n_2421),
.Y(n_2461)
);

AOI21xp5_ASAP7_75t_L g2462 ( 
.A1(n_2435),
.A2(n_110),
.B(n_111),
.Y(n_2462)
);

O2A1O1Ixp33_ASAP7_75t_L g2463 ( 
.A1(n_2443),
.A2(n_114),
.B(n_112),
.C(n_113),
.Y(n_2463)
);

NOR2xp67_ASAP7_75t_L g2464 ( 
.A(n_2415),
.B(n_112),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_SL g2465 ( 
.A(n_2412),
.B(n_113),
.Y(n_2465)
);

OAI22xp5_ASAP7_75t_L g2466 ( 
.A1(n_2430),
.A2(n_2228),
.B1(n_1988),
.B2(n_1986),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2434),
.Y(n_2467)
);

AOI211xp5_ASAP7_75t_L g2468 ( 
.A1(n_2424),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_2468)
);

OAI22xp33_ASAP7_75t_L g2469 ( 
.A1(n_2411),
.A2(n_2212),
.B1(n_118),
.B2(n_115),
.Y(n_2469)
);

NAND4xp25_ASAP7_75t_L g2470 ( 
.A(n_2436),
.B(n_119),
.C(n_116),
.D(n_118),
.Y(n_2470)
);

O2A1O1Ixp33_ASAP7_75t_SL g2471 ( 
.A1(n_2429),
.A2(n_122),
.B(n_120),
.C(n_121),
.Y(n_2471)
);

AOI221xp5_ASAP7_75t_L g2472 ( 
.A1(n_2418),
.A2(n_123),
.B1(n_120),
.B2(n_121),
.C(n_124),
.Y(n_2472)
);

OAI22xp5_ASAP7_75t_L g2473 ( 
.A1(n_2431),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_2473)
);

AOI221xp5_ASAP7_75t_L g2474 ( 
.A1(n_2444),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.C(n_128),
.Y(n_2474)
);

AOI21xp5_ASAP7_75t_L g2475 ( 
.A1(n_2434),
.A2(n_2439),
.B(n_2416),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2433),
.Y(n_2476)
);

AOI21xp5_ASAP7_75t_L g2477 ( 
.A1(n_2423),
.A2(n_127),
.B(n_128),
.Y(n_2477)
);

OAI21xp33_ASAP7_75t_L g2478 ( 
.A1(n_2417),
.A2(n_129),
.B(n_130),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2442),
.Y(n_2479)
);

BUFx4f_ASAP7_75t_SL g2480 ( 
.A(n_2417),
.Y(n_2480)
);

AO21x1_ASAP7_75t_L g2481 ( 
.A1(n_2417),
.A2(n_139),
.B(n_131),
.Y(n_2481)
);

HB1xp67_ASAP7_75t_L g2482 ( 
.A(n_2445),
.Y(n_2482)
);

NOR4xp25_ASAP7_75t_L g2483 ( 
.A(n_2419),
.B(n_133),
.C(n_131),
.D(n_132),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2445),
.Y(n_2484)
);

OAI22xp5_ASAP7_75t_L g2485 ( 
.A1(n_2417),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2467),
.B(n_134),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2461),
.B(n_135),
.Y(n_2487)
);

AOI22xp5_ASAP7_75t_L g2488 ( 
.A1(n_2452),
.A2(n_2080),
.B1(n_138),
.B2(n_136),
.Y(n_2488)
);

NOR2xp33_ASAP7_75t_L g2489 ( 
.A(n_2482),
.B(n_137),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2483),
.B(n_136),
.Y(n_2490)
);

OAI22xp5_ASAP7_75t_L g2491 ( 
.A1(n_2480),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_2491)
);

AOI221xp5_ASAP7_75t_L g2492 ( 
.A1(n_2473),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.C(n_144),
.Y(n_2492)
);

OAI21xp33_ASAP7_75t_SL g2493 ( 
.A1(n_2448),
.A2(n_144),
.B(n_143),
.Y(n_2493)
);

AOI221x1_ASAP7_75t_L g2494 ( 
.A1(n_2484),
.A2(n_146),
.B1(n_142),
.B2(n_145),
.C(n_148),
.Y(n_2494)
);

OAI221xp5_ASAP7_75t_L g2495 ( 
.A1(n_2478),
.A2(n_148),
.B1(n_145),
.B2(n_146),
.C(n_149),
.Y(n_2495)
);

OAI221xp5_ASAP7_75t_L g2496 ( 
.A1(n_2472),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.C(n_153),
.Y(n_2496)
);

AOI222xp33_ASAP7_75t_L g2497 ( 
.A1(n_2464),
.A2(n_152),
.B1(n_154),
.B2(n_150),
.C1(n_151),
.C2(n_153),
.Y(n_2497)
);

OAI21xp5_ASAP7_75t_SL g2498 ( 
.A1(n_2470),
.A2(n_154),
.B(n_155),
.Y(n_2498)
);

NAND2x1_ASAP7_75t_L g2499 ( 
.A(n_2450),
.B(n_156),
.Y(n_2499)
);

AOI211xp5_ASAP7_75t_L g2500 ( 
.A1(n_2481),
.A2(n_2451),
.B(n_2471),
.C(n_2474),
.Y(n_2500)
);

OAI21xp33_ASAP7_75t_SL g2501 ( 
.A1(n_2465),
.A2(n_156),
.B(n_157),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2457),
.Y(n_2502)
);

AOI221xp5_ASAP7_75t_L g2503 ( 
.A1(n_2475),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.C(n_161),
.Y(n_2503)
);

NOR4xp75_ASAP7_75t_L g2504 ( 
.A(n_2456),
.B(n_162),
.C(n_158),
.D(n_159),
.Y(n_2504)
);

OAI22xp5_ASAP7_75t_L g2505 ( 
.A1(n_2476),
.A2(n_2468),
.B1(n_2479),
.B2(n_2477),
.Y(n_2505)
);

AOI21xp33_ASAP7_75t_L g2506 ( 
.A1(n_2463),
.A2(n_162),
.B(n_163),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2458),
.B(n_164),
.Y(n_2507)
);

AOI221xp5_ASAP7_75t_L g2508 ( 
.A1(n_2455),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.C(n_168),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2460),
.Y(n_2509)
);

AOI21xp33_ASAP7_75t_L g2510 ( 
.A1(n_2462),
.A2(n_165),
.B(n_166),
.Y(n_2510)
);

AOI21xp5_ASAP7_75t_L g2511 ( 
.A1(n_2485),
.A2(n_167),
.B(n_168),
.Y(n_2511)
);

OAI322xp33_ASAP7_75t_L g2512 ( 
.A1(n_2466),
.A2(n_177),
.A3(n_176),
.B1(n_174),
.B2(n_169),
.C1(n_173),
.C2(n_175),
.Y(n_2512)
);

AOI211xp5_ASAP7_75t_L g2513 ( 
.A1(n_2469),
.A2(n_174),
.B(n_169),
.C(n_173),
.Y(n_2513)
);

OAI22xp5_ASAP7_75t_L g2514 ( 
.A1(n_2459),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_2514)
);

AOI211xp5_ASAP7_75t_L g2515 ( 
.A1(n_2454),
.A2(n_180),
.B(n_178),
.C(n_179),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2453),
.B(n_178),
.Y(n_2516)
);

AOI21xp5_ASAP7_75t_L g2517 ( 
.A1(n_2449),
.A2(n_180),
.B(n_181),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2467),
.B(n_181),
.Y(n_2518)
);

AOI221x1_ASAP7_75t_L g2519 ( 
.A1(n_2467),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.C(n_185),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2467),
.B(n_182),
.Y(n_2520)
);

NAND4xp25_ASAP7_75t_L g2521 ( 
.A(n_2452),
.B(n_185),
.C(n_183),
.D(n_184),
.Y(n_2521)
);

OAI21xp33_ASAP7_75t_L g2522 ( 
.A1(n_2452),
.A2(n_186),
.B(n_187),
.Y(n_2522)
);

AOI21xp5_ASAP7_75t_L g2523 ( 
.A1(n_2467),
.A2(n_186),
.B(n_187),
.Y(n_2523)
);

AOI21xp5_ASAP7_75t_L g2524 ( 
.A1(n_2467),
.A2(n_188),
.B(n_189),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2467),
.B(n_188),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2467),
.B(n_189),
.Y(n_2526)
);

O2A1O1Ixp5_ASAP7_75t_SL g2527 ( 
.A1(n_2467),
.A2(n_192),
.B(n_190),
.C(n_191),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2467),
.B(n_191),
.Y(n_2528)
);

NOR3xp33_ASAP7_75t_L g2529 ( 
.A(n_2452),
.B(n_192),
.C(n_193),
.Y(n_2529)
);

NOR2xp33_ASAP7_75t_R g2530 ( 
.A(n_2480),
.B(n_195),
.Y(n_2530)
);

AOI211xp5_ASAP7_75t_L g2531 ( 
.A1(n_2467),
.A2(n_197),
.B(n_195),
.C(n_196),
.Y(n_2531)
);

OAI22xp5_ASAP7_75t_L g2532 ( 
.A1(n_2480),
.A2(n_199),
.B1(n_196),
.B2(n_198),
.Y(n_2532)
);

AOI21x1_ASAP7_75t_L g2533 ( 
.A1(n_2448),
.A2(n_198),
.B(n_199),
.Y(n_2533)
);

AOI221x1_ASAP7_75t_L g2534 ( 
.A1(n_2467),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.C(n_203),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2467),
.B(n_200),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2481),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2467),
.B(n_201),
.Y(n_2537)
);

AOI21xp33_ASAP7_75t_L g2538 ( 
.A1(n_2448),
.A2(n_202),
.B(n_203),
.Y(n_2538)
);

AOI21xp33_ASAP7_75t_L g2539 ( 
.A1(n_2448),
.A2(n_204),
.B(n_205),
.Y(n_2539)
);

AOI22xp33_ASAP7_75t_L g2540 ( 
.A1(n_2484),
.A2(n_2152),
.B1(n_207),
.B2(n_204),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2481),
.Y(n_2541)
);

AOI21xp5_ASAP7_75t_L g2542 ( 
.A1(n_2467),
.A2(n_206),
.B(n_207),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2481),
.Y(n_2543)
);

OAI221xp5_ASAP7_75t_L g2544 ( 
.A1(n_2467),
.A2(n_209),
.B1(n_206),
.B2(n_208),
.C(n_210),
.Y(n_2544)
);

AOI22xp5_ASAP7_75t_L g2545 ( 
.A1(n_2452),
.A2(n_211),
.B1(n_208),
.B2(n_209),
.Y(n_2545)
);

AOI321xp33_ASAP7_75t_L g2546 ( 
.A1(n_2467),
.A2(n_215),
.A3(n_217),
.B1(n_213),
.B2(n_214),
.C(n_216),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2481),
.Y(n_2547)
);

AOI221xp5_ASAP7_75t_L g2548 ( 
.A1(n_2467),
.A2(n_217),
.B1(n_213),
.B2(n_214),
.C(n_218),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_L g2549 ( 
.A(n_2467),
.B(n_218),
.Y(n_2549)
);

OAI21xp5_ASAP7_75t_SL g2550 ( 
.A1(n_2498),
.A2(n_219),
.B(n_220),
.Y(n_2550)
);

OAI21xp33_ASAP7_75t_L g2551 ( 
.A1(n_2521),
.A2(n_219),
.B(n_220),
.Y(n_2551)
);

NAND2x1_ASAP7_75t_SL g2552 ( 
.A(n_2520),
.B(n_221),
.Y(n_2552)
);

AOI221xp5_ASAP7_75t_L g2553 ( 
.A1(n_2549),
.A2(n_2541),
.B1(n_2547),
.B2(n_2543),
.C(n_2536),
.Y(n_2553)
);

NOR3xp33_ASAP7_75t_L g2554 ( 
.A(n_2486),
.B(n_2525),
.C(n_2518),
.Y(n_2554)
);

OAI321xp33_ASAP7_75t_L g2555 ( 
.A1(n_2505),
.A2(n_224),
.A3(n_226),
.B1(n_221),
.B2(n_223),
.C(n_225),
.Y(n_2555)
);

OAI221xp5_ASAP7_75t_L g2556 ( 
.A1(n_2526),
.A2(n_2537),
.B1(n_2535),
.B2(n_2528),
.C(n_2531),
.Y(n_2556)
);

NAND3xp33_ASAP7_75t_L g2557 ( 
.A(n_2489),
.B(n_223),
.C(n_224),
.Y(n_2557)
);

OAI211xp5_ASAP7_75t_L g2558 ( 
.A1(n_2519),
.A2(n_227),
.B(n_225),
.C(n_226),
.Y(n_2558)
);

NOR3xp33_ASAP7_75t_L g2559 ( 
.A(n_2502),
.B(n_227),
.C(n_228),
.Y(n_2559)
);

NAND4xp25_ASAP7_75t_L g2560 ( 
.A(n_2500),
.B(n_230),
.C(n_228),
.D(n_229),
.Y(n_2560)
);

NAND4xp25_ASAP7_75t_L g2561 ( 
.A(n_2534),
.B(n_231),
.C(n_229),
.D(n_230),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2490),
.Y(n_2562)
);

AOI211xp5_ASAP7_75t_L g2563 ( 
.A1(n_2523),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_2563)
);

NAND3xp33_ASAP7_75t_L g2564 ( 
.A(n_2503),
.B(n_232),
.C(n_233),
.Y(n_2564)
);

AOI221xp5_ASAP7_75t_L g2565 ( 
.A1(n_2510),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.C(n_237),
.Y(n_2565)
);

AOI321xp33_ASAP7_75t_L g2566 ( 
.A1(n_2509),
.A2(n_238),
.A3(n_240),
.B1(n_236),
.B2(n_237),
.C(n_239),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2533),
.Y(n_2567)
);

NAND5xp2_ASAP7_75t_L g2568 ( 
.A(n_2513),
.B(n_241),
.C(n_238),
.D(n_239),
.E(n_242),
.Y(n_2568)
);

AOI22xp5_ASAP7_75t_L g2569 ( 
.A1(n_2529),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_2569)
);

AOI22xp5_ASAP7_75t_L g2570 ( 
.A1(n_2488),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.Y(n_2570)
);

AOI221xp5_ASAP7_75t_L g2571 ( 
.A1(n_2524),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.C(n_247),
.Y(n_2571)
);

AOI311xp33_ASAP7_75t_L g2572 ( 
.A1(n_2515),
.A2(n_249),
.A3(n_247),
.B(n_248),
.C(n_250),
.Y(n_2572)
);

OAI211xp5_ASAP7_75t_SL g2573 ( 
.A1(n_2493),
.A2(n_251),
.B(n_248),
.C(n_249),
.Y(n_2573)
);

NOR2xp33_ASAP7_75t_L g2574 ( 
.A(n_2499),
.B(n_251),
.Y(n_2574)
);

A2O1A1Ixp33_ASAP7_75t_L g2575 ( 
.A1(n_2542),
.A2(n_254),
.B(n_252),
.C(n_253),
.Y(n_2575)
);

NOR2xp33_ASAP7_75t_SL g2576 ( 
.A(n_2487),
.B(n_252),
.Y(n_2576)
);

AOI221xp5_ASAP7_75t_L g2577 ( 
.A1(n_2522),
.A2(n_257),
.B1(n_253),
.B2(n_255),
.C(n_258),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2546),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_SL g2579 ( 
.A(n_2546),
.B(n_255),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2497),
.B(n_257),
.Y(n_2580)
);

AOI221xp5_ASAP7_75t_L g2581 ( 
.A1(n_2506),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.C(n_261),
.Y(n_2581)
);

O2A1O1Ixp33_ASAP7_75t_L g2582 ( 
.A1(n_2538),
.A2(n_263),
.B(n_261),
.C(n_262),
.Y(n_2582)
);

AOI22x1_ASAP7_75t_SL g2583 ( 
.A1(n_2530),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.Y(n_2583)
);

NOR2x1_ASAP7_75t_L g2584 ( 
.A(n_2544),
.B(n_264),
.Y(n_2584)
);

OAI322xp33_ASAP7_75t_L g2585 ( 
.A1(n_2507),
.A2(n_271),
.A3(n_270),
.B1(n_268),
.B2(n_266),
.C1(n_267),
.C2(n_269),
.Y(n_2585)
);

AOI21xp33_ASAP7_75t_L g2586 ( 
.A1(n_2501),
.A2(n_268),
.B(n_270),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2527),
.B(n_271),
.Y(n_2587)
);

OAI21xp33_ASAP7_75t_SL g2588 ( 
.A1(n_2545),
.A2(n_272),
.B(n_273),
.Y(n_2588)
);

OAI221xp5_ASAP7_75t_L g2589 ( 
.A1(n_2492),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.C(n_277),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2504),
.Y(n_2590)
);

AOI21xp5_ASAP7_75t_L g2591 ( 
.A1(n_2539),
.A2(n_274),
.B(n_276),
.Y(n_2591)
);

AOI222xp33_ASAP7_75t_L g2592 ( 
.A1(n_2514),
.A2(n_279),
.B1(n_281),
.B2(n_277),
.C1(n_278),
.C2(n_280),
.Y(n_2592)
);

OAI211xp5_ASAP7_75t_L g2593 ( 
.A1(n_2548),
.A2(n_281),
.B(n_279),
.C(n_280),
.Y(n_2593)
);

OAI221xp5_ASAP7_75t_L g2594 ( 
.A1(n_2495),
.A2(n_2508),
.B1(n_2496),
.B2(n_2511),
.C(n_2516),
.Y(n_2594)
);

AOI221xp5_ASAP7_75t_L g2595 ( 
.A1(n_2512),
.A2(n_2517),
.B1(n_2532),
.B2(n_2491),
.C(n_2540),
.Y(n_2595)
);

OAI221xp5_ASAP7_75t_L g2596 ( 
.A1(n_2494),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.C(n_285),
.Y(n_2596)
);

NOR2xp33_ASAP7_75t_SL g2597 ( 
.A(n_2487),
.B(n_282),
.Y(n_2597)
);

A2O1A1Ixp33_ASAP7_75t_L g2598 ( 
.A1(n_2549),
.A2(n_287),
.B(n_285),
.C(n_286),
.Y(n_2598)
);

OAI22xp5_ASAP7_75t_L g2599 ( 
.A1(n_2486),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.Y(n_2599)
);

OAI221xp5_ASAP7_75t_L g2600 ( 
.A1(n_2486),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.C(n_291),
.Y(n_2600)
);

AOI22xp5_ASAP7_75t_L g2601 ( 
.A1(n_2549),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_2601)
);

AOI221xp5_ASAP7_75t_L g2602 ( 
.A1(n_2549),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.C(n_295),
.Y(n_2602)
);

NOR3xp33_ASAP7_75t_SL g2603 ( 
.A(n_2549),
.B(n_294),
.C(n_296),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2490),
.Y(n_2604)
);

OAI21xp33_ASAP7_75t_SL g2605 ( 
.A1(n_2503),
.A2(n_296),
.B(n_297),
.Y(n_2605)
);

INVx2_ASAP7_75t_SL g2606 ( 
.A(n_2499),
.Y(n_2606)
);

NOR4xp25_ASAP7_75t_L g2607 ( 
.A(n_2486),
.B(n_299),
.C(n_297),
.D(n_298),
.Y(n_2607)
);

O2A1O1Ixp33_ASAP7_75t_L g2608 ( 
.A1(n_2486),
.A2(n_300),
.B(n_298),
.C(n_299),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2490),
.B(n_301),
.Y(n_2609)
);

AOI21xp5_ASAP7_75t_L g2610 ( 
.A1(n_2486),
.A2(n_301),
.B(n_302),
.Y(n_2610)
);

NAND4xp25_ASAP7_75t_L g2611 ( 
.A(n_2549),
.B(n_304),
.C(n_302),
.D(n_303),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2490),
.B(n_303),
.Y(n_2612)
);

AOI221xp5_ASAP7_75t_L g2613 ( 
.A1(n_2549),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.C(n_308),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2490),
.Y(n_2614)
);

O2A1O1Ixp33_ASAP7_75t_L g2615 ( 
.A1(n_2486),
.A2(n_308),
.B(n_305),
.C(n_306),
.Y(n_2615)
);

AOI33xp33_ASAP7_75t_L g2616 ( 
.A1(n_2520),
.A2(n_311),
.A3(n_314),
.B1(n_309),
.B2(n_310),
.B3(n_312),
.Y(n_2616)
);

AOI21xp33_ASAP7_75t_L g2617 ( 
.A1(n_2502),
.A2(n_309),
.B(n_311),
.Y(n_2617)
);

A2O1A1Ixp33_ASAP7_75t_L g2618 ( 
.A1(n_2549),
.A2(n_315),
.B(n_312),
.C(n_314),
.Y(n_2618)
);

AOI221xp5_ASAP7_75t_L g2619 ( 
.A1(n_2549),
.A2(n_317),
.B1(n_315),
.B2(n_316),
.C(n_318),
.Y(n_2619)
);

AOI221xp5_ASAP7_75t_L g2620 ( 
.A1(n_2549),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.C(n_320),
.Y(n_2620)
);

AOI221xp5_ASAP7_75t_L g2621 ( 
.A1(n_2549),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.C(n_323),
.Y(n_2621)
);

OAI21xp5_ASAP7_75t_SL g2622 ( 
.A1(n_2498),
.A2(n_322),
.B(n_323),
.Y(n_2622)
);

OAI211xp5_ASAP7_75t_SL g2623 ( 
.A1(n_2536),
.A2(n_326),
.B(n_324),
.C(n_325),
.Y(n_2623)
);

AOI21xp5_ASAP7_75t_L g2624 ( 
.A1(n_2486),
.A2(n_324),
.B(n_325),
.Y(n_2624)
);

AOI221xp5_ASAP7_75t_L g2625 ( 
.A1(n_2549),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.C(n_329),
.Y(n_2625)
);

AOI221xp5_ASAP7_75t_L g2626 ( 
.A1(n_2549),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.C(n_330),
.Y(n_2626)
);

NOR2xp67_ASAP7_75t_L g2627 ( 
.A(n_2555),
.B(n_330),
.Y(n_2627)
);

NOR2x1_ASAP7_75t_L g2628 ( 
.A(n_2560),
.B(n_331),
.Y(n_2628)
);

OAI211xp5_ASAP7_75t_SL g2629 ( 
.A1(n_2553),
.A2(n_2562),
.B(n_2614),
.C(n_2604),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2566),
.B(n_331),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_SL g2631 ( 
.A(n_2578),
.B(n_332),
.Y(n_2631)
);

NOR2xp33_ASAP7_75t_L g2632 ( 
.A(n_2567),
.B(n_332),
.Y(n_2632)
);

NAND3xp33_ASAP7_75t_L g2633 ( 
.A(n_2554),
.B(n_333),
.C(n_334),
.Y(n_2633)
);

OAI211xp5_ASAP7_75t_SL g2634 ( 
.A1(n_2556),
.A2(n_336),
.B(n_333),
.C(n_334),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2606),
.B(n_336),
.Y(n_2635)
);

NOR3xp33_ASAP7_75t_L g2636 ( 
.A(n_2609),
.B(n_2612),
.C(n_2574),
.Y(n_2636)
);

A2O1A1Ixp33_ASAP7_75t_L g2637 ( 
.A1(n_2608),
.A2(n_339),
.B(n_337),
.C(n_338),
.Y(n_2637)
);

OAI21xp5_ASAP7_75t_L g2638 ( 
.A1(n_2579),
.A2(n_337),
.B(n_338),
.Y(n_2638)
);

AOI21xp5_ASAP7_75t_L g2639 ( 
.A1(n_2587),
.A2(n_339),
.B(n_340),
.Y(n_2639)
);

AOI21xp33_ASAP7_75t_L g2640 ( 
.A1(n_2590),
.A2(n_340),
.B(n_341),
.Y(n_2640)
);

AOI22xp5_ASAP7_75t_L g2641 ( 
.A1(n_2551),
.A2(n_343),
.B1(n_341),
.B2(n_342),
.Y(n_2641)
);

NOR2xp33_ASAP7_75t_L g2642 ( 
.A(n_2552),
.B(n_342),
.Y(n_2642)
);

NAND3xp33_ASAP7_75t_L g2643 ( 
.A(n_2576),
.B(n_343),
.C(n_344),
.Y(n_2643)
);

OAI211xp5_ASAP7_75t_L g2644 ( 
.A1(n_2571),
.A2(n_346),
.B(n_344),
.C(n_345),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_SL g2645 ( 
.A(n_2607),
.B(n_347),
.Y(n_2645)
);

NOR2xp33_ASAP7_75t_L g2646 ( 
.A(n_2597),
.B(n_2583),
.Y(n_2646)
);

NAND3xp33_ASAP7_75t_L g2647 ( 
.A(n_2603),
.B(n_348),
.C(n_349),
.Y(n_2647)
);

NOR2xp33_ASAP7_75t_L g2648 ( 
.A(n_2573),
.B(n_349),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2558),
.Y(n_2649)
);

OAI221xp5_ASAP7_75t_L g2650 ( 
.A1(n_2550),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.C(n_353),
.Y(n_2650)
);

AOI21xp33_ASAP7_75t_L g2651 ( 
.A1(n_2615),
.A2(n_352),
.B(n_354),
.Y(n_2651)
);

NAND3xp33_ASAP7_75t_L g2652 ( 
.A(n_2559),
.B(n_355),
.C(n_356),
.Y(n_2652)
);

NAND4xp25_ASAP7_75t_SL g2653 ( 
.A(n_2577),
.B(n_2592),
.C(n_2581),
.D(n_2595),
.Y(n_2653)
);

AOI211x1_ASAP7_75t_L g2654 ( 
.A1(n_2596),
.A2(n_358),
.B(n_356),
.C(n_357),
.Y(n_2654)
);

OAI211xp5_ASAP7_75t_SL g2655 ( 
.A1(n_2586),
.A2(n_359),
.B(n_357),
.C(n_358),
.Y(n_2655)
);

OAI221xp5_ASAP7_75t_SL g2656 ( 
.A1(n_2622),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.C(n_364),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_SL g2657 ( 
.A(n_2572),
.B(n_360),
.Y(n_2657)
);

NAND3xp33_ASAP7_75t_L g2658 ( 
.A(n_2563),
.B(n_2557),
.C(n_2610),
.Y(n_2658)
);

OR2x2_ASAP7_75t_L g2659 ( 
.A(n_2561),
.B(n_364),
.Y(n_2659)
);

NAND3xp33_ASAP7_75t_L g2660 ( 
.A(n_2624),
.B(n_366),
.C(n_367),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2616),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2580),
.Y(n_2662)
);

NOR3xp33_ASAP7_75t_L g2663 ( 
.A(n_2623),
.B(n_367),
.C(n_368),
.Y(n_2663)
);

OAI31xp33_ASAP7_75t_L g2664 ( 
.A1(n_2593),
.A2(n_370),
.A3(n_368),
.B(n_369),
.Y(n_2664)
);

O2A1O1Ixp33_ASAP7_75t_L g2665 ( 
.A1(n_2575),
.A2(n_373),
.B(n_371),
.C(n_372),
.Y(n_2665)
);

NOR4xp25_ASAP7_75t_L g2666 ( 
.A(n_2588),
.B(n_373),
.C(n_371),
.D(n_372),
.Y(n_2666)
);

AND4x1_ASAP7_75t_L g2667 ( 
.A(n_2565),
.B(n_376),
.C(n_374),
.D(n_375),
.Y(n_2667)
);

NOR2x1_ASAP7_75t_L g2668 ( 
.A(n_2611),
.B(n_374),
.Y(n_2668)
);

NAND3xp33_ASAP7_75t_SL g2669 ( 
.A(n_2582),
.B(n_377),
.C(n_378),
.Y(n_2669)
);

NAND4xp25_ASAP7_75t_L g2670 ( 
.A(n_2568),
.B(n_379),
.C(n_377),
.D(n_378),
.Y(n_2670)
);

AOI311xp33_ASAP7_75t_L g2671 ( 
.A1(n_2594),
.A2(n_382),
.A3(n_380),
.B(n_381),
.C(n_383),
.Y(n_2671)
);

NOR2x1_ASAP7_75t_L g2672 ( 
.A(n_2585),
.B(n_380),
.Y(n_2672)
);

NOR2xp33_ASAP7_75t_L g2673 ( 
.A(n_2600),
.B(n_381),
.Y(n_2673)
);

NOR2x1_ASAP7_75t_L g2674 ( 
.A(n_2599),
.B(n_382),
.Y(n_2674)
);

AOI221xp5_ASAP7_75t_L g2675 ( 
.A1(n_2605),
.A2(n_385),
.B1(n_383),
.B2(n_384),
.C(n_386),
.Y(n_2675)
);

NAND3xp33_ASAP7_75t_SL g2676 ( 
.A(n_2591),
.B(n_2601),
.C(n_2602),
.Y(n_2676)
);

NOR2xp33_ASAP7_75t_SL g2677 ( 
.A(n_2617),
.B(n_384),
.Y(n_2677)
);

NAND3xp33_ASAP7_75t_L g2678 ( 
.A(n_2613),
.B(n_388),
.C(n_389),
.Y(n_2678)
);

NAND3xp33_ASAP7_75t_L g2679 ( 
.A(n_2619),
.B(n_390),
.C(n_391),
.Y(n_2679)
);

HB1xp67_ASAP7_75t_L g2680 ( 
.A(n_2584),
.Y(n_2680)
);

NAND4xp75_ASAP7_75t_L g2681 ( 
.A(n_2569),
.B(n_392),
.C(n_390),
.D(n_391),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2598),
.Y(n_2682)
);

INVxp33_ASAP7_75t_L g2683 ( 
.A(n_2620),
.Y(n_2683)
);

INVxp67_ASAP7_75t_L g2684 ( 
.A(n_2564),
.Y(n_2684)
);

O2A1O1Ixp33_ASAP7_75t_L g2685 ( 
.A1(n_2618),
.A2(n_395),
.B(n_393),
.C(n_394),
.Y(n_2685)
);

NOR3xp33_ASAP7_75t_L g2686 ( 
.A(n_2621),
.B(n_394),
.C(n_395),
.Y(n_2686)
);

NOR2xp67_ASAP7_75t_SL g2687 ( 
.A(n_2589),
.B(n_396),
.Y(n_2687)
);

NAND4xp25_ASAP7_75t_L g2688 ( 
.A(n_2570),
.B(n_398),
.C(n_396),
.D(n_397),
.Y(n_2688)
);

AOI221xp5_ASAP7_75t_L g2689 ( 
.A1(n_2625),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.C(n_400),
.Y(n_2689)
);

NAND4xp25_ASAP7_75t_L g2690 ( 
.A(n_2626),
.B(n_402),
.C(n_399),
.D(n_401),
.Y(n_2690)
);

NAND3xp33_ASAP7_75t_SL g2691 ( 
.A(n_2553),
.B(n_403),
.C(n_404),
.Y(n_2691)
);

NOR3xp33_ASAP7_75t_L g2692 ( 
.A(n_2553),
.B(n_403),
.C(n_404),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2562),
.B(n_405),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2562),
.B(n_405),
.Y(n_2694)
);

OAI211xp5_ASAP7_75t_L g2695 ( 
.A1(n_2553),
.A2(n_408),
.B(n_406),
.C(n_407),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2642),
.Y(n_2696)
);

AND3x2_ASAP7_75t_L g2697 ( 
.A(n_2680),
.B(n_406),
.C(n_407),
.Y(n_2697)
);

AOI211xp5_ASAP7_75t_L g2698 ( 
.A1(n_2629),
.A2(n_410),
.B(n_408),
.C(n_409),
.Y(n_2698)
);

NOR4xp75_ASAP7_75t_L g2699 ( 
.A(n_2638),
.B(n_2657),
.C(n_2691),
.D(n_2631),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2646),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2659),
.Y(n_2701)
);

AOI221xp5_ASAP7_75t_L g2702 ( 
.A1(n_2649),
.A2(n_412),
.B1(n_409),
.B2(n_410),
.C(n_413),
.Y(n_2702)
);

AOI221xp5_ASAP7_75t_L g2703 ( 
.A1(n_2632),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.C(n_417),
.Y(n_2703)
);

HB1xp67_ASAP7_75t_L g2704 ( 
.A(n_2627),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2645),
.Y(n_2705)
);

NAND3xp33_ASAP7_75t_L g2706 ( 
.A(n_2636),
.B(n_414),
.C(n_415),
.Y(n_2706)
);

NAND3xp33_ASAP7_75t_SL g2707 ( 
.A(n_2662),
.B(n_416),
.C(n_417),
.Y(n_2707)
);

NOR3xp33_ASAP7_75t_L g2708 ( 
.A(n_2693),
.B(n_418),
.C(n_419),
.Y(n_2708)
);

OR2x2_ASAP7_75t_L g2709 ( 
.A(n_2670),
.B(n_418),
.Y(n_2709)
);

NAND4xp25_ASAP7_75t_L g2710 ( 
.A(n_2639),
.B(n_421),
.C(n_419),
.D(n_420),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2630),
.Y(n_2711)
);

NOR4xp25_ASAP7_75t_L g2712 ( 
.A(n_2653),
.B(n_424),
.C(n_422),
.D(n_423),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2671),
.B(n_2152),
.Y(n_2713)
);

NOR3xp33_ASAP7_75t_L g2714 ( 
.A(n_2694),
.B(n_422),
.C(n_423),
.Y(n_2714)
);

OAI22xp5_ASAP7_75t_L g2715 ( 
.A1(n_2641),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_2715)
);

NAND5xp2_ASAP7_75t_L g2716 ( 
.A(n_2677),
.B(n_425),
.C(n_427),
.D(n_428),
.E(n_429),
.Y(n_2716)
);

NAND3xp33_ASAP7_75t_L g2717 ( 
.A(n_2692),
.B(n_2684),
.C(n_2643),
.Y(n_2717)
);

NAND3xp33_ASAP7_75t_SL g2718 ( 
.A(n_2666),
.B(n_427),
.C(n_428),
.Y(n_2718)
);

NAND4xp25_ASAP7_75t_L g2719 ( 
.A(n_2647),
.B(n_431),
.C(n_429),
.D(n_430),
.Y(n_2719)
);

OAI21xp5_ASAP7_75t_L g2720 ( 
.A1(n_2628),
.A2(n_431),
.B(n_432),
.Y(n_2720)
);

NAND3xp33_ASAP7_75t_SL g2721 ( 
.A(n_2695),
.B(n_432),
.C(n_433),
.Y(n_2721)
);

AOI21xp5_ASAP7_75t_L g2722 ( 
.A1(n_2640),
.A2(n_434),
.B(n_435),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_SL g2723 ( 
.A(n_2664),
.B(n_435),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2668),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2635),
.Y(n_2725)
);

NOR2x1_ASAP7_75t_L g2726 ( 
.A(n_2633),
.B(n_436),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2661),
.B(n_437),
.Y(n_2727)
);

NOR2x1_ASAP7_75t_L g2728 ( 
.A(n_2660),
.B(n_437),
.Y(n_2728)
);

NOR3xp33_ASAP7_75t_SL g2729 ( 
.A(n_2655),
.B(n_438),
.C(n_439),
.Y(n_2729)
);

OAI321xp33_ASAP7_75t_L g2730 ( 
.A1(n_2669),
.A2(n_439),
.A3(n_440),
.B1(n_441),
.B2(n_442),
.C(n_443),
.Y(n_2730)
);

NAND4xp25_ASAP7_75t_L g2731 ( 
.A(n_2648),
.B(n_443),
.C(n_440),
.D(n_442),
.Y(n_2731)
);

NOR3xp33_ASAP7_75t_L g2732 ( 
.A(n_2634),
.B(n_444),
.C(n_445),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2663),
.B(n_444),
.Y(n_2733)
);

NAND3xp33_ASAP7_75t_L g2734 ( 
.A(n_2682),
.B(n_445),
.C(n_446),
.Y(n_2734)
);

AND3x4_ASAP7_75t_L g2735 ( 
.A(n_2667),
.B(n_446),
.C(n_447),
.Y(n_2735)
);

NAND3xp33_ASAP7_75t_L g2736 ( 
.A(n_2675),
.B(n_448),
.C(n_449),
.Y(n_2736)
);

OAI21xp5_ASAP7_75t_L g2737 ( 
.A1(n_2672),
.A2(n_448),
.B(n_449),
.Y(n_2737)
);

AO22x2_ASAP7_75t_L g2738 ( 
.A1(n_2654),
.A2(n_452),
.B1(n_450),
.B2(n_451),
.Y(n_2738)
);

NAND4xp25_ASAP7_75t_L g2739 ( 
.A(n_2658),
.B(n_452),
.C(n_450),
.D(n_451),
.Y(n_2739)
);

NAND3xp33_ASAP7_75t_SL g2740 ( 
.A(n_2683),
.B(n_453),
.C(n_454),
.Y(n_2740)
);

NAND3xp33_ASAP7_75t_L g2741 ( 
.A(n_2652),
.B(n_453),
.C(n_454),
.Y(n_2741)
);

OAI221xp5_ASAP7_75t_L g2742 ( 
.A1(n_2650),
.A2(n_455),
.B1(n_456),
.B2(n_457),
.C(n_458),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2674),
.B(n_455),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2673),
.B(n_457),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2650),
.Y(n_2745)
);

AOI21xp5_ASAP7_75t_L g2746 ( 
.A1(n_2656),
.A2(n_458),
.B(n_459),
.Y(n_2746)
);

OAI221xp5_ASAP7_75t_SL g2747 ( 
.A1(n_2637),
.A2(n_2665),
.B1(n_2685),
.B2(n_2644),
.C(n_2689),
.Y(n_2747)
);

NAND5xp2_ASAP7_75t_L g2748 ( 
.A(n_2651),
.B(n_459),
.C(n_460),
.D(n_461),
.E(n_462),
.Y(n_2748)
);

NAND3xp33_ASAP7_75t_L g2749 ( 
.A(n_2686),
.B(n_460),
.C(n_463),
.Y(n_2749)
);

AOI221x1_ASAP7_75t_L g2750 ( 
.A1(n_2690),
.A2(n_463),
.B1(n_464),
.B2(n_465),
.C(n_466),
.Y(n_2750)
);

AND2x2_ASAP7_75t_L g2751 ( 
.A(n_2704),
.B(n_2681),
.Y(n_2751)
);

NOR2x1_ASAP7_75t_L g2752 ( 
.A(n_2724),
.B(n_2688),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2738),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2697),
.Y(n_2754)
);

AOI22xp5_ASAP7_75t_L g2755 ( 
.A1(n_2700),
.A2(n_2676),
.B1(n_2687),
.B2(n_2679),
.Y(n_2755)
);

NOR3xp33_ASAP7_75t_L g2756 ( 
.A(n_2725),
.B(n_2678),
.C(n_464),
.Y(n_2756)
);

AO22x2_ASAP7_75t_L g2757 ( 
.A1(n_2705),
.A2(n_467),
.B1(n_465),
.B2(n_466),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2743),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2738),
.Y(n_2759)
);

NOR2x1_ASAP7_75t_L g2760 ( 
.A(n_2711),
.B(n_467),
.Y(n_2760)
);

AND3x4_ASAP7_75t_L g2761 ( 
.A(n_2699),
.B(n_2712),
.C(n_2729),
.Y(n_2761)
);

NOR2x1_ASAP7_75t_L g2762 ( 
.A(n_2696),
.B(n_468),
.Y(n_2762)
);

NOR2x1_ASAP7_75t_L g2763 ( 
.A(n_2727),
.B(n_2717),
.Y(n_2763)
);

NOR4xp25_ASAP7_75t_L g2764 ( 
.A(n_2701),
.B(n_471),
.C(n_469),
.D(n_470),
.Y(n_2764)
);

OA22x2_ASAP7_75t_L g2765 ( 
.A1(n_2735),
.A2(n_472),
.B1(n_470),
.B2(n_471),
.Y(n_2765)
);

NOR2xp67_ASAP7_75t_L g2766 ( 
.A(n_2716),
.B(n_2718),
.Y(n_2766)
);

NAND2x1p5_ASAP7_75t_L g2767 ( 
.A(n_2728),
.B(n_473),
.Y(n_2767)
);

INVx1_ASAP7_75t_SL g2768 ( 
.A(n_2709),
.Y(n_2768)
);

AOI22xp5_ASAP7_75t_L g2769 ( 
.A1(n_2745),
.A2(n_475),
.B1(n_473),
.B2(n_474),
.Y(n_2769)
);

NOR2x1_ASAP7_75t_L g2770 ( 
.A(n_2737),
.B(n_474),
.Y(n_2770)
);

AND2x2_ASAP7_75t_L g2771 ( 
.A(n_2720),
.B(n_2231),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2726),
.Y(n_2772)
);

OR2x2_ASAP7_75t_L g2773 ( 
.A(n_2748),
.B(n_475),
.Y(n_2773)
);

OAI22xp5_ASAP7_75t_L g2774 ( 
.A1(n_2698),
.A2(n_479),
.B1(n_476),
.B2(n_477),
.Y(n_2774)
);

NOR2x1_ASAP7_75t_L g2775 ( 
.A(n_2740),
.B(n_477),
.Y(n_2775)
);

HB1xp67_ASAP7_75t_L g2776 ( 
.A(n_2744),
.Y(n_2776)
);

AND3x4_ASAP7_75t_L g2777 ( 
.A(n_2708),
.B(n_479),
.C(n_480),
.Y(n_2777)
);

AND3x4_ASAP7_75t_L g2778 ( 
.A(n_2714),
.B(n_480),
.C(n_481),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2707),
.B(n_481),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2713),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2733),
.Y(n_2781)
);

NOR2x1_ASAP7_75t_L g2782 ( 
.A(n_2734),
.B(n_482),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2723),
.Y(n_2783)
);

INVxp33_ASAP7_75t_SL g2784 ( 
.A(n_2722),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2706),
.Y(n_2785)
);

NOR2x1_ASAP7_75t_L g2786 ( 
.A(n_2731),
.B(n_482),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2750),
.Y(n_2787)
);

NOR2x1_ASAP7_75t_L g2788 ( 
.A(n_2739),
.B(n_483),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_L g2789 ( 
.A(n_2710),
.B(n_484),
.Y(n_2789)
);

NOR2x1_ASAP7_75t_L g2790 ( 
.A(n_2719),
.B(n_485),
.Y(n_2790)
);

NOR2x1_ASAP7_75t_L g2791 ( 
.A(n_2721),
.B(n_486),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2741),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2732),
.Y(n_2793)
);

AOI22xp5_ASAP7_75t_L g2794 ( 
.A1(n_2715),
.A2(n_486),
.B1(n_487),
.B2(n_488),
.Y(n_2794)
);

NOR2xp33_ASAP7_75t_L g2795 ( 
.A(n_2730),
.B(n_487),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2742),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2749),
.Y(n_2797)
);

NOR2xp33_ASAP7_75t_L g2798 ( 
.A(n_2747),
.B(n_489),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2736),
.Y(n_2799)
);

NAND3xp33_ASAP7_75t_L g2800 ( 
.A(n_2759),
.B(n_2703),
.C(n_2702),
.Y(n_2800)
);

NOR2x1_ASAP7_75t_L g2801 ( 
.A(n_2763),
.B(n_2746),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2761),
.Y(n_2802)
);

NAND5xp2_ASAP7_75t_L g2803 ( 
.A(n_2767),
.B(n_490),
.C(n_491),
.D(n_492),
.E(n_493),
.Y(n_2803)
);

NOR3xp33_ASAP7_75t_L g2804 ( 
.A(n_2780),
.B(n_491),
.C(n_492),
.Y(n_2804)
);

INVxp67_ASAP7_75t_L g2805 ( 
.A(n_2776),
.Y(n_2805)
);

AND2x2_ASAP7_75t_L g2806 ( 
.A(n_2753),
.B(n_2231),
.Y(n_2806)
);

NOR3xp33_ASAP7_75t_SL g2807 ( 
.A(n_2758),
.B(n_493),
.C(n_495),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2768),
.B(n_495),
.Y(n_2808)
);

NOR3xp33_ASAP7_75t_L g2809 ( 
.A(n_2781),
.B(n_2754),
.C(n_2772),
.Y(n_2809)
);

NAND4xp25_ASAP7_75t_SL g2810 ( 
.A(n_2794),
.B(n_496),
.C(n_497),
.D(n_498),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2787),
.Y(n_2811)
);

NAND3x1_ASAP7_75t_SL g2812 ( 
.A(n_2752),
.B(n_497),
.C(n_498),
.Y(n_2812)
);

NOR4xp25_ASAP7_75t_L g2813 ( 
.A(n_2751),
.B(n_499),
.C(n_500),
.D(n_501),
.Y(n_2813)
);

NAND4xp75_ASAP7_75t_L g2814 ( 
.A(n_2762),
.B(n_501),
.C(n_502),
.D(n_503),
.Y(n_2814)
);

AND3x4_ASAP7_75t_L g2815 ( 
.A(n_2766),
.B(n_502),
.C(n_503),
.Y(n_2815)
);

NOR3xp33_ASAP7_75t_L g2816 ( 
.A(n_2798),
.B(n_504),
.C(n_505),
.Y(n_2816)
);

NAND2x1p5_ASAP7_75t_L g2817 ( 
.A(n_2770),
.B(n_504),
.Y(n_2817)
);

OAI21xp5_ASAP7_75t_SL g2818 ( 
.A1(n_2755),
.A2(n_506),
.B(n_507),
.Y(n_2818)
);

NAND4xp25_ASAP7_75t_L g2819 ( 
.A(n_2795),
.B(n_508),
.C(n_509),
.D(n_510),
.Y(n_2819)
);

NOR2x1_ASAP7_75t_L g2820 ( 
.A(n_2760),
.B(n_508),
.Y(n_2820)
);

INVxp67_ASAP7_75t_SL g2821 ( 
.A(n_2784),
.Y(n_2821)
);

OAI221xp5_ASAP7_75t_L g2822 ( 
.A1(n_2764),
.A2(n_2773),
.B1(n_2779),
.B2(n_2789),
.C(n_2783),
.Y(n_2822)
);

OR3x1_ASAP7_75t_L g2823 ( 
.A(n_2785),
.B(n_509),
.C(n_510),
.Y(n_2823)
);

NOR3xp33_ASAP7_75t_SL g2824 ( 
.A(n_2793),
.B(n_511),
.C(n_512),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2775),
.B(n_511),
.Y(n_2825)
);

NAND3xp33_ASAP7_75t_L g2826 ( 
.A(n_2799),
.B(n_512),
.C(n_513),
.Y(n_2826)
);

NOR3xp33_ASAP7_75t_SL g2827 ( 
.A(n_2792),
.B(n_513),
.C(n_514),
.Y(n_2827)
);

NAND3x1_ASAP7_75t_L g2828 ( 
.A(n_2791),
.B(n_514),
.C(n_515),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2786),
.B(n_515),
.Y(n_2829)
);

AND2x4_ASAP7_75t_L g2830 ( 
.A(n_2797),
.B(n_516),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2811),
.Y(n_2831)
);

NOR3x2_ASAP7_75t_L g2832 ( 
.A(n_2814),
.B(n_2765),
.C(n_2777),
.Y(n_2832)
);

NAND4xp75_ASAP7_75t_L g2833 ( 
.A(n_2801),
.B(n_2782),
.C(n_2790),
.D(n_2788),
.Y(n_2833)
);

BUFx2_ASAP7_75t_L g2834 ( 
.A(n_2805),
.Y(n_2834)
);

OR2x2_ASAP7_75t_L g2835 ( 
.A(n_2802),
.B(n_2796),
.Y(n_2835)
);

INVx1_ASAP7_75t_SL g2836 ( 
.A(n_2825),
.Y(n_2836)
);

NAND3xp33_ASAP7_75t_SL g2837 ( 
.A(n_2809),
.B(n_2778),
.C(n_2756),
.Y(n_2837)
);

NOR2xp67_ASAP7_75t_L g2838 ( 
.A(n_2803),
.B(n_2769),
.Y(n_2838)
);

AOI221xp5_ASAP7_75t_L g2839 ( 
.A1(n_2821),
.A2(n_2774),
.B1(n_2757),
.B2(n_2771),
.C(n_519),
.Y(n_2839)
);

NAND3x2_ASAP7_75t_L g2840 ( 
.A(n_2830),
.B(n_2757),
.C(n_516),
.Y(n_2840)
);

BUFx2_ASAP7_75t_L g2841 ( 
.A(n_2820),
.Y(n_2841)
);

OAI211xp5_ASAP7_75t_SL g2842 ( 
.A1(n_2822),
.A2(n_517),
.B(n_518),
.C(n_520),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2823),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2817),
.Y(n_2844)
);

OR2x2_ASAP7_75t_L g2845 ( 
.A(n_2829),
.B(n_517),
.Y(n_2845)
);

AND4x1_ASAP7_75t_L g2846 ( 
.A(n_2824),
.B(n_2827),
.C(n_2807),
.D(n_2813),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2808),
.Y(n_2847)
);

INVxp33_ASAP7_75t_SL g2848 ( 
.A(n_2800),
.Y(n_2848)
);

O2A1O1Ixp33_ASAP7_75t_L g2849 ( 
.A1(n_2804),
.A2(n_518),
.B(n_520),
.C(n_521),
.Y(n_2849)
);

NAND5xp2_ASAP7_75t_L g2850 ( 
.A(n_2816),
.B(n_521),
.C(n_522),
.D(n_523),
.E(n_524),
.Y(n_2850)
);

HB1xp67_ASAP7_75t_L g2851 ( 
.A(n_2815),
.Y(n_2851)
);

AND3x2_ASAP7_75t_L g2852 ( 
.A(n_2830),
.B(n_524),
.C(n_525),
.Y(n_2852)
);

OR2x6_ASAP7_75t_L g2853 ( 
.A(n_2828),
.B(n_2818),
.Y(n_2853)
);

AOI21xp5_ASAP7_75t_L g2854 ( 
.A1(n_2819),
.A2(n_526),
.B(n_527),
.Y(n_2854)
);

OAI31xp33_ASAP7_75t_L g2855 ( 
.A1(n_2810),
.A2(n_526),
.A3(n_527),
.B(n_528),
.Y(n_2855)
);

AOI21xp33_ASAP7_75t_L g2856 ( 
.A1(n_2826),
.A2(n_528),
.B(n_529),
.Y(n_2856)
);

HB1xp67_ASAP7_75t_L g2857 ( 
.A(n_2812),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2806),
.Y(n_2858)
);

A2O1A1Ixp33_ASAP7_75t_L g2859 ( 
.A1(n_2805),
.A2(n_529),
.B(n_530),
.C(n_531),
.Y(n_2859)
);

AOI211xp5_ASAP7_75t_L g2860 ( 
.A1(n_2805),
.A2(n_530),
.B(n_532),
.C(n_533),
.Y(n_2860)
);

NOR4xp75_ASAP7_75t_L g2861 ( 
.A(n_2822),
.B(n_533),
.C(n_535),
.D(n_536),
.Y(n_2861)
);

NOR2x1_ASAP7_75t_L g2862 ( 
.A(n_2811),
.B(n_536),
.Y(n_2862)
);

NAND2x1p5_ASAP7_75t_L g2863 ( 
.A(n_2811),
.B(n_537),
.Y(n_2863)
);

NAND4xp25_ASAP7_75t_L g2864 ( 
.A(n_2809),
.B(n_538),
.C(n_539),
.D(n_540),
.Y(n_2864)
);

NAND2x1p5_ASAP7_75t_L g2865 ( 
.A(n_2811),
.B(n_538),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2811),
.Y(n_2866)
);

AOI221xp5_ASAP7_75t_L g2867 ( 
.A1(n_2805),
.A2(n_539),
.B1(n_540),
.B2(n_541),
.C(n_542),
.Y(n_2867)
);

AND2x2_ASAP7_75t_L g2868 ( 
.A(n_2811),
.B(n_2231),
.Y(n_2868)
);

OAI22xp5_ASAP7_75t_SL g2869 ( 
.A1(n_2843),
.A2(n_541),
.B1(n_542),
.B2(n_545),
.Y(n_2869)
);

NOR2xp67_ASAP7_75t_L g2870 ( 
.A(n_2831),
.B(n_545),
.Y(n_2870)
);

NOR4xp25_ASAP7_75t_L g2871 ( 
.A(n_2866),
.B(n_546),
.C(n_547),
.D(n_548),
.Y(n_2871)
);

INVx3_ASAP7_75t_L g2872 ( 
.A(n_2834),
.Y(n_2872)
);

NAND4xp25_ASAP7_75t_L g2873 ( 
.A(n_2848),
.B(n_547),
.C(n_548),
.D(n_549),
.Y(n_2873)
);

AND2x2_ASAP7_75t_L g2874 ( 
.A(n_2841),
.B(n_549),
.Y(n_2874)
);

INVx2_ASAP7_75t_SL g2875 ( 
.A(n_2835),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2833),
.Y(n_2876)
);

AND2x4_ASAP7_75t_L g2877 ( 
.A(n_2844),
.B(n_550),
.Y(n_2877)
);

BUFx2_ASAP7_75t_L g2878 ( 
.A(n_2851),
.Y(n_2878)
);

AOI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2837),
.A2(n_551),
.B(n_552),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2857),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2836),
.B(n_551),
.Y(n_2881)
);

OAI22xp5_ASAP7_75t_L g2882 ( 
.A1(n_2853),
.A2(n_554),
.B1(n_555),
.B2(n_556),
.Y(n_2882)
);

NOR3xp33_ASAP7_75t_SL g2883 ( 
.A(n_2847),
.B(n_554),
.C(n_557),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2832),
.Y(n_2884)
);

OR2x2_ASAP7_75t_L g2885 ( 
.A(n_2840),
.B(n_558),
.Y(n_2885)
);

NOR3xp33_ASAP7_75t_L g2886 ( 
.A(n_2858),
.B(n_558),
.C(n_559),
.Y(n_2886)
);

AND3x4_ASAP7_75t_L g2887 ( 
.A(n_2846),
.B(n_559),
.C(n_560),
.Y(n_2887)
);

AND2x4_ASAP7_75t_L g2888 ( 
.A(n_2838),
.B(n_560),
.Y(n_2888)
);

XOR2x1_ASAP7_75t_L g2889 ( 
.A(n_2863),
.B(n_561),
.Y(n_2889)
);

NAND4xp75_ASAP7_75t_L g2890 ( 
.A(n_2862),
.B(n_561),
.C(n_562),
.D(n_563),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_SL g2891 ( 
.A(n_2839),
.B(n_562),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2853),
.B(n_564),
.Y(n_2892)
);

OR2x2_ASAP7_75t_L g2893 ( 
.A(n_2865),
.B(n_564),
.Y(n_2893)
);

AND2x2_ASAP7_75t_SL g2894 ( 
.A(n_2872),
.B(n_2845),
.Y(n_2894)
);

HB1xp67_ASAP7_75t_L g2895 ( 
.A(n_2875),
.Y(n_2895)
);

HB1xp67_ASAP7_75t_L g2896 ( 
.A(n_2878),
.Y(n_2896)
);

HB1xp67_ASAP7_75t_L g2897 ( 
.A(n_2880),
.Y(n_2897)
);

INVxp67_ASAP7_75t_SL g2898 ( 
.A(n_2876),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2889),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2884),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2870),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2893),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2885),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2888),
.Y(n_2904)
);

HB1xp67_ASAP7_75t_L g2905 ( 
.A(n_2892),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2887),
.Y(n_2906)
);

INVx1_ASAP7_75t_SL g2907 ( 
.A(n_2891),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2881),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2890),
.Y(n_2909)
);

BUFx2_ASAP7_75t_L g2910 ( 
.A(n_2874),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2883),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2877),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2886),
.Y(n_2913)
);

CKINVDCx5p33_ASAP7_75t_R g2914 ( 
.A(n_2896),
.Y(n_2914)
);

NOR2xp33_ASAP7_75t_R g2915 ( 
.A(n_2899),
.B(n_2852),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2897),
.B(n_2871),
.Y(n_2916)
);

NOR2x1_ASAP7_75t_L g2917 ( 
.A(n_2900),
.B(n_2850),
.Y(n_2917)
);

INVxp67_ASAP7_75t_SL g2918 ( 
.A(n_2895),
.Y(n_2918)
);

INVx3_ASAP7_75t_L g2919 ( 
.A(n_2894),
.Y(n_2919)
);

AOI22xp5_ASAP7_75t_L g2920 ( 
.A1(n_2898),
.A2(n_2864),
.B1(n_2842),
.B2(n_2873),
.Y(n_2920)
);

BUFx8_ASAP7_75t_L g2921 ( 
.A(n_2910),
.Y(n_2921)
);

NAND4xp75_ASAP7_75t_L g2922 ( 
.A(n_2901),
.B(n_2879),
.C(n_2855),
.D(n_2854),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2902),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2904),
.Y(n_2924)
);

OAI22xp5_ASAP7_75t_L g2925 ( 
.A1(n_2911),
.A2(n_2849),
.B1(n_2860),
.B2(n_2859),
.Y(n_2925)
);

OAI22x1_ASAP7_75t_L g2926 ( 
.A1(n_2912),
.A2(n_2861),
.B1(n_2868),
.B2(n_2856),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2918),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2919),
.Y(n_2928)
);

OAI22xp5_ASAP7_75t_L g2929 ( 
.A1(n_2914),
.A2(n_2923),
.B1(n_2924),
.B2(n_2916),
.Y(n_2929)
);

OA22x2_ASAP7_75t_L g2930 ( 
.A1(n_2920),
.A2(n_2905),
.B1(n_2906),
.B2(n_2926),
.Y(n_2930)
);

HB1xp67_ASAP7_75t_L g2931 ( 
.A(n_2921),
.Y(n_2931)
);

INVxp67_ASAP7_75t_L g2932 ( 
.A(n_2917),
.Y(n_2932)
);

AND2x4_ASAP7_75t_L g2933 ( 
.A(n_2915),
.B(n_2903),
.Y(n_2933)
);

XNOR2xp5_ASAP7_75t_L g2934 ( 
.A(n_2931),
.B(n_2908),
.Y(n_2934)
);

AOI22x1_ASAP7_75t_L g2935 ( 
.A1(n_2927),
.A2(n_2907),
.B1(n_2909),
.B2(n_2913),
.Y(n_2935)
);

A2O1A1Ixp33_ASAP7_75t_L g2936 ( 
.A1(n_2928),
.A2(n_2925),
.B(n_2867),
.C(n_2882),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_SL g2937 ( 
.A(n_2933),
.B(n_2869),
.Y(n_2937)
);

INVxp33_ASAP7_75t_SL g2938 ( 
.A(n_2929),
.Y(n_2938)
);

AND2x2_ASAP7_75t_L g2939 ( 
.A(n_2932),
.B(n_2922),
.Y(n_2939)
);

XNOR2x1_ASAP7_75t_L g2940 ( 
.A(n_2930),
.B(n_565),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2938),
.B(n_565),
.Y(n_2941)
);

OAI22xp5_ASAP7_75t_L g2942 ( 
.A1(n_2934),
.A2(n_566),
.B1(n_567),
.B2(n_568),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2939),
.Y(n_2943)
);

OAI22xp5_ASAP7_75t_L g2944 ( 
.A1(n_2935),
.A2(n_568),
.B1(n_569),
.B2(n_570),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2943),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_2941),
.Y(n_2946)
);

OAI21xp5_ASAP7_75t_L g2947 ( 
.A1(n_2944),
.A2(n_2937),
.B(n_2940),
.Y(n_2947)
);

OAI22xp5_ASAP7_75t_L g2948 ( 
.A1(n_2945),
.A2(n_2936),
.B1(n_2942),
.B2(n_571),
.Y(n_2948)
);

INVx3_ASAP7_75t_SL g2949 ( 
.A(n_2946),
.Y(n_2949)
);

HB1xp67_ASAP7_75t_L g2950 ( 
.A(n_2947),
.Y(n_2950)
);

AOI221xp5_ASAP7_75t_L g2951 ( 
.A1(n_2950),
.A2(n_569),
.B1(n_570),
.B2(n_572),
.C(n_573),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2949),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2952),
.Y(n_2953)
);

OAI21xp5_ASAP7_75t_SL g2954 ( 
.A1(n_2953),
.A2(n_2948),
.B(n_2951),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2954),
.Y(n_2955)
);

AOI221xp5_ASAP7_75t_L g2956 ( 
.A1(n_2955),
.A2(n_572),
.B1(n_574),
.B2(n_575),
.C(n_576),
.Y(n_2956)
);

OAI221xp5_ASAP7_75t_R g2957 ( 
.A1(n_2956),
.A2(n_574),
.B1(n_575),
.B2(n_576),
.C(n_577),
.Y(n_2957)
);

AOI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_2957),
.A2(n_577),
.B(n_578),
.Y(n_2958)
);

AOI211xp5_ASAP7_75t_L g2959 ( 
.A1(n_2958),
.A2(n_580),
.B(n_581),
.C(n_582),
.Y(n_2959)
);


endmodule