module fake_jpeg_6144_n_323 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_13),
.B(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_38),
.B(n_49),
.Y(n_81)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_25),
.Y(n_41)
);

AO22x1_ASAP7_75t_L g82 ( 
.A1(n_41),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_13),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_13),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_46),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_50),
.Y(n_89)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_21),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_0),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_20),
.B(n_23),
.C(n_21),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_53),
.Y(n_94)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_20),
.B1(n_23),
.B2(n_29),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_54),
.A2(n_60),
.B1(n_73),
.B2(n_75),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_19),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_63),
.Y(n_107)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_57),
.B(n_67),
.Y(n_122)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_58),
.B(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_20),
.B1(n_23),
.B2(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_61),
.B(n_66),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_33),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_29),
.B1(n_28),
.B2(n_24),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_64),
.A2(n_72),
.B1(n_90),
.B2(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_68),
.Y(n_132)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_69),
.B(n_85),
.Y(n_131)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_70),
.B(n_84),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_28),
.B1(n_30),
.B2(n_24),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_39),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_77),
.B1(n_79),
.B2(n_93),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_22),
.B1(n_31),
.B2(n_19),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_22),
.B1(n_26),
.B2(n_17),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_26),
.B1(n_17),
.B2(n_35),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_27),
.B1(n_14),
.B2(n_26),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_88),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_48),
.A2(n_41),
.B1(n_53),
.B2(n_27),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_92),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_36),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_8),
.B(n_9),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_36),
.B(n_27),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_45),
.A2(n_37),
.B1(n_36),
.B2(n_38),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_38),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_45),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_37),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_37),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_8),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_38),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_42),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_43),
.B(n_7),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_8),
.Y(n_109)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_111),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_109),
.B(n_58),
.Y(n_145)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_113),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_114),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_76),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_126),
.A2(n_59),
.B1(n_56),
.B2(n_63),
.Y(n_167)
);

CKINVDCx6p67_ASAP7_75t_R g128 ( 
.A(n_84),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_84),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_9),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_102),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_55),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_133),
.B(n_140),
.Y(n_193)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_142),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_116),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_136),
.B(n_141),
.C(n_155),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_138),
.B(n_145),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_112),
.A2(n_87),
.B1(n_71),
.B2(n_100),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_139),
.A2(n_149),
.B1(n_166),
.B2(n_167),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_81),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_107),
.B(n_55),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_68),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_159),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_71),
.B1(n_65),
.B2(n_90),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_131),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_154),
.Y(n_177)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_92),
.C(n_85),
.Y(n_155)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_160),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_89),
.Y(n_159)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

AND2x6_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_120),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_78),
.C(n_69),
.Y(n_196)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

BUFx24_ASAP7_75t_SL g179 ( 
.A(n_162),
.Y(n_179)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_79),
.B1(n_77),
.B2(n_96),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_165),
.A2(n_119),
.B1(n_118),
.B2(n_105),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_127),
.A2(n_65),
.B1(n_91),
.B2(n_101),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_168),
.Y(n_171)
);

OAI21x1_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_114),
.B(n_116),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_169),
.A2(n_174),
.B(n_191),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_170),
.B(n_199),
.Y(n_225)
);

AO22x1_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_114),
.B1(n_123),
.B2(n_93),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g218 ( 
.A1(n_173),
.A2(n_62),
.B(n_160),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_155),
.B(n_119),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_176),
.A2(n_198),
.B1(n_199),
.B2(n_158),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_105),
.B(n_132),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_189),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_135),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_183),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_184),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_139),
.A2(n_118),
.B1(n_107),
.B2(n_65),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_186),
.B1(n_170),
.B2(n_178),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_107),
.B1(n_91),
.B2(n_86),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_190),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_168),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_188),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_142),
.A2(n_132),
.B(n_109),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_138),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_147),
.A2(n_125),
.B(n_94),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_195),
.Y(n_230)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_202),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_141),
.B(n_117),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_203),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_157),
.A2(n_57),
.B1(n_108),
.B2(n_70),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_157),
.A2(n_76),
.B1(n_62),
.B2(n_117),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_137),
.B(n_84),
.C(n_78),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_137),
.C(n_168),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_153),
.A2(n_11),
.B(n_12),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_11),
.Y(n_203)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_216),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_218),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_211),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_76),
.C(n_140),
.Y(n_211)
);

AO21x2_ASAP7_75t_L g212 ( 
.A1(n_173),
.A2(n_150),
.B(n_143),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_219),
.B1(n_186),
.B2(n_191),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_143),
.C(n_150),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_213),
.B(n_174),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_195),
.A2(n_62),
.B1(n_164),
.B2(n_111),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_215),
.A2(n_220),
.B1(n_223),
.B2(n_176),
.Y(n_237)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_204),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_221),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_173),
.A2(n_111),
.B1(n_134),
.B2(n_154),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_177),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_229),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_169),
.A2(n_178),
.B1(n_185),
.B2(n_196),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_225),
.A2(n_193),
.B(n_205),
.Y(n_252)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_181),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_182),
.B(n_189),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_231),
.B(n_233),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_242),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_249),
.B1(n_255),
.B2(n_209),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_197),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_239),
.A2(n_252),
.B(n_256),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_243),
.B1(n_201),
.B2(n_203),
.Y(n_273)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_212),
.A2(n_187),
.B1(n_190),
.B2(n_175),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_215),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_246),
.Y(n_268)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_228),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_248),
.B(n_250),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_212),
.A2(n_183),
.B1(n_217),
.B2(n_200),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_226),
.B(n_184),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_253),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_213),
.C(n_211),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_216),
.B(n_205),
.Y(n_255)
);

XNOR2x2_ASAP7_75t_SL g256 ( 
.A(n_212),
.B(n_202),
.Y(n_256)
);

AOI221xp5_ASAP7_75t_L g282 ( 
.A1(n_257),
.A2(n_256),
.B1(n_240),
.B2(n_243),
.C(n_234),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_262),
.C(n_263),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_237),
.A2(n_218),
.B1(n_223),
.B2(n_220),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_272),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_207),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_207),
.C(n_232),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_218),
.B1(n_214),
.B2(n_224),
.Y(n_264)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_210),
.C(n_227),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_269),
.C(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_227),
.C(n_229),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_239),
.C(n_234),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_236),
.A2(n_231),
.B1(n_214),
.B2(n_224),
.Y(n_272)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_263),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_282),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_275),
.A2(n_276),
.B(n_281),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_256),
.B(n_248),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_255),
.Y(n_278)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_269),
.B(n_235),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_284),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_260),
.B(n_228),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_242),
.C(n_272),
.Y(n_296)
);

BUFx12f_ASAP7_75t_SL g281 ( 
.A(n_258),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_252),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_260),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_259),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_294),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_266),
.C(n_262),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_291),
.A2(n_292),
.B(n_296),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_271),
.C(n_273),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_208),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_276),
.B(n_238),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_261),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_297),
.A2(n_299),
.B(n_278),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_268),
.C(n_239),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_292),
.B(n_179),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_300),
.B(n_308),
.Y(n_310)
);

NOR3xp33_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_281),
.C(n_285),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_307),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_290),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_299),
.C(n_294),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_295),
.A2(n_283),
.B1(n_270),
.B2(n_245),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_286),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_247),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_244),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_313),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_180),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_180),
.Y(n_317)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g318 ( 
.A1(n_315),
.A2(n_311),
.B(n_238),
.C(n_310),
.D(n_309),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_307),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_318),
.A2(n_319),
.A3(n_308),
.B1(n_247),
.B2(n_303),
.C1(n_316),
.C2(n_312),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_301),
.C(n_291),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_321),
.B(n_171),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_171),
.Y(n_323)
);


endmodule