module fake_jpeg_11370_n_576 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_576);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_576;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_16),
.B(n_14),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_67),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_62),
.A2(n_36),
.B1(n_33),
.B2(n_50),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_8),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_73),
.B(n_77),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_28),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_28),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_79),
.B(n_81),
.Y(n_151)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_80),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_17),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_8),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_83),
.B(n_84),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_6),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_88),
.Y(n_179)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_10),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_90),
.B(n_98),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_28),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_94),
.Y(n_133)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_17),
.Y(n_97)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_21),
.B(n_10),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_21),
.B(n_10),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_100),
.B(n_107),
.Y(n_150)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_24),
.Y(n_101)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_102),
.Y(n_180)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_17),
.Y(n_103)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_106),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_33),
.B(n_5),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_19),
.Y(n_108)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_30),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_109),
.B(n_45),
.Y(n_173)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_27),
.Y(n_110)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_81),
.A2(n_51),
.B1(n_49),
.B2(n_25),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_118),
.A2(n_167),
.B1(n_37),
.B2(n_44),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_130),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_56),
.B(n_29),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_131),
.B(n_173),
.Y(n_218)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

INVx6_ASAP7_75t_SL g146 ( 
.A(n_82),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_146),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_75),
.A2(n_35),
.B(n_34),
.C(n_40),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_149),
.B(n_174),
.Y(n_205)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_72),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

BUFx12_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_57),
.B(n_52),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_169),
.Y(n_206)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_65),
.Y(n_166)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_58),
.B(n_34),
.Y(n_169)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_63),
.Y(n_170)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_64),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_65),
.Y(n_172)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_85),
.Y(n_174)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_74),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_61),
.B(n_36),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_117),
.Y(n_214)
);

INVx4_ASAP7_75t_SL g183 ( 
.A(n_103),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_105),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_71),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_184),
.B(n_186),
.Y(n_207)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_86),
.Y(n_185)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_88),
.B(n_37),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_192),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_193),
.Y(n_280)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_114),
.Y(n_195)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_195),
.Y(n_256)
);

CKINVDCx12_ASAP7_75t_R g196 ( 
.A(n_133),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_196),
.Y(n_276)
);

CKINVDCx12_ASAP7_75t_R g197 ( 
.A(n_125),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_197),
.Y(n_309)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_115),
.Y(n_198)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_198),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_199),
.B(n_204),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_164),
.A2(n_169),
.B1(n_112),
.B2(n_87),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_201),
.A2(n_211),
.B1(n_232),
.B2(n_254),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_130),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_202),
.B(n_214),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_203),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_137),
.B(n_29),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_208),
.B(n_219),
.Y(n_298)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_209),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_210),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_153),
.A2(n_101),
.B1(n_111),
.B2(n_110),
.Y(n_211)
);

CKINVDCx12_ASAP7_75t_R g212 ( 
.A(n_152),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_212),
.Y(n_288)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_116),
.Y(n_213)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_213),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_150),
.B(n_50),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_215),
.B(n_220),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_216),
.A2(n_121),
.B1(n_93),
.B2(n_92),
.Y(n_270)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_120),
.Y(n_217)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_137),
.B(n_52),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_117),
.B(n_139),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_131),
.B(n_165),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_221),
.B(n_239),
.Y(n_265)
);

AND2x2_ASAP7_75t_SL g222 ( 
.A(n_126),
.B(n_160),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_222),
.B(n_247),
.Y(n_295)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_154),
.Y(n_224)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_123),
.Y(n_226)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_226),
.Y(n_299)
);

BUFx12f_ASAP7_75t_L g228 ( 
.A(n_135),
.Y(n_228)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_228),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_141),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_230),
.B(n_231),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_165),
.B(n_44),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_156),
.A2(n_76),
.B1(n_102),
.B2(n_96),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_170),
.A2(n_49),
.B1(n_51),
.B2(n_25),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_233),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_122),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

CKINVDCx12_ASAP7_75t_R g235 ( 
.A(n_163),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_235),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_145),
.B(n_38),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_236),
.B(n_246),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_176),
.B(n_113),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_237),
.B(n_245),
.Y(n_258)
);

AO22x1_ASAP7_75t_L g238 ( 
.A1(n_167),
.A2(n_47),
.B1(n_40),
.B2(n_32),
.Y(n_238)
);

O2A1O1Ixp33_ASAP7_75t_L g282 ( 
.A1(n_238),
.A2(n_251),
.B(n_161),
.C(n_144),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_143),
.B(n_47),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_159),
.Y(n_241)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_241),
.Y(n_272)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_147),
.Y(n_242)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_242),
.Y(n_285)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_168),
.Y(n_243)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_243),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_118),
.A2(n_106),
.B1(n_80),
.B2(n_38),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_66),
.B1(n_95),
.B2(n_127),
.Y(n_255)
);

AOI21xp33_ASAP7_75t_L g245 ( 
.A1(n_122),
.A2(n_32),
.B(n_144),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_183),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_132),
.B(n_0),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_157),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_248),
.B(n_249),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_128),
.B(n_119),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_140),
.Y(n_250)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_250),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_124),
.A2(n_91),
.B(n_70),
.C(n_104),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_175),
.A2(n_48),
.B1(n_54),
.B2(n_51),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_180),
.B1(n_148),
.B2(n_140),
.Y(n_273)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_129),
.Y(n_253)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_253),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_175),
.A2(n_49),
.B1(n_48),
.B2(n_53),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_255),
.A2(n_259),
.B1(n_269),
.B2(n_270),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_199),
.A2(n_129),
.B1(n_134),
.B2(n_124),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_204),
.A2(n_205),
.B1(n_221),
.B2(n_206),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_267),
.A2(n_273),
.B1(n_278),
.B2(n_281),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_238),
.A2(n_134),
.B1(n_119),
.B2(n_180),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_247),
.A2(n_148),
.B1(n_177),
.B2(n_53),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_277),
.A2(n_279),
.B1(n_290),
.B2(n_294),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_252),
.A2(n_158),
.B1(n_138),
.B2(n_171),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_218),
.A2(n_138),
.B1(n_158),
.B2(n_3),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_208),
.A2(n_219),
.B1(n_207),
.B2(n_239),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_289),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_190),
.A2(n_250),
.B1(n_189),
.B2(n_194),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_190),
.A2(n_161),
.B1(n_0),
.B2(n_3),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_189),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_210),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_194),
.A2(n_4),
.B1(n_5),
.B2(n_11),
.Y(n_291)
);

A2O1A1Ixp33_ASAP7_75t_SL g351 ( 
.A1(n_291),
.A2(n_304),
.B(n_284),
.C(n_271),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_222),
.A2(n_4),
.B1(n_12),
.B2(n_13),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_222),
.A2(n_0),
.B1(n_15),
.B2(n_210),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_195),
.Y(n_305)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_305),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_198),
.B(n_217),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_306),
.A2(n_193),
.B(n_188),
.Y(n_339)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_225),
.Y(n_307)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_251),
.A2(n_209),
.B1(n_229),
.B2(n_213),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_311),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_203),
.A2(n_226),
.B1(n_253),
.B2(n_240),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_312),
.A2(n_192),
.B1(n_187),
.B2(n_188),
.Y(n_338)
);

AND2x6_ASAP7_75t_L g313 ( 
.A(n_258),
.B(n_227),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_313),
.B(n_347),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_265),
.B(n_242),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_315),
.B(n_323),
.Y(n_395)
);

INVx13_ASAP7_75t_L g316 ( 
.A(n_280),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_316),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_264),
.B(n_191),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_317),
.B(n_353),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_223),
.C(n_200),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_318),
.B(n_340),
.C(n_339),
.Y(n_396)
);

INVx6_ASAP7_75t_SL g319 ( 
.A(n_276),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_319),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_308),
.A2(n_229),
.B1(n_234),
.B2(n_187),
.Y(n_321)
);

OAI22x1_ASAP7_75t_L g373 ( 
.A1(n_321),
.A2(n_310),
.B1(n_303),
.B2(n_296),
.Y(n_373)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_272),
.Y(n_322)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_322),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_224),
.Y(n_323)
);

INVx11_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g368 ( 
.A(n_324),
.Y(n_368)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_272),
.Y(n_325)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_325),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_261),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_326),
.B(n_327),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_295),
.B(n_191),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_328),
.Y(n_381)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_292),
.Y(n_329)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_329),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_275),
.B(n_301),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_330),
.B(n_332),
.Y(n_388)
);

INVx13_ASAP7_75t_L g331 ( 
.A(n_309),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_331),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_286),
.B(n_200),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_307),
.Y(n_334)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_334),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_293),
.B(n_188),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_335),
.B(n_341),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_338),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_339),
.B(n_349),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_281),
.B(n_193),
.C(n_228),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_293),
.B(n_228),
.Y(n_341)
);

INVx13_ASAP7_75t_L g342 ( 
.A(n_288),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_342),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_298),
.B(n_258),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_344),
.B(n_348),
.Y(n_401)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_302),
.Y(n_345)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_345),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_299),
.Y(n_346)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_346),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_306),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_295),
.B(n_298),
.Y(n_348)
);

INVx13_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_299),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_350),
.B(n_354),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_351),
.A2(n_289),
.B1(n_283),
.B2(n_312),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_304),
.B(n_287),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_294),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_300),
.B(n_263),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_302),
.Y(n_354)
);

AND2x6_ASAP7_75t_L g355 ( 
.A(n_282),
.B(n_270),
.Y(n_355)
);

MAJx2_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_360),
.C(n_256),
.Y(n_382)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_306),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_357),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_300),
.B(n_263),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_257),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_359),
.A2(n_285),
.B(n_274),
.Y(n_378)
);

AND2x6_ASAP7_75t_L g360 ( 
.A(n_308),
.B(n_277),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_348),
.B(n_305),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_361),
.B(n_379),
.C(n_389),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_362),
.B(n_396),
.Y(n_405)
);

OAI32xp33_ASAP7_75t_L g363 ( 
.A1(n_352),
.A2(n_262),
.A3(n_266),
.B1(n_257),
.B2(n_285),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_363),
.B(n_378),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_333),
.A2(n_255),
.B1(n_273),
.B2(n_278),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_371),
.A2(n_376),
.B1(n_387),
.B2(n_390),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_373),
.A2(n_380),
.B(n_346),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_374),
.A2(n_377),
.B1(n_384),
.B2(n_351),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_333),
.A2(n_303),
.B1(n_296),
.B2(n_262),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_336),
.A2(n_262),
.B1(n_266),
.B2(n_296),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_315),
.B(n_256),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_337),
.A2(n_260),
.B(n_268),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_382),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_336),
.A2(n_358),
.B1(n_351),
.B2(n_337),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_343),
.A2(n_274),
.B1(n_268),
.B2(n_260),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_318),
.B(n_327),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_343),
.A2(n_351),
.B1(n_360),
.B2(n_323),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_351),
.A2(n_355),
.B1(n_340),
.B2(n_347),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_397),
.A2(n_358),
.B1(n_346),
.B2(n_320),
.Y(n_427)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_366),
.Y(n_402)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_402),
.Y(n_452)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_366),
.Y(n_403)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_403),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_397),
.B(n_356),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_404),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_406),
.B(n_407),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_393),
.Y(n_407)
);

BUFx10_ASAP7_75t_L g409 ( 
.A(n_385),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_409),
.Y(n_446)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_370),
.Y(n_410)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_410),
.Y(n_463)
);

INVx13_ASAP7_75t_L g412 ( 
.A(n_365),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_412),
.Y(n_449)
);

AOI32xp33_ASAP7_75t_L g413 ( 
.A1(n_401),
.A2(n_313),
.A3(n_317),
.B1(n_319),
.B2(n_324),
.Y(n_413)
);

AOI21xp33_ASAP7_75t_L g458 ( 
.A1(n_413),
.A2(n_419),
.B(n_428),
.Y(n_458)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_370),
.Y(n_414)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_414),
.Y(n_466)
);

NOR3xp33_ASAP7_75t_L g415 ( 
.A(n_364),
.B(n_331),
.C(n_342),
.Y(n_415)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_431),
.C(n_435),
.Y(n_444)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_367),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_416),
.B(n_418),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_375),
.Y(n_418)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_382),
.B(n_331),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_381),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_420),
.B(n_422),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_421),
.A2(n_380),
.B(n_398),
.Y(n_453)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_381),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_375),
.B(n_334),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_423),
.B(n_424),
.Y(n_447)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_391),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_425),
.B(n_429),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_427),
.A2(n_434),
.B1(n_374),
.B2(n_384),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_390),
.A2(n_329),
.B(n_328),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_363),
.B(n_325),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_399),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_430),
.B(n_436),
.Y(n_448)
);

OAI21xp33_ASAP7_75t_L g431 ( 
.A1(n_372),
.A2(n_322),
.B(n_320),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_361),
.B(n_314),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_432),
.B(n_433),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_395),
.B(n_314),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_371),
.A2(n_350),
.B1(n_359),
.B2(n_354),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_388),
.B(n_345),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_386),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_418),
.B(n_369),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_438),
.B(n_442),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_439),
.A2(n_443),
.B1(n_455),
.B2(n_406),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_417),
.B(n_389),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_440),
.B(n_445),
.C(n_450),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_423),
.B(n_369),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_408),
.A2(n_377),
.B1(n_395),
.B2(n_398),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_417),
.B(n_396),
.C(n_379),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_405),
.B(n_362),
.C(n_383),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_407),
.B(n_386),
.Y(n_451)
);

INVxp33_ASAP7_75t_L g470 ( 
.A(n_451),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_453),
.A2(n_461),
.B(n_411),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_408),
.A2(n_387),
.B1(n_376),
.B2(n_392),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_436),
.B(n_392),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_456),
.B(n_457),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_426),
.B(n_368),
.Y(n_457)
);

AO22x1_ASAP7_75t_L g461 ( 
.A1(n_428),
.A2(n_378),
.B1(n_394),
.B2(n_400),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_432),
.B(n_383),
.C(n_367),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_467),
.C(n_404),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_383),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_464),
.B(n_429),
.Y(n_468)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_468),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_437),
.A2(n_427),
.B1(n_411),
.B2(n_426),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_471),
.A2(n_439),
.B1(n_443),
.B2(n_467),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_472),
.B(n_481),
.Y(n_502)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_447),
.Y(n_473)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_473),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_464),
.B(n_447),
.Y(n_476)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_476),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_477),
.B(n_465),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_448),
.B(n_410),
.Y(n_478)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_478),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_479),
.A2(n_482),
.B1(n_484),
.B2(n_485),
.Y(n_514)
);

A2O1A1Ixp33_ASAP7_75t_L g480 ( 
.A1(n_437),
.A2(n_404),
.B(n_421),
.C(n_419),
.Y(n_480)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_480),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_438),
.B(n_404),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_462),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_440),
.B(n_434),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_483),
.B(n_487),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_442),
.B(n_444),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_409),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_462),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_486),
.A2(n_488),
.B1(n_490),
.B2(n_466),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_454),
.B(n_425),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_460),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_460),
.B(n_424),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_489),
.B(n_492),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_449),
.B(n_409),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_445),
.B(n_403),
.C(n_420),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_491),
.B(n_493),
.C(n_441),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_458),
.A2(n_409),
.B(n_394),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_450),
.B(n_402),
.C(n_414),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_495),
.B(n_482),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_496),
.A2(n_503),
.B1(n_479),
.B2(n_486),
.Y(n_519)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_497),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_474),
.A2(n_453),
.B1(n_466),
.B2(n_459),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_498),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_472),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_491),
.B(n_441),
.C(n_455),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_500),
.B(n_501),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_469),
.B(n_446),
.C(n_459),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_471),
.A2(n_461),
.B1(n_446),
.B2(n_452),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_469),
.B(n_446),
.C(n_463),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_504),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_474),
.A2(n_463),
.B1(n_452),
.B2(n_422),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_505),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_461),
.C(n_400),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_511),
.B(n_512),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_483),
.B(n_416),
.C(n_373),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_477),
.B(n_449),
.C(n_349),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_490),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_519),
.A2(n_529),
.B1(n_515),
.B2(n_488),
.Y(n_546)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_507),
.Y(n_520)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_520),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_521),
.A2(n_500),
.B(n_492),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_522),
.B(n_513),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_523),
.B(n_501),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_502),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_527),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_514),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_506),
.Y(n_528)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_528),
.Y(n_541)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_494),
.Y(n_529)
);

FAx1_ASAP7_75t_SL g530 ( 
.A(n_511),
.B(n_481),
.CI(n_476),
.CON(n_530),
.SN(n_530)
);

BUFx24_ASAP7_75t_SL g545 ( 
.A(n_530),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_508),
.B(n_470),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_532),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_521),
.B(n_495),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_533),
.B(n_534),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_531),
.B(n_504),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_535),
.B(n_536),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_525),
.A2(n_496),
.B1(n_503),
.B2(n_473),
.Y(n_536)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_539),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_517),
.B(n_499),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_542),
.B(n_543),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_516),
.B(n_509),
.C(n_512),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_544),
.B(n_522),
.C(n_524),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_546),
.B(n_530),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_550),
.B(n_551),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_538),
.B(n_478),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_553),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_545),
.A2(n_525),
.B1(n_518),
.B2(n_520),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_554),
.A2(n_541),
.B1(n_537),
.B2(n_528),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_534),
.B(n_475),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_555),
.B(n_475),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_533),
.B(n_518),
.C(n_509),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_556),
.B(n_544),
.C(n_542),
.Y(n_561)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_558),
.Y(n_566)
);

INVx11_ASAP7_75t_L g559 ( 
.A(n_548),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_559),
.B(n_561),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_SL g560 ( 
.A1(n_552),
.A2(n_540),
.B(n_529),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_560),
.A2(n_562),
.B1(n_468),
.B2(n_489),
.Y(n_567)
);

AOI322xp5_ASAP7_75t_L g564 ( 
.A1(n_563),
.A2(n_547),
.A3(n_530),
.B1(n_553),
.B2(n_480),
.C1(n_539),
.C2(n_549),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_564),
.B(n_557),
.Y(n_569)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_567),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_569),
.B(n_556),
.Y(n_571)
);

AOI321xp33_ASAP7_75t_L g570 ( 
.A1(n_568),
.A2(n_566),
.A3(n_565),
.B1(n_549),
.B2(n_563),
.C(n_560),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g572 ( 
.A1(n_570),
.A2(n_571),
.B(n_487),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_572),
.A2(n_510),
.B1(n_412),
.B2(n_349),
.Y(n_573)
);

BUFx24_ASAP7_75t_SL g574 ( 
.A(n_573),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_574),
.B(n_510),
.C(n_316),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_575),
.B(n_316),
.Y(n_576)
);


endmodule