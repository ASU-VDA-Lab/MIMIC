module fake_jpeg_8798_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_1),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_30),
.Y(n_61)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_48),
.B(n_27),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_22),
.B1(n_48),
.B2(n_46),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_49),
.A2(n_46),
.B1(n_48),
.B2(n_45),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_22),
.B1(n_34),
.B2(n_30),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_58),
.B1(n_62),
.B2(n_34),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_20),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_43),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_22),
.B1(n_34),
.B2(n_35),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_34),
.B1(n_35),
.B2(n_30),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_39),
.C(n_42),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_32),
.Y(n_120)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_92),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_74),
.A2(n_37),
.B1(n_40),
.B2(n_33),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_79),
.B(n_87),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_88),
.B(n_91),
.Y(n_110)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_56),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g93 ( 
.A1(n_50),
.A2(n_42),
.B(n_30),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_98),
.B(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_97),
.B1(n_57),
.B2(n_69),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_40),
.B1(n_52),
.B2(n_64),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_63),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_45),
.B1(n_48),
.B2(n_57),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_99),
.A2(n_100),
.B1(n_89),
.B2(n_85),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_45),
.B1(n_48),
.B2(n_57),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_112),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_63),
.B(n_65),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_104),
.A2(n_114),
.B(n_32),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_116),
.B1(n_118),
.B2(n_121),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_65),
.B1(n_35),
.B2(n_56),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_71),
.Y(n_108)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_31),
.B1(n_29),
.B2(n_32),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_19),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_119),
.B(n_31),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_78),
.B(n_75),
.Y(n_129)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_123),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_75),
.A2(n_40),
.B1(n_66),
.B2(n_44),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_111),
.B1(n_122),
.B2(n_113),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_128),
.A2(n_146),
.B1(n_152),
.B2(n_147),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_129),
.A2(n_137),
.B(n_142),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_91),
.C(n_77),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_139),
.C(n_31),
.Y(n_162)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_144),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_40),
.B1(n_92),
.B2(n_89),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_135),
.A2(n_143),
.B1(n_148),
.B2(n_72),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_104),
.A2(n_44),
.B(n_33),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_77),
.C(n_76),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_141),
.B(n_143),
.Y(n_176)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_148),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_89),
.B1(n_76),
.B2(n_70),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_156),
.Y(n_159)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_85),
.B(n_26),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_60),
.B1(n_47),
.B2(n_41),
.Y(n_175)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_155),
.A2(n_123),
.B1(n_103),
.B2(n_60),
.Y(n_168)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_157),
.B(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_160),
.B(n_172),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_120),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_162),
.C(n_173),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_109),
.B1(n_111),
.B2(n_103),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_163),
.A2(n_175),
.B1(n_132),
.B2(n_155),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_167),
.B1(n_170),
.B2(n_179),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_119),
.B(n_20),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_165),
.A2(n_166),
.B(n_171),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_26),
.B(n_20),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_134),
.A2(n_44),
.B1(n_72),
.B2(n_109),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_168),
.A2(n_125),
.B1(n_115),
.B2(n_102),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_134),
.A2(n_142),
.B1(n_131),
.B2(n_154),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_1),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_139),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_47),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_185),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_47),
.C(n_41),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_160),
.C(n_174),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_140),
.A2(n_29),
.B1(n_26),
.B2(n_83),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_136),
.Y(n_201)
);

AO21x2_ASAP7_75t_SL g181 ( 
.A1(n_153),
.A2(n_41),
.B(n_127),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_136),
.B1(n_27),
.B2(n_127),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_182),
.A2(n_25),
.B1(n_28),
.B2(n_27),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_29),
.B(n_23),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_184),
.A2(n_18),
.B(n_24),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_156),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx3_ASAP7_75t_SL g192 ( 
.A(n_186),
.Y(n_192)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_185),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_189),
.Y(n_232)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_169),
.B(n_28),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_193),
.B(n_207),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_102),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_198),
.C(n_213),
.Y(n_224)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

BUFx24_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_190),
.B1(n_211),
.B2(n_191),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_208),
.B(n_183),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_203),
.A2(n_206),
.B1(n_212),
.B2(n_184),
.Y(n_227)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_18),
.B1(n_19),
.B2(n_24),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_205),
.A2(n_209),
.B1(n_214),
.B2(n_17),
.Y(n_240)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_172),
.A2(n_18),
.A3(n_28),
.B1(n_24),
.B2(n_25),
.C1(n_23),
.C2(n_27),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_158),
.B1(n_164),
.B2(n_181),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_167),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_210),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_162),
.B(n_125),
.C(n_95),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_25),
.B1(n_125),
.B2(n_82),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_95),
.C(n_82),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_177),
.C(n_179),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_157),
.Y(n_218)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_218),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_219),
.B(n_244),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_169),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_17),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_222),
.A2(n_223),
.B1(n_227),
.B2(n_229),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_200),
.A2(n_175),
.B1(n_183),
.B2(n_186),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_236),
.C(n_238),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_171),
.Y(n_226)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_199),
.A2(n_196),
.B1(n_209),
.B2(n_193),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_171),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_L g246 ( 
.A1(n_230),
.A2(n_233),
.B(n_215),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_165),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_192),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_2),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_165),
.C(n_166),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_166),
.C(n_28),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_203),
.B1(n_212),
.B2(n_199),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_214),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_242),
.A2(n_208),
.B1(n_213),
.B2(n_11),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_17),
.C(n_3),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_2),
.C(n_3),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_192),
.Y(n_244)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_230),
.B(n_196),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_247),
.B(n_250),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_249),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_221),
.B(n_215),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_237),
.B1(n_228),
.B2(n_241),
.Y(n_251)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_266),
.Y(n_270)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_256),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_17),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_258),
.C(n_259),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_17),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_218),
.A2(n_9),
.B(n_15),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_233),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_262),
.C(n_219),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_10),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_10),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_265),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_234),
.B(n_9),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_223),
.Y(n_266)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

NOR2x1_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_226),
.Y(n_268)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_241),
.B1(n_231),
.B2(n_232),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_269),
.A2(n_275),
.B1(n_282),
.B2(n_261),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_220),
.B1(n_234),
.B2(n_235),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_276),
.B(n_13),
.Y(n_299)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_248),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_284),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_225),
.C(n_238),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_258),
.C(n_245),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_253),
.A2(n_220),
.B1(n_236),
.B2(n_243),
.Y(n_282)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_254),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_246),
.Y(n_285)
);

NAND3xp33_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_269),
.C(n_282),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_247),
.B(n_250),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_287),
.A2(n_281),
.B(n_275),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_273),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_259),
.C(n_257),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_299),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_262),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_297),
.Y(n_312)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_292),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_239),
.B1(n_4),
.B2(n_5),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_294),
.A2(n_295),
.B1(n_279),
.B2(n_283),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_239),
.B1(n_4),
.B2(n_5),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_11),
.Y(n_296)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_12),
.C(n_15),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_270),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_298)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_298),
.Y(n_304)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_311),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_277),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_308),
.Y(n_317)
);

O2A1O1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_288),
.B(n_297),
.C(n_287),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_286),
.B(n_267),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_276),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_310),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_273),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_319),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_289),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_320),
.B(n_322),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_291),
.B1(n_295),
.B2(n_294),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_301),
.C(n_312),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_304),
.A2(n_290),
.B1(n_14),
.B2(n_16),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_305),
.A2(n_14),
.B(n_6),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_5),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_329),
.C(n_322),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_314),
.B(n_306),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_325),
.B(n_6),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_313),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_317),
.Y(n_331)
);

OAI21x1_ASAP7_75t_L g328 ( 
.A1(n_316),
.A2(n_312),
.B(n_311),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_328),
.A2(n_7),
.B(n_8),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_304),
.C(n_14),
.Y(n_329)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_331),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_334),
.A2(n_326),
.B(n_333),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_323),
.C(n_332),
.Y(n_337)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_337),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_335),
.B(n_7),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_8),
.C(n_306),
.Y(n_340)
);


endmodule