module fake_netlist_5_1916_n_88 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_88);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_88;

wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_38;
wire n_80;
wire n_35;
wire n_73;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_85;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_81;
wire n_28;
wire n_70;
wire n_68;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_5),
.Y(n_20)
);

OA21x2_ASAP7_75t_L g21 ( 
.A1(n_15),
.A2(n_7),
.B(n_16),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g22 ( 
.A1(n_14),
.A2(n_4),
.B(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

AND2x4_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

AO22x1_ASAP7_75t_L g29 ( 
.A1(n_8),
.A2(n_2),
.B1(n_10),
.B2(n_6),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_0),
.Y(n_31)
);

OAI21x1_ASAP7_75t_L g32 ( 
.A1(n_0),
.A2(n_3),
.B(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_24),
.Y(n_36)
);

NAND2x1p5_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_22),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_23),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_27),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_22),
.A2(n_33),
.B1(n_35),
.B2(n_28),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_23),
.B(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

OAI21x1_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_32),
.B(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx11_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_27),
.B(n_29),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_42),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_20),
.Y(n_51)
);

OAI21x1_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_37),
.B(n_32),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_47),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_48),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_54),
.Y(n_62)
);

AOI311xp33_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_35),
.A3(n_28),
.B(n_31),
.C(n_20),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_57),
.B(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_54),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_55),
.Y(n_68)
);

AOI211xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_29),
.B(n_31),
.C(n_30),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_60),
.B1(n_21),
.B2(n_22),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_27),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_33),
.B(n_25),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_21),
.B(n_22),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_25),
.B1(n_34),
.B2(n_65),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_63),
.B(n_25),
.C(n_34),
.Y(n_76)
);

OAI221xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_25),
.B1(n_34),
.B2(n_72),
.C(n_75),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_25),
.Y(n_78)
);

NOR4xp25_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_25),
.C(n_34),
.D(n_74),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_34),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_34),
.B1(n_76),
.B2(n_80),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

OA21x2_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_82),
.B(n_81),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_85),
.A2(n_84),
.B1(n_67),
.B2(n_62),
.Y(n_87)
);

AOI31xp33_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_85),
.A3(n_86),
.B(n_84),
.Y(n_88)
);


endmodule