module real_jpeg_24131_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_164;
wire n_48;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_191;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_2),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_2),
.A2(n_25),
.B1(n_33),
.B2(n_36),
.Y(n_79)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_5),
.A2(n_21),
.B1(n_24),
.B2(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_5),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_6),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_6),
.A2(n_35),
.B1(n_51),
.B2(n_53),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_6),
.A2(n_35),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_6),
.A2(n_21),
.B1(n_24),
.B2(n_35),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_8),
.A2(n_33),
.B1(n_36),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_8),
.A2(n_44),
.B1(n_51),
.B2(n_53),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_8),
.A2(n_44),
.B1(n_61),
.B2(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_8),
.A2(n_21),
.B1(n_24),
.B2(n_44),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_8),
.B(n_53),
.C(n_66),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_8),
.B(n_67),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_8),
.B(n_33),
.C(n_49),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_8),
.B(n_21),
.C(n_39),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_8),
.B(n_159),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_8),
.B(n_42),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_8),
.B(n_113),
.Y(n_201)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_9),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_11),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_117),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_116),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_97),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_16),
.B(n_97),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_72),
.C(n_82),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_17),
.B(n_72),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_45),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_SL g115 ( 
.A(n_18),
.B(n_58),
.C(n_70),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_30),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_19),
.A2(n_30),
.B1(n_31),
.B2(n_230),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_19),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_20),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_20),
.B(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_20),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_21),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_21),
.A2(n_24),
.B1(n_39),
.B2(n_40),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_21),
.B(n_191),
.Y(n_190)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_23),
.A2(n_76),
.B(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_28),
.B(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_30),
.A2(n_31),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_30),
.A2(n_31),
.B1(n_170),
.B2(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_31),
.B(n_164),
.C(n_170),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_31),
.B(n_140),
.C(n_201),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_31)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

OA22x2_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_33),
.B(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_43),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_37),
.A2(n_42),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_37),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_41),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_41),
.A2(n_80),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_41),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_43),
.B(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_58),
.B1(n_70),
.B2(n_71),
.Y(n_45)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_46),
.A2(n_70),
.B1(n_128),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_46),
.A2(n_70),
.B1(n_89),
.B2(n_124),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_46),
.B(n_89),
.C(n_208),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B(n_54),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_47),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_47),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_56)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_51),
.Y(n_53)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_53),
.B1(n_65),
.B2(n_66),
.Y(n_67)
);

CKINVDCx6p67_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_53),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_55),
.A2(n_57),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_57),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_58),
.A2(n_71),
.B1(n_111),
.B2(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_58),
.B(n_111),
.C(n_134),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_63),
.B1(n_67),
.B2(n_68),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_67),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_127),
.C(n_128),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_77),
.B1(n_78),
.B2(n_81),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_73),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_73),
.A2(n_81),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_78),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_75),
.B(n_145),
.Y(n_175)
);

INVx3_ASAP7_75t_SL g159 ( 
.A(n_76),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_82),
.B(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_91),
.C(n_94),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_83),
.A2(n_84),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_85),
.A2(n_89),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_85),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_87),
.A2(n_142),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_89),
.A2(n_124),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_89),
.B(n_187),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_91),
.A2(n_94),
.B1(n_127),
.B2(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_91),
.Y(n_227)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_94),
.A2(n_127),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_115),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_106),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_105),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_111),
.B(n_114),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_111),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_157),
.C(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_111),
.A2(n_147),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_233),
.B(n_237),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_160),
.B(n_219),
.C(n_232),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_149),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_120),
.B(n_149),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_133),
.B2(n_148),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_126),
.B1(n_131),
.B2(n_132),
.Y(n_122)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_123),
.B(n_132),
.C(n_148),
.Y(n_220)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_146),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_136),
.B1(n_139),
.B2(n_140),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_139),
.A2(n_140),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_140),
.B(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_140),
.B(n_193),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_140)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_155),
.C(n_156),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_150),
.A2(n_151),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_156),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_158),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_157),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_158),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_218),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_179),
.B(n_217),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_176),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_163),
.B(n_176),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_164),
.A2(n_165),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_169),
.B(n_184),
.Y(n_195)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_210),
.B(n_216),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_204),
.B(n_209),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_196),
.B(n_203),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_188),
.B(n_195),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_185),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_192),
.B(n_194),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_197),
.B(n_198),
.Y(n_203)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_205),
.B(n_206),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_211),
.B(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_221),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_231),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_228),
.B2(n_229),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_229),
.C(n_231),
.Y(n_234)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_235),
.Y(n_237)
);


endmodule