module real_jpeg_14286_n_16 (n_5, n_4, n_8, n_0, n_12, n_324, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_324;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_4),
.A2(n_48),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_4),
.A2(n_32),
.B1(n_35),
.B2(n_48),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_4),
.A2(n_48),
.B1(n_74),
.B2(n_75),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_5),
.A2(n_74),
.B1(n_75),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_5),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_135),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_135),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_5),
.A2(n_32),
.B1(n_35),
.B2(n_135),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_6),
.A2(n_56),
.B1(n_62),
.B2(n_63),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_6),
.A2(n_32),
.B1(n_35),
.B2(n_56),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_6),
.A2(n_56),
.B1(n_74),
.B2(n_75),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_7),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_7),
.A2(n_34),
.B1(n_74),
.B2(n_75),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_7),
.A2(n_34),
.B1(n_45),
.B2(n_46),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_7),
.A2(n_34),
.B1(n_62),
.B2(n_63),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_10),
.A2(n_73),
.B(n_74),
.C(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_10),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_10),
.A2(n_74),
.B1(n_75),
.B2(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_10),
.B(n_84),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_149),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_10),
.A2(n_102),
.B1(n_103),
.B2(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_10),
.B(n_90),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_11),
.A2(n_74),
.B1(n_75),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_11),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_11),
.A2(n_62),
.B1(n_63),
.B2(n_158),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_158),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_11),
.A2(n_32),
.B1(n_35),
.B2(n_158),
.Y(n_237)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_13),
.A2(n_32),
.B1(n_35),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_13),
.A2(n_39),
.B1(n_62),
.B2(n_63),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_13),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_13),
.A2(n_39),
.B1(n_74),
.B2(n_75),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_14),
.A2(n_74),
.B1(n_75),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_14),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_14),
.A2(n_62),
.B1(n_63),
.B2(n_82),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_82),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_14),
.A2(n_32),
.B1(n_35),
.B2(n_82),
.Y(n_231)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_317),
.C(n_321),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_315),
.B(n_319),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_307),
.B(n_314),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_273),
.B(n_304),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_136),
.B(n_272),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_116),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_22),
.B(n_116),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_86),
.B2(n_115),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_23),
.B(n_87),
.C(n_99),
.Y(n_302)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_57),
.C(n_69),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_25),
.A2(n_26),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_41),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_27),
.A2(n_28),
.B1(n_41),
.B2(n_42),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_36),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_29),
.A2(n_102),
.B(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_30),
.A2(n_40),
.B1(n_126),
.B2(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_30),
.A2(n_40),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_31),
.A2(n_40),
.B(n_128),
.Y(n_202)
);

CKINVDCx6p67_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_35),
.B1(n_51),
.B2(n_52),
.Y(n_53)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_35),
.B(n_52),
.C(n_149),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_35),
.B(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_36),
.A2(n_103),
.B(n_146),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_38),
.B(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_44),
.A2(n_53),
.B(n_95),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

OA22x2_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_46),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_SL g198 ( 
.A1(n_45),
.A2(n_59),
.B(n_199),
.C(n_201),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_45),
.B(n_221),
.Y(n_220)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

NOR3xp33_ASAP7_75t_L g201 ( 
.A(n_46),
.B(n_60),
.C(n_62),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_49),
.A2(n_55),
.B(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_49),
.A2(n_94),
.B(n_107),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_49),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_49),
.A2(n_54),
.B1(n_206),
.B2(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_49),
.A2(n_54),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_49),
.A2(n_54),
.B1(n_214),
.B2(n_224),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_49),
.A2(n_54),
.B(n_94),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_53),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_53),
.B(n_149),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_57),
.B(n_69),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_61),
.B(n_64),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_58),
.B(n_68),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_58),
.A2(n_153),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_63),
.B1(n_73),
.B2(n_78),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_62),
.A2(n_78),
.B(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

HAxp5_ASAP7_75t_SL g200 ( 
.A(n_63),
.B(n_149),
.CON(n_200),
.SN(n_200)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_64),
.B(n_154),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_65),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_65),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_65),
.A2(n_90),
.B1(n_152),
.B2(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_65),
.A2(n_90),
.B1(n_187),
.B2(n_200),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_65),
.A2(n_90),
.B(n_131),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_80),
.B(n_83),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_70),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_70),
.A2(n_79),
.B1(n_156),
.B2(n_159),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_70),
.A2(n_113),
.B(n_311),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_71),
.A2(n_81),
.B1(n_84),
.B2(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_71),
.A2(n_84),
.B1(n_157),
.B2(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_71),
.B(n_114),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_71),
.A2(n_84),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_71),
.A2(n_84),
.B(n_85),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_79),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_78),
.Y(n_72)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_79),
.A2(n_286),
.B(n_287),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_83),
.B(n_287),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_85),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_99),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_92),
.B(n_98),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_92),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_90),
.B(n_131),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_91),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_93),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_98),
.B(n_276),
.C(n_289),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g303 ( 
.A(n_98),
.B(n_276),
.CI(n_289),
.CON(n_303),
.SN(n_303)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_108),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g289 ( 
.A1(n_100),
.A2(n_101),
.B(n_110),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_101),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_105),
.B1(n_106),
.B2(n_109),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B(n_104),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_102),
.A2(n_103),
.B1(n_229),
.B2(n_237),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_103),
.B(n_149),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_122),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_121),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_122),
.B(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_130),
.C(n_133),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_129),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_133),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_132),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_134),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_266),
.B(n_271),
.Y(n_136)
);

AOI221xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_175),
.B1(n_191),
.B2(n_265),
.C(n_324),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_164),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_139),
.B(n_164),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_160),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_140),
.B(n_161),
.C(n_162),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_150),
.C(n_155),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_142),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_144),
.B1(n_147),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_150),
.B(n_155),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_153),
.B(n_154),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g280 ( 
.A1(n_153),
.A2(n_281),
.B(n_282),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.C(n_174),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_174),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.C(n_172),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_170),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_171),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_189),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_176),
.B(n_189),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.C(n_181),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_177),
.B(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_179),
.B(n_181),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.C(n_185),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_185),
.B(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_264),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_259),
.B(n_263),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_215),
.B(n_258),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_210),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_195),
.B(n_210),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_207),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_203),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_197),
.B(n_203),
.C(n_207),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_198),
.B(n_202),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.C(n_213),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_213),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_253),
.B(n_257),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_243),
.B(n_252),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_232),
.B(n_242),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_227),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_227),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_219)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_220),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_225),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_238),
.B(n_241),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_240),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_245),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_248),
.C(n_251),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_256),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_262),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_301),
.Y(n_273)
);

AOI21xp33_ASAP7_75t_L g304 ( 
.A1(n_274),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_290),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_290),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_285),
.B2(n_288),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_283),
.B2(n_284),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_284),
.C(n_285),
.Y(n_291)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_284),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_294),
.C(n_299),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_285),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_285),
.A2(n_288),
.B1(n_293),
.B2(n_300),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_291),
.C(n_300),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_286),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_297),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_296),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_298),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_303),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_313),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_308),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_317),
.Y(n_320)
);

FAx1_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_310),
.CI(n_312),
.CON(n_308),
.SN(n_308)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_318),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);


endmodule