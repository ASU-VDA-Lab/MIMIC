module fake_jpeg_16116_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_0),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_16),
.Y(n_56)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_43),
.Y(n_49)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_17),
.B1(n_31),
.B2(n_19),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_61),
.B1(n_25),
.B2(n_20),
.Y(n_76)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_58),
.Y(n_83)
);

CKINVDCx6p67_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_63),
.Y(n_81)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_59),
.Y(n_93)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_35),
.A2(n_19),
.B1(n_16),
.B2(n_27),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_27),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_27),
.B1(n_22),
.B2(n_24),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_64),
.A2(n_68),
.B1(n_25),
.B2(n_20),
.Y(n_73)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_22),
.B1(n_20),
.B2(n_24),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_70),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_35),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_73),
.A2(n_0),
.B(n_1),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_78),
.B1(n_18),
.B2(n_32),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_53),
.B(n_35),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_24),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_22),
.B1(n_31),
.B2(n_17),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVxp67_ASAP7_75t_SL g108 ( 
.A(n_85),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_43),
.B1(n_39),
.B2(n_36),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_96)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_46),
.B(n_38),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_59),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_43),
.B1(n_39),
.B2(n_33),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_39),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_18),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_46),
.A2(n_36),
.B1(n_41),
.B2(n_34),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_55),
.A2(n_17),
.B1(n_31),
.B2(n_32),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVxp67_ASAP7_75t_SL g117 ( 
.A(n_94),
.Y(n_117)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_100),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_97),
.A2(n_106),
.B(n_118),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_47),
.B1(n_44),
.B2(n_66),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_98),
.A2(n_116),
.B1(n_79),
.B2(n_72),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_30),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_102),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_21),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_109),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_115),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_25),
.B(n_32),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_107),
.B(n_119),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_77),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_111),
.B1(n_29),
.B2(n_93),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_18),
.A3(n_29),
.B1(n_30),
.B2(n_41),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_21),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_112),
.B(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_44),
.B1(n_52),
.B2(n_58),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_81),
.B(n_87),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_82),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_93),
.Y(n_146)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_111),
.A2(n_89),
.B1(n_86),
.B2(n_52),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_128),
.A2(n_104),
.B1(n_28),
.B2(n_117),
.Y(n_171)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_80),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_130),
.A2(n_136),
.B(n_29),
.Y(n_167)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_132),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_96),
.A2(n_91),
.B1(n_82),
.B2(n_72),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_137),
.B1(n_139),
.B2(n_143),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_97),
.B(n_79),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_96),
.A2(n_71),
.B1(n_48),
.B2(n_42),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_113),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_145),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_114),
.A2(n_71),
.B1(n_41),
.B2(n_50),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_116),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_146),
.Y(n_158)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_114),
.A2(n_50),
.B1(n_93),
.B2(n_94),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_148),
.A2(n_95),
.B1(n_105),
.B2(n_115),
.Y(n_153)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_109),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_162),
.C(n_124),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_118),
.B(n_112),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_151),
.A2(n_152),
.B(n_165),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_140),
.A2(n_106),
.B(n_107),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_153),
.B(n_160),
.Y(n_201)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_146),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_103),
.C(n_59),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_126),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_0),
.B(n_1),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_138),
.B(n_130),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_171),
.A2(n_176),
.B1(n_131),
.B2(n_122),
.Y(n_189)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_175),
.Y(n_177)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_125),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_145),
.A2(n_104),
.B1(n_84),
.B2(n_85),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_168),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_178),
.B(n_184),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_182),
.C(n_183),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_134),
.Y(n_181)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_127),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_136),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_135),
.C(n_138),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_144),
.B1(n_128),
.B2(n_133),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_189),
.B1(n_192),
.B2(n_199),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_148),
.Y(n_190)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_143),
.C(n_132),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_198),
.C(n_200),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_168),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_195),
.A2(n_197),
.B(n_203),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_137),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_139),
.C(n_141),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_156),
.A2(n_142),
.B1(n_125),
.B2(n_131),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_166),
.C(n_165),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_122),
.Y(n_202)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_157),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_171),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_164),
.B1(n_154),
.B2(n_172),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_222),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_161),
.Y(n_206)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_200),
.A2(n_161),
.B1(n_174),
.B2(n_157),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_195),
.A2(n_155),
.B1(n_159),
.B2(n_170),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_153),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_203),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_167),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_220),
.C(n_223),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_197),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_23),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_193),
.A2(n_201),
.B(n_190),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_181),
.B(n_192),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_193),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_159),
.Y(n_221)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_163),
.B1(n_176),
.B2(n_84),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_202),
.Y(n_225)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_199),
.A2(n_30),
.B1(n_3),
.B2(n_4),
.Y(n_228)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_230),
.A2(n_215),
.B(n_216),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_185),
.Y(n_231)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_238),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_188),
.Y(n_233)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_198),
.C(n_188),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_240),
.C(n_243),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_187),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_189),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_242),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_196),
.C(n_191),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_196),
.C(n_191),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_30),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_247),
.C(n_21),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_21),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_221),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_206),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_249),
.B(n_224),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_235),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_258),
.Y(n_276)
);

XNOR2x2_ASAP7_75t_SL g254 ( 
.A(n_247),
.B(n_219),
.Y(n_254)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_263),
.C(n_239),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_207),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_262),
.C(n_267),
.Y(n_271)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_257),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_214),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

INVx13_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_250),
.B1(n_240),
.B2(n_4),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_218),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_264),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_229),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_211),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_236),
.A2(n_204),
.B1(n_216),
.B2(n_222),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_232),
.C(n_243),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_242),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_275),
.Y(n_289)
);

NOR2x1_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_204),
.Y(n_277)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_284),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_246),
.C(n_23),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_282),
.C(n_283),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_10),
.C(n_14),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_10),
.C(n_14),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_9),
.C(n_13),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_9),
.C(n_12),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_286),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_2),
.C(n_3),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_268),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_293),
.C(n_12),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_259),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_275),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_286),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_274),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_263),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_273),
.A2(n_253),
.B(n_255),
.Y(n_297)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_297),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_281),
.A2(n_261),
.B1(n_260),
.B2(n_270),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_298),
.A2(n_300),
.B1(n_12),
.B2(n_15),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_10),
.Y(n_299)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_277),
.A2(n_254),
.B1(n_8),
.B2(n_11),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_304),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_303),
.C(n_310),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_2),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_8),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_11),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_294),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_11),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_308),
.Y(n_315)
);

INVx6_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_294),
.Y(n_317)
);

NOR2x1_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_291),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_316),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_289),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_317),
.B(n_319),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_308),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_295),
.Y(n_319)
);

NAND4xp25_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_290),
.C(n_15),
.D(n_4),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_15),
.B(n_3),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_321),
.A2(n_323),
.B(n_324),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_318),
.B(n_302),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_313),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_2),
.C(n_5),
.Y(n_329)
);

AOI321xp33_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_312),
.A3(n_314),
.B1(n_315),
.B2(n_2),
.C(n_4),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_327),
.A2(n_329),
.B(n_326),
.Y(n_330)
);

NAND3xp33_ASAP7_75t_SL g331 ( 
.A(n_330),
.B(n_328),
.C(n_5),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_5),
.Y(n_333)
);


endmodule