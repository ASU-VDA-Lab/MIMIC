module real_aes_3016_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_453;
wire n_379;
wire n_374;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_504;
wire n_455;
wire n_231;
wire n_547;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_246;
wire n_412;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_613;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_498;
wire n_481;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_472;
wire n_452;
wire n_262;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_294;
wire n_393;
wire n_258;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_0), .A2(n_93), .B1(n_468), .B2(n_486), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_1), .A2(n_206), .B1(n_293), .B2(n_382), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_2), .A2(n_199), .B1(n_300), .B2(n_301), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_3), .A2(n_169), .B1(n_432), .B2(n_598), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_4), .A2(n_122), .B1(n_300), .B2(n_301), .Y(n_560) );
AO22x2_ASAP7_75t_L g243 ( .A1(n_5), .A2(n_158), .B1(n_240), .B2(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g576 ( .A(n_5), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_6), .A2(n_94), .B1(n_287), .B2(n_291), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_7), .A2(n_62), .B1(n_434), .B2(n_435), .Y(n_433) );
AOI221xp5_ASAP7_75t_SL g222 ( .A1(n_8), .A2(n_223), .B1(n_567), .B2(n_578), .C(n_584), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_9), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_10), .A2(n_69), .B1(n_341), .B2(n_344), .Y(n_340) );
AO22x2_ASAP7_75t_L g239 ( .A1(n_11), .A2(n_47), .B1(n_240), .B2(n_241), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_11), .B(n_575), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_12), .Y(n_551) );
AOI22xp33_ASAP7_75t_SL g427 ( .A1(n_13), .A2(n_149), .B1(n_313), .B2(n_428), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_14), .A2(n_121), .B1(n_265), .B2(n_426), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_15), .A2(n_180), .B1(n_297), .B2(n_298), .Y(n_296) );
AO222x2_ASAP7_75t_SL g520 ( .A1(n_16), .A2(n_32), .B1(n_130), .B2(n_237), .C1(n_253), .C2(n_258), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_17), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_18), .A2(n_102), .B1(n_438), .B2(n_439), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_19), .A2(n_219), .B1(n_366), .B2(n_421), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_20), .A2(n_135), .B1(n_509), .B2(n_512), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_21), .A2(n_48), .B1(n_336), .B2(n_339), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_22), .B(n_456), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_23), .A2(n_124), .B1(n_277), .B2(n_282), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_24), .A2(n_198), .B1(n_398), .B2(n_399), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_25), .A2(n_125), .B1(n_293), .B2(n_294), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_26), .A2(n_101), .B1(n_424), .B2(n_426), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_27), .A2(n_155), .B1(n_265), .B2(n_371), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_28), .A2(n_112), .B1(n_300), .B2(n_301), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_29), .A2(n_172), .B1(n_402), .B2(n_453), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_30), .A2(n_110), .B1(n_265), .B2(n_426), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_31), .A2(n_114), .B1(n_297), .B2(n_298), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_33), .A2(n_150), .B1(n_297), .B2(n_298), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_34), .A2(n_156), .B1(n_344), .B2(n_384), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_35), .A2(n_63), .B1(n_301), .B2(n_406), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_36), .A2(n_144), .B1(n_311), .B2(n_424), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_37), .A2(n_91), .B1(n_313), .B2(n_315), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_38), .A2(n_92), .B1(n_277), .B2(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_39), .A2(n_74), .B1(n_398), .B2(n_399), .Y(n_523) );
AOI22xp33_ASAP7_75t_SL g431 ( .A1(n_40), .A2(n_193), .B1(n_379), .B2(n_432), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_41), .A2(n_138), .B1(n_298), .B2(n_410), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_42), .A2(n_105), .B1(n_398), .B2(n_399), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_43), .A2(n_96), .B1(n_311), .B2(n_424), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_44), .A2(n_123), .B1(n_237), .B2(n_253), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_45), .A2(n_140), .B1(n_334), .B2(n_539), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_46), .A2(n_214), .B1(n_467), .B2(n_468), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_49), .A2(n_209), .B1(n_442), .B2(n_443), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_50), .A2(n_56), .B1(n_438), .B2(n_488), .Y(n_487) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_51), .A2(n_90), .B1(n_282), .B2(n_453), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_52), .A2(n_77), .B1(n_351), .B2(n_438), .Y(n_601) );
AO222x2_ASAP7_75t_SL g500 ( .A1(n_53), .A2(n_151), .B1(n_167), .B2(n_237), .C1(n_253), .C2(n_258), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_54), .A2(n_113), .B1(n_621), .B2(n_622), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_55), .A2(n_205), .B1(n_319), .B2(n_421), .Y(n_624) );
OA22x2_ASAP7_75t_L g231 ( .A1(n_57), .A2(n_232), .B1(n_233), .B2(n_303), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_57), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_58), .A2(n_98), .B1(n_432), .B2(n_464), .Y(n_463) );
INVx3_ASAP7_75t_L g240 ( .A(n_59), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_60), .A2(n_84), .B1(n_442), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_61), .A2(n_80), .B1(n_329), .B2(n_333), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_64), .A2(n_118), .B1(n_298), .B2(n_410), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_65), .A2(n_207), .B1(n_237), .B2(n_253), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_66), .A2(n_188), .B1(n_237), .B2(n_253), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_67), .A2(n_162), .B1(n_294), .B2(n_509), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_68), .A2(n_127), .B1(n_313), .B2(n_428), .Y(n_591) );
OAI22xp33_ASAP7_75t_L g306 ( .A1(n_70), .A2(n_307), .B1(n_352), .B2(n_353), .Y(n_306) );
INVx1_ASAP7_75t_L g352 ( .A(n_70), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_71), .A2(n_195), .B1(n_300), .B2(n_301), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_72), .A2(n_78), .B1(n_287), .B2(n_294), .Y(n_541) );
INVx1_ASAP7_75t_SL g248 ( .A(n_73), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_73), .B(n_109), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_75), .A2(n_202), .B1(n_333), .B2(n_378), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_76), .A2(n_97), .B1(n_277), .B2(n_402), .Y(n_547) );
INVx2_ASAP7_75t_L g583 ( .A(n_79), .Y(n_583) );
XOR2x2_ASAP7_75t_L g355 ( .A(n_81), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_82), .B(n_417), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_83), .A2(n_174), .B1(n_398), .B2(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_85), .A2(n_183), .B1(n_461), .B2(n_600), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_86), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_87), .A2(n_186), .B1(n_442), .B2(n_461), .Y(n_481) );
OA22x2_ASAP7_75t_L g610 ( .A1(n_88), .A2(n_611), .B1(n_612), .B2(n_613), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_88), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_89), .A2(n_117), .B1(n_310), .B2(n_311), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_95), .A2(n_194), .B1(n_321), .B2(n_366), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_99), .A2(n_159), .B1(n_293), .B2(n_294), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_100), .A2(n_210), .B1(n_336), .B2(n_376), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_103), .A2(n_212), .B1(n_365), .B2(n_367), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_104), .A2(n_160), .B1(n_348), .B2(n_381), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_106), .A2(n_141), .B1(n_464), .B2(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_107), .A2(n_192), .B1(n_313), .B2(n_315), .Y(n_625) );
AOI22xp33_ASAP7_75t_SL g626 ( .A1(n_108), .A2(n_189), .B1(n_310), .B2(n_311), .Y(n_626) );
AO22x2_ASAP7_75t_L g251 ( .A1(n_109), .A2(n_168), .B1(n_240), .B2(n_252), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_111), .A2(n_204), .B1(n_319), .B2(n_321), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_115), .A2(n_218), .B1(n_459), .B2(n_461), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_116), .A2(n_179), .B1(n_293), .B2(n_294), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_119), .A2(n_153), .B1(n_319), .B2(n_321), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_120), .A2(n_136), .B1(n_282), .B2(n_453), .Y(n_556) );
INVx1_ASAP7_75t_L g249 ( .A(n_126), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_128), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_129), .B(n_324), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_131), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_132), .B(n_417), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_133), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_134), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_137), .A2(n_154), .B1(n_420), .B2(n_421), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_139), .A2(n_181), .B1(n_359), .B2(n_361), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_142), .B(n_417), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_143), .B(n_324), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_145), .B(n_324), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_146), .A2(n_152), .B1(n_341), .B2(n_616), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_147), .A2(n_201), .B1(n_443), .B2(n_618), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_148), .A2(n_164), .B1(n_298), .B2(n_410), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_157), .A2(n_208), .B1(n_539), .B2(n_540), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_161), .A2(n_165), .B1(n_293), .B2(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_163), .A2(n_177), .B1(n_291), .B2(n_543), .Y(n_542) );
OA22x2_ASAP7_75t_L g448 ( .A1(n_166), .A2(n_449), .B1(n_469), .B2(n_470), .Y(n_448) );
INVx1_ASAP7_75t_L g469 ( .A(n_166), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_170), .A2(n_221), .B1(n_348), .B2(n_350), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_171), .A2(n_203), .B1(n_313), .B2(n_428), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_173), .B(n_363), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_175), .A2(n_216), .B1(n_287), .B2(n_294), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_176), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g571 ( .A(n_178), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_178), .B(n_583), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_182), .A2(n_187), .B1(n_287), .B2(n_382), .Y(n_562) );
INVx1_ASAP7_75t_L g572 ( .A(n_184), .Y(n_572) );
AND2x2_ASAP7_75t_R g604 ( .A(n_184), .B(n_571), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_185), .B(n_257), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_190), .A2(n_215), .B1(n_319), .B2(n_421), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_191), .B(n_582), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_196), .Y(n_280) );
AOI22x1_ASAP7_75t_SL g472 ( .A1(n_197), .A2(n_473), .B1(n_474), .B2(n_489), .Y(n_472) );
INVx1_ASAP7_75t_L g489 ( .A(n_197), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_200), .A2(n_217), .B1(n_298), .B2(n_410), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_211), .A2(n_586), .B1(n_587), .B2(n_602), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g602 ( .A(n_211), .Y(n_602) );
XOR2x2_ASAP7_75t_L g412 ( .A(n_213), .B(n_413), .Y(n_412) );
AOI22x1_ASAP7_75t_L g497 ( .A1(n_220), .A2(n_498), .B1(n_514), .B2(n_515), .Y(n_497) );
INVx1_ASAP7_75t_L g515 ( .A(n_220), .Y(n_515) );
OR2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_390), .Y(n_223) );
AOI21xp33_ASAP7_75t_L g567 ( .A1(n_224), .A2(n_390), .B(n_568), .Y(n_567) );
BUFx2_ASAP7_75t_SL g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
OAI22x1_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_354), .B1(n_387), .B2(n_388), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_304), .Y(n_227) );
OA21x2_ASAP7_75t_L g387 ( .A1(n_228), .A2(n_304), .B(n_385), .Y(n_387) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g386 ( .A(n_231), .Y(n_386) );
INVx1_ASAP7_75t_L g303 ( .A(n_233), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_284), .Y(n_233) );
NOR3xp33_ASAP7_75t_L g234 ( .A(n_235), .B(n_262), .C(n_274), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_236), .B(n_256), .Y(n_235) );
AND2x4_ASAP7_75t_L g237 ( .A(n_238), .B(n_245), .Y(n_237) );
AND2x2_ASAP7_75t_L g277 ( .A(n_238), .B(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g291 ( .A(n_238), .B(n_290), .Y(n_291) );
AND2x4_ASAP7_75t_L g314 ( .A(n_238), .B(n_278), .Y(n_314) );
AND2x2_ASAP7_75t_L g320 ( .A(n_238), .B(n_245), .Y(n_320) );
AND2x2_ASAP7_75t_L g453 ( .A(n_238), .B(n_278), .Y(n_453) );
AND2x2_ASAP7_75t_L g512 ( .A(n_238), .B(n_290), .Y(n_512) );
AND2x4_ASAP7_75t_L g238 ( .A(n_239), .B(n_242), .Y(n_238) );
AND2x2_ASAP7_75t_L g255 ( .A(n_239), .B(n_243), .Y(n_255) );
INVx1_ASAP7_75t_L g261 ( .A(n_239), .Y(n_261) );
INVx1_ASAP7_75t_L g268 ( .A(n_239), .Y(n_268) );
INVx2_ASAP7_75t_L g241 ( .A(n_240), .Y(n_241) );
INVx1_ASAP7_75t_L g244 ( .A(n_240), .Y(n_244) );
OAI22x1_ASAP7_75t_L g246 ( .A1(n_240), .A2(n_247), .B1(n_248), .B2(n_249), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_240), .Y(n_247) );
INVx1_ASAP7_75t_L g252 ( .A(n_240), .Y(n_252) );
AND2x4_ASAP7_75t_L g260 ( .A(n_242), .B(n_261), .Y(n_260) );
INVxp67_ASAP7_75t_L g283 ( .A(n_242), .Y(n_283) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g267 ( .A(n_243), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g266 ( .A(n_245), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g297 ( .A(n_245), .B(n_260), .Y(n_297) );
AND2x4_ASAP7_75t_L g338 ( .A(n_245), .B(n_260), .Y(n_338) );
AND2x4_ASAP7_75t_L g398 ( .A(n_245), .B(n_267), .Y(n_398) );
AND2x2_ASAP7_75t_L g410 ( .A(n_245), .B(n_260), .Y(n_410) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_250), .Y(n_245) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_246), .Y(n_254) );
AND2x2_ASAP7_75t_L g259 ( .A(n_246), .B(n_251), .Y(n_259) );
INVx2_ASAP7_75t_L g279 ( .A(n_246), .Y(n_279) );
AND2x4_ASAP7_75t_L g290 ( .A(n_250), .B(n_279), .Y(n_290) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g278 ( .A(n_251), .B(n_279), .Y(n_278) );
BUFx2_ASAP7_75t_L g302 ( .A(n_251), .Y(n_302) );
AND2x2_ASAP7_75t_SL g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g322 ( .A(n_254), .B(n_255), .Y(n_322) );
AND2x4_ASAP7_75t_L g298 ( .A(n_255), .B(n_290), .Y(n_298) );
AND2x4_ASAP7_75t_L g301 ( .A(n_255), .B(n_302), .Y(n_301) );
AND2x4_ASAP7_75t_L g334 ( .A(n_255), .B(n_302), .Y(n_334) );
AND2x4_ASAP7_75t_L g351 ( .A(n_255), .B(n_290), .Y(n_351) );
BUFx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
AND2x4_ASAP7_75t_L g271 ( .A(n_259), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g282 ( .A(n_259), .B(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g317 ( .A(n_259), .B(n_283), .Y(n_317) );
AND2x2_ASAP7_75t_L g326 ( .A(n_259), .B(n_260), .Y(n_326) );
AND2x2_ASAP7_75t_L g399 ( .A(n_259), .B(n_272), .Y(n_399) );
AND2x2_ASAP7_75t_L g402 ( .A(n_259), .B(n_283), .Y(n_402) );
AND2x2_ASAP7_75t_L g504 ( .A(n_259), .B(n_272), .Y(n_504) );
AND2x4_ASAP7_75t_L g289 ( .A(n_260), .B(n_290), .Y(n_289) );
AND2x6_ASAP7_75t_L g293 ( .A(n_260), .B(n_278), .Y(n_293) );
AND2x2_ASAP7_75t_L g343 ( .A(n_260), .B(n_278), .Y(n_343) );
AND2x2_ASAP7_75t_L g509 ( .A(n_260), .B(n_290), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_264), .B1(n_269), .B2(n_270), .Y(n_262) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_266), .Y(n_310) );
INVx3_ASAP7_75t_L g425 ( .A(n_266), .Y(n_425) );
AND2x6_ASAP7_75t_L g294 ( .A(n_267), .B(n_290), .Y(n_294) );
AND2x2_ASAP7_75t_SL g300 ( .A(n_267), .B(n_278), .Y(n_300) );
AND2x2_ASAP7_75t_L g332 ( .A(n_267), .B(n_278), .Y(n_332) );
AND2x4_ASAP7_75t_L g346 ( .A(n_267), .B(n_290), .Y(n_346) );
AND2x2_ASAP7_75t_L g406 ( .A(n_267), .B(n_278), .Y(n_406) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_268), .Y(n_273) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
BUFx4f_ASAP7_75t_L g311 ( .A(n_271), .Y(n_311) );
INVx2_ASAP7_75t_L g373 ( .A(n_271), .Y(n_373) );
BUFx6f_ASAP7_75t_SL g426 ( .A(n_271), .Y(n_426) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B1(n_280), .B2(n_281), .Y(n_274) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVxp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_295), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_292), .Y(n_285) );
INVx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx4_ASAP7_75t_L g349 ( .A(n_288), .Y(n_349) );
INVx2_ASAP7_75t_SL g442 ( .A(n_288), .Y(n_442) );
INVx3_ASAP7_75t_SL g467 ( .A(n_288), .Y(n_467) );
INVx2_ASAP7_75t_SL g618 ( .A(n_288), .Y(n_618) );
INVx8_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx3_ASAP7_75t_L g339 ( .A(n_291), .Y(n_339) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_291), .Y(n_382) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_291), .Y(n_443) );
INVx2_ASAP7_75t_L g462 ( .A(n_291), .Y(n_462) );
INVx1_ASAP7_75t_L g460 ( .A(n_293), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_299), .Y(n_295) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_306), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g353 ( .A(n_307), .Y(n_353) );
NOR2xp67_ASAP7_75t_L g307 ( .A(n_308), .B(n_327), .Y(n_307) );
NAND4xp25_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .C(n_318), .D(n_323), .Y(n_308) );
BUFx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_314), .Y(n_360) );
INVx2_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g361 ( .A(n_316), .Y(n_361) );
INVx2_ASAP7_75t_L g428 ( .A(n_316), .Y(n_428) );
INVx6_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx5_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx3_ASAP7_75t_L g366 ( .A(n_320), .Y(n_366) );
BUFx3_ASAP7_75t_L g420 ( .A(n_320), .Y(n_420) );
BUFx12f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx3_ASAP7_75t_L g369 ( .A(n_322), .Y(n_369) );
BUFx2_ASAP7_75t_L g363 ( .A(n_324), .Y(n_363) );
INVx4_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
INVx4_ASAP7_75t_SL g417 ( .A(n_325), .Y(n_417) );
INVx3_ASAP7_75t_SL g456 ( .A(n_325), .Y(n_456) );
INVx6_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND4xp25_ASAP7_75t_L g327 ( .A(n_328), .B(n_335), .C(n_340), .D(n_347), .Y(n_327) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g379 ( .A(n_331), .Y(n_379) );
INVx1_ASAP7_75t_L g464 ( .A(n_331), .Y(n_464) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_332), .Y(n_539) );
BUFx3_ASAP7_75t_L g598 ( .A(n_332), .Y(n_598) );
BUFx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx2_ASAP7_75t_L g432 ( .A(n_334), .Y(n_432) );
INVx5_ASAP7_75t_SL g484 ( .A(n_334), .Y(n_484) );
BUFx3_ASAP7_75t_L g540 ( .A(n_334), .Y(n_540) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g621 ( .A(n_337), .Y(n_621) );
INVx6_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx3_ASAP7_75t_L g438 ( .A(n_338), .Y(n_438) );
INVx2_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_SL g384 ( .A(n_342), .Y(n_384) );
INVx2_ASAP7_75t_L g434 ( .A(n_342), .Y(n_434) );
INVx2_ASAP7_75t_L g600 ( .A(n_342), .Y(n_600) );
INVx3_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g486 ( .A(n_343), .Y(n_486) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g435 ( .A(n_345), .Y(n_435) );
INVx2_ASAP7_75t_SL g468 ( .A(n_345), .Y(n_468) );
INVx2_ASAP7_75t_L g596 ( .A(n_345), .Y(n_596) );
INVx1_ASAP7_75t_SL g616 ( .A(n_345), .Y(n_616) );
INVx8_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
BUFx2_ASAP7_75t_SL g376 ( .A(n_351), .Y(n_376) );
INVx2_ASAP7_75t_L g440 ( .A(n_351), .Y(n_440) );
BUFx3_ASAP7_75t_L g488 ( .A(n_351), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_385), .Y(n_354) );
INVx5_ASAP7_75t_L g389 ( .A(n_355), .Y(n_389) );
NOR2x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_374), .Y(n_356) );
NAND4xp25_ASAP7_75t_L g357 ( .A(n_358), .B(n_362), .C(n_364), .D(n_370), .Y(n_357) );
BUFx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx6f_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g421 ( .A(n_369), .Y(n_421) );
INVx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND4xp25_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .C(n_380), .D(n_383), .Y(n_374) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
XNOR2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_494), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_393), .B1(n_444), .B2(n_445), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
XNOR2x1_ASAP7_75t_L g393 ( .A(n_394), .B(n_412), .Y(n_393) );
XNOR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_411), .Y(n_394) );
NOR2x1_ASAP7_75t_L g395 ( .A(n_396), .B(n_404), .Y(n_395) );
NAND4xp25_ASAP7_75t_L g396 ( .A(n_397), .B(n_400), .C(n_401), .D(n_403), .Y(n_396) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .C(n_408), .D(n_409), .Y(n_404) );
NAND2x1_ASAP7_75t_L g413 ( .A(n_414), .B(n_429), .Y(n_413) );
NOR2x1_ASAP7_75t_L g414 ( .A(n_415), .B(n_422), .Y(n_414) );
OAI21xp5_ASAP7_75t_SL g415 ( .A1(n_416), .A2(n_418), .B(n_419), .Y(n_415) );
INVx1_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_427), .Y(n_422) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NOR2x1_ASAP7_75t_L g429 ( .A(n_430), .B(n_436), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_433), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_441), .Y(n_436) );
INVx2_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_SL g622 ( .A(n_440), .Y(n_622) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_471), .B1(n_490), .B2(n_493), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g492 ( .A(n_447), .Y(n_492) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g470 ( .A(n_449), .Y(n_470) );
NOR2x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_457), .Y(n_449) );
NAND4xp25_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .C(n_454), .D(n_455), .Y(n_450) );
NAND4xp25_ASAP7_75t_L g457 ( .A(n_458), .B(n_463), .C(n_465), .D(n_466), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g543 ( .A(n_460), .Y(n_543) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g493 ( .A(n_471), .Y(n_493) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_480), .Y(n_474) );
NAND4xp25_ASAP7_75t_SL g475 ( .A(n_476), .B(n_477), .C(n_478), .D(n_479), .Y(n_475) );
NAND4xp25_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .C(n_485), .D(n_487), .Y(n_480) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AOI22xp33_ASAP7_75t_R g494 ( .A1(n_495), .A2(n_533), .B1(n_565), .B2(n_566), .Y(n_494) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g565 ( .A(n_496), .Y(n_565) );
AO22x2_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_516), .B1(n_517), .B2(n_532), .Y(n_496) );
INVx1_ASAP7_75t_L g532 ( .A(n_497), .Y(n_532) );
INVx1_ASAP7_75t_L g514 ( .A(n_498), .Y(n_514) );
NAND2x1_ASAP7_75t_SL g498 ( .A(n_499), .B(n_505), .Y(n_498) );
NOR2xp67_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
NOR2x1_ASAP7_75t_L g505 ( .A(n_506), .B(n_510), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_513), .Y(n_510) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
XOR2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_531), .Y(n_517) );
NAND2x1_ASAP7_75t_L g518 ( .A(n_519), .B(n_524), .Y(n_518) );
NOR2x1_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
NOR2x1_ASAP7_75t_L g524 ( .A(n_525), .B(n_528), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g566 ( .A(n_533), .Y(n_566) );
AO22x2_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_550), .B1(n_563), .B2(n_564), .Y(n_533) );
INVx1_ASAP7_75t_SL g563 ( .A(n_534), .Y(n_563) );
XNOR2x1_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_545), .Y(n_536) );
NAND4xp25_ASAP7_75t_L g537 ( .A(n_538), .B(n_541), .C(n_542), .D(n_544), .Y(n_537) );
NAND4xp25_ASAP7_75t_SL g545 ( .A(n_546), .B(n_547), .C(n_548), .D(n_549), .Y(n_545) );
INVx2_ASAP7_75t_SL g564 ( .A(n_550), .Y(n_564) );
XNOR2x1_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NOR2x1_ASAP7_75t_L g552 ( .A(n_553), .B(n_558), .Y(n_552) );
NAND4xp25_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .C(n_556), .D(n_557), .Y(n_553) );
NAND4xp25_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .C(n_561), .D(n_562), .Y(n_558) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_570), .B(n_574), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g580 ( .A(n_572), .Y(n_580) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_SL g578 ( .A(n_579), .B(n_581), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g628 ( .A(n_580), .B(n_581), .Y(n_628) );
OAI222xp33_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_603), .B1(n_605), .B2(n_610), .C1(n_611), .C2(n_628), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_587), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_594), .Y(n_588) );
NAND4xp25_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .C(n_592), .D(n_593), .Y(n_589) );
NAND4xp25_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .C(n_599), .D(n_601), .Y(n_594) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_606), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_607), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_608), .Y(n_607) );
CKINVDCx6p67_ASAP7_75t_R g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NOR2x1_ASAP7_75t_L g613 ( .A(n_614), .B(n_623), .Y(n_613) );
NAND4xp25_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .C(n_619), .D(n_620), .Y(n_614) );
NAND4xp25_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .C(n_626), .D(n_627), .Y(n_623) );
endmodule