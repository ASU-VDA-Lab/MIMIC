module real_jpeg_17536_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_578;
wire n_366;
wire n_149;
wire n_332;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_634;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_586;
wire n_405;
wire n_120;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_641;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_1),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_1),
.Y(n_126)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_1),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_2),
.Y(n_83)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_2),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_2),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_3),
.A2(n_117),
.B1(n_121),
.B2(n_122),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_3),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_3),
.A2(n_121),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_3),
.A2(n_101),
.B1(n_121),
.B2(n_351),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g573 ( 
.A1(n_3),
.A2(n_121),
.B1(n_148),
.B2(n_574),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_4),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_4),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g473 ( 
.A(n_4),
.Y(n_473)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_4),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_5),
.A2(n_21),
.B(n_23),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_6),
.Y(n_114)
);

BUFx4f_ASAP7_75t_L g120 ( 
.A(n_6),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_6),
.Y(n_131)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_6),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_7),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_147)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_7),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_7),
.A2(n_33),
.B1(n_152),
.B2(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_7),
.A2(n_152),
.B1(n_495),
.B2(n_496),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_7),
.A2(n_152),
.B1(n_535),
.B2(n_536),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_8),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_8),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_8),
.A2(n_157),
.B1(n_273),
.B2(n_275),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_8),
.A2(n_157),
.B1(n_380),
.B2(n_429),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_SL g516 ( 
.A1(n_8),
.A2(n_157),
.B1(n_312),
.B2(n_517),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_9),
.B(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_9),
.A2(n_89),
.B(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_9),
.Y(n_319)
);

OAI32xp33_ASAP7_75t_L g410 ( 
.A1(n_9),
.A2(n_411),
.A3(n_412),
.B1(n_415),
.B2(n_416),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_SL g436 ( 
.A1(n_9),
.A2(n_319),
.B1(n_437),
.B2(n_440),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_9),
.B(n_75),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_9),
.A2(n_107),
.B1(n_534),
.B2(n_540),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_10),
.A2(n_211),
.B1(n_213),
.B2(n_215),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_10),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_10),
.A2(n_215),
.B1(n_330),
.B2(n_334),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_10),
.A2(n_215),
.B1(n_263),
.B2(n_578),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_SL g617 ( 
.A1(n_10),
.A2(n_215),
.B1(n_618),
.B2(n_622),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_11),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_11),
.A2(n_69),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_11),
.A2(n_69),
.B1(n_346),
.B2(n_348),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_11),
.A2(n_69),
.B1(n_419),
.B2(n_422),
.Y(n_418)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_12),
.A2(n_33),
.B1(n_39),
.B2(n_40),
.Y(n_32)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_12),
.A2(n_39),
.B1(n_252),
.B2(n_255),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_12),
.A2(n_39),
.B1(n_384),
.B2(n_433),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_12),
.A2(n_39),
.B1(n_500),
.B2(n_503),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_14),
.A2(n_128),
.B1(n_132),
.B2(n_134),
.Y(n_127)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_14),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_14),
.A2(n_134),
.B1(n_181),
.B2(n_185),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_14),
.A2(n_134),
.B1(n_368),
.B2(n_373),
.Y(n_367)
);

OAI22xp33_ASAP7_75t_SL g585 ( 
.A1(n_14),
.A2(n_134),
.B1(n_586),
.B2(n_587),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_15),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_15),
.Y(n_189)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_15),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_15),
.Y(n_202)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_15),
.Y(n_237)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_15),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_15),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_16),
.A2(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_16),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_16),
.A2(n_227),
.B1(n_380),
.B2(n_384),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_16),
.A2(n_227),
.B1(n_373),
.B2(n_591),
.Y(n_590)
);

AO22x1_ASAP7_75t_L g630 ( 
.A1(n_16),
.A2(n_227),
.B1(n_631),
.B2(n_632),
.Y(n_630)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_17),
.A2(n_233),
.B1(n_238),
.B2(n_239),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_17),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_17),
.A2(n_238),
.B1(n_260),
.B2(n_263),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_17),
.A2(n_238),
.B1(n_309),
.B2(n_312),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_17),
.A2(n_238),
.B1(n_398),
.B2(n_400),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_19),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_19),
.Y(n_160)
);

BUFx8_ASAP7_75t_L g254 ( 
.A(n_19),
.Y(n_254)
);

BUFx12f_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_641),
.B(n_643),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_564),
.B(n_634),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_405),
.B(n_559),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_322),
.C(n_358),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_264),
.B(n_295),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_29),
.B(n_264),
.C(n_561),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_161),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_30),
.B(n_162),
.C(n_228),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_77),
.C(n_135),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_31),
.A2(n_135),
.B1(n_136),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_31),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_44),
.B1(n_67),
.B2(n_75),
.Y(n_31)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_32),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_37),
.Y(n_143)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_37),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_38),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx2_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_43),
.Y(n_414)
);

INVx3_ASAP7_75t_SL g258 ( 
.A(n_44),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_44),
.A2(n_75),
.B1(n_365),
.B2(n_366),
.Y(n_364)
);

OAI21xp33_ASAP7_75t_SL g613 ( 
.A1(n_44),
.A2(n_75),
.B(n_614),
.Y(n_613)
);

OA21x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_52),
.B(n_59),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_49),
.Y(n_439)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_51),
.Y(n_144)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_51),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_51),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_51),
.Y(n_375)
);

INVxp33_ASAP7_75t_L g416 ( 
.A(n_52),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_65),
.Y(n_288)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_67),
.Y(n_257)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_72),
.Y(n_263)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_76),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_76),
.A2(n_258),
.B1(n_272),
.B2(n_278),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_76),
.A2(n_258),
.B1(n_272),
.B2(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_76),
.A2(n_258),
.B1(n_259),
.B2(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_76),
.A2(n_258),
.B1(n_302),
.B2(n_436),
.Y(n_435)
);

OAI22x1_ASAP7_75t_L g576 ( 
.A1(n_76),
.A2(n_258),
.B1(n_367),
.B2(n_577),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_76),
.A2(n_258),
.B1(n_577),
.B2(n_590),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_77),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_106),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_78),
.B(n_106),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_88),
.B1(n_93),
.B2(n_100),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_86),
.Y(n_274)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_92),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_92),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_92),
.Y(n_347)
);

AO21x2_ASAP7_75t_SL g137 ( 
.A1(n_93),
.A2(n_138),
.B(n_142),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g399 ( 
.A(n_95),
.Y(n_399)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_95),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AO22x2_ASAP7_75t_L g142 ( 
.A1(n_98),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_142)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_104),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_104),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_115),
.B1(n_124),
.B2(n_127),
.Y(n_106)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_107),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_107),
.A2(n_127),
.B1(n_210),
.B2(n_246),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_107),
.A2(n_223),
.B(n_340),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_107),
.A2(n_499),
.B1(n_505),
.B2(n_506),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_107),
.A2(n_516),
.B1(n_531),
.B2(n_534),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_109),
.Y(n_317)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_110),
.Y(n_248)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_112),
.Y(n_224)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_113),
.Y(n_311)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_113),
.Y(n_502)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_114),
.Y(n_212)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_114),
.Y(n_214)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_114),
.Y(n_226)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_114),
.Y(n_539)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_116),
.A2(n_216),
.B1(n_308),
.B2(n_315),
.Y(n_307)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_120),
.Y(n_423)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_120),
.Y(n_468)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_126),
.Y(n_340)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_131),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_147),
.B1(n_153),
.B2(n_154),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_137),
.A2(n_153),
.B1(n_154),
.B2(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_137),
.A2(n_147),
.B1(n_153),
.B2(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_137),
.A2(n_153),
.B1(n_251),
.B2(n_345),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_137),
.A2(n_153),
.B1(n_345),
.B2(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_137),
.A2(n_153),
.B1(n_397),
.B2(n_573),
.Y(n_572)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_137),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_137),
.A2(n_153),
.B1(n_616),
.B2(n_617),
.Y(n_615)
);

OAI22xp33_ASAP7_75t_L g628 ( 
.A1(n_137),
.A2(n_153),
.B1(n_617),
.B2(n_629),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx6_ASAP7_75t_L g586 ( 
.A(n_140),
.Y(n_586)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_142),
.A2(n_583),
.B1(n_584),
.B2(n_585),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_SL g642 ( 
.A1(n_142),
.A2(n_584),
.B(n_630),
.Y(n_642)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_149),
.Y(n_255)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_150),
.Y(n_401)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_150),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_153),
.B(n_319),
.Y(n_318)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_155),
.Y(n_622)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_160),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_228),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_208),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_190),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_164),
.A2(n_190),
.B(n_208),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_179),
.Y(n_164)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_165),
.Y(n_244)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_165),
.Y(n_293)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_166),
.B(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_170),
.B1(n_174),
.B2(n_176),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_172),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_173),
.Y(n_314)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_174),
.Y(n_421)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_180),
.A2(n_285),
.B1(n_293),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_203),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_191),
.A2(n_203),
.B1(n_232),
.B2(n_243),
.Y(n_231)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_191),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_191),
.A2(n_377),
.B1(n_378),
.B2(n_379),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_191),
.A2(n_378),
.B1(n_428),
.B2(n_432),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_191),
.A2(n_243),
.B1(n_491),
.B2(n_494),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_191),
.A2(n_243),
.B1(n_428),
.B2(n_494),
.Y(n_510)
);

OA21x2_ASAP7_75t_L g570 ( 
.A1(n_191),
.A2(n_243),
.B(n_379),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_196),
.B1(n_199),
.B2(n_201),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_195),
.Y(n_337)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_201),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_202),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_202),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_206),
.B(n_319),
.Y(n_415)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_216),
.B1(n_217),
.B2(n_222),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_216),
.A2(n_308),
.B1(n_418),
.B2(n_424),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_216),
.A2(n_515),
.B1(n_520),
.B2(n_524),
.Y(n_514)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_SL g505 ( 
.A(n_219),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_219),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_221),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_249),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_229),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_245),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_230),
.A2(n_231),
.B1(n_245),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_232),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_235),
.Y(n_433)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_237),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_237),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_237),
.Y(n_383)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_239),
.Y(n_495)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_256),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_250),
.B(n_256),
.C(n_325),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_254),
.Y(n_575)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_254),
.Y(n_631)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_255),
.Y(n_587)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_261),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_262),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.C(n_270),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_265),
.B(n_321),
.Y(n_320)
);

XNOR2x1_ASAP7_75t_SL g321 ( 
.A(n_268),
.B(n_270),
.Y(n_321)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_279),
.C(n_284),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_284),
.Y(n_298)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_279),
.B(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_293),
.B2(n_294),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_285),
.A2(n_286),
.B1(n_293),
.B2(n_454),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_292),
.Y(n_431)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_293),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_R g543 ( 
.A(n_293),
.B(n_319),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_320),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_296),
.B(n_320),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.C(n_300),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_297),
.B(n_556),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_299),
.B(n_300),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_306),
.C(n_318),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_301),
.B(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_306),
.A2(n_307),
.B1(n_318),
.B2(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_311),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx5_ASAP7_75t_L g424 ( 
.A(n_316),
.Y(n_424)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_318),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_319),
.B(n_475),
.Y(n_474)
);

OAI21xp33_ASAP7_75t_SL g491 ( 
.A1(n_319),
.A2(n_474),
.B(n_492),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_319),
.B(n_531),
.Y(n_530)
);

A2O1A1O1Ixp25_ASAP7_75t_L g559 ( 
.A1(n_322),
.A2(n_358),
.B(n_560),
.C(n_562),
.D(n_563),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_357),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_323),
.B(n_357),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_326),
.Y(n_323)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_324),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_342),
.B1(n_355),
.B2(n_356),
.Y(n_326)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_327),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_327),
.B(n_356),
.C(n_404),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_328),
.A2(n_338),
.B1(n_339),
.B2(n_341),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_328),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_328),
.B(n_339),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_329),
.Y(n_377)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_333),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_338),
.A2(n_339),
.B1(n_395),
.B2(n_396),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_338),
.A2(n_396),
.B(n_402),
.Y(n_602)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_342),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_354),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_349),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_344),
.B(n_354),
.C(n_361),
.Y(n_360)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_349),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_350),
.Y(n_365)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_403),
.Y(n_358)
);

NOR2xp67_ASAP7_75t_L g563 ( 
.A(n_359),
.B(n_403),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_362),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_360),
.B(n_605),
.C(n_606),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_391),
.Y(n_362)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_363),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_364),
.A2(n_376),
.B(n_390),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_364),
.B(n_376),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_388),
.Y(n_464)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_390),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_390),
.A2(n_598),
.B1(n_601),
.B2(n_609),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_391),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_392),
.A2(n_393),
.B1(n_394),
.B2(n_402),
.Y(n_391)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_392),
.Y(n_402)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx3_ASAP7_75t_SL g400 ( 
.A(n_401),
.Y(n_400)
);

AOI21x1_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_554),
.B(n_558),
.Y(n_405)
);

OAI21x1_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_457),
.B(n_553),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_445),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_408),
.B(n_445),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_427),
.C(n_434),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_409),
.B(n_550),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_417),
.B1(n_425),
.B2(n_426),
.Y(n_409)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_410),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_410),
.B(n_426),
.Y(n_452)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_417),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_418),
.Y(n_506)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_419),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_427),
.A2(n_434),
.B1(n_435),
.B2(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_427),
.Y(n_551)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_431),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_432),
.Y(n_454)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx5_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_446),
.A2(n_447),
.B1(n_450),
.B2(n_451),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_446),
.B(n_453),
.C(n_455),
.Y(n_557)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_452),
.A2(n_453),
.B1(n_455),
.B2(n_456),
.Y(n_451)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_452),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_453),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_547),
.B(n_552),
.Y(n_457)
);

OAI21x1_ASAP7_75t_L g458 ( 
.A1(n_459),
.A2(n_512),
.B(n_546),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_497),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_460),
.B(n_497),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_489),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_461),
.A2(n_489),
.B1(n_490),
.B2(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_461),
.Y(n_526)
);

OAI32xp33_ASAP7_75t_L g461 ( 
.A1(n_462),
.A2(n_465),
.A3(n_469),
.B1(n_474),
.B2(n_477),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_466),
.B(n_530),
.Y(n_529)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_483),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_507),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_498),
.B(n_509),
.C(n_511),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_499),
.Y(n_524)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_508),
.A2(n_509),
.B1(n_510),
.B2(n_511),
.Y(n_507)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_508),
.Y(n_511)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_513),
.A2(n_527),
.B(n_545),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_525),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_514),
.B(n_525),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_528),
.A2(n_541),
.B(n_544),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_533),
.Y(n_528)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_532),
.Y(n_540)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_543),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_542),
.B(n_543),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_548),
.B(n_549),
.Y(n_547)
);

NOR2xp67_ASAP7_75t_SL g552 ( 
.A(n_548),
.B(n_549),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_555),
.B(n_557),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_555),
.B(n_557),
.Y(n_558)
);

NOR3xp33_ASAP7_75t_L g564 ( 
.A(n_565),
.B(n_610),
.C(n_626),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_566),
.B(n_603),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_567),
.A2(n_637),
.B(n_638),
.Y(n_636)
);

NOR2x1_ASAP7_75t_L g567 ( 
.A(n_568),
.B(n_597),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_568),
.B(n_597),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_569),
.B(n_580),
.Y(n_568)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_569),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_570),
.B(n_571),
.C(n_576),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_570),
.A2(n_589),
.B1(n_594),
.B2(n_595),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_570),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_570),
.B(n_576),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_570),
.B(n_582),
.C(n_595),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_571),
.A2(n_572),
.B1(n_581),
.B2(n_596),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_571),
.A2(n_572),
.B1(n_599),
.B2(n_600),
.Y(n_598)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_572),
.B(n_581),
.C(n_625),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_573),
.Y(n_583)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_581),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_582),
.B(n_588),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_585),
.Y(n_616)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_589),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_590),
.Y(n_614)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_598),
.B(n_601),
.C(n_602),
.Y(n_597)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_598),
.Y(n_609)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_599),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_602),
.B(n_608),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_604),
.B(n_607),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_604),
.B(n_607),
.Y(n_637)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

A2O1A1O1Ixp25_ASAP7_75t_L g635 ( 
.A1(n_611),
.A2(n_627),
.B(n_636),
.C(n_639),
.D(n_640),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_612),
.B(n_624),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_612),
.B(n_624),
.Y(n_639)
);

BUFx24_ASAP7_75t_SL g646 ( 
.A(n_612),
.Y(n_646)
);

FAx1_ASAP7_75t_SL g612 ( 
.A(n_613),
.B(n_615),
.CI(n_623),
.CON(n_612),
.SN(n_612)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_613),
.B(n_615),
.C(n_623),
.Y(n_633)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_628),
.B(n_633),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_628),
.B(n_633),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_628),
.B(n_642),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_628),
.B(n_642),
.Y(n_644)
);

CKINVDCx6p67_ASAP7_75t_R g629 ( 
.A(n_630),
.Y(n_629)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_635),
.Y(n_634)
);

CKINVDCx14_ASAP7_75t_R g643 ( 
.A(n_644),
.Y(n_643)
);


endmodule