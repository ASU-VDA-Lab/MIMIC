module fake_jpeg_5240_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_SL g10 ( 
.A(n_8),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_7),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_14),
.B(n_18),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_14),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_16),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_19),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_10),
.B1(n_19),
.B2(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_24),
.C(n_23),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_41),
.C(n_48),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_33),
.A2(n_35),
.B(n_32),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_47),
.B(n_14),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_17),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_18),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_28),
.C(n_15),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_46),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_27),
.B1(n_13),
.B2(n_21),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_53),
.B1(n_38),
.B2(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_54),
.B(n_56),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_56),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_60),
.B1(n_49),
.B2(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_57),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_40),
.B1(n_42),
.B2(n_27),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_22),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_54),
.C(n_22),
.Y(n_65)
);

INVxp33_ASAP7_75t_SL g63 ( 
.A(n_60),
.Y(n_63)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_66),
.B1(n_67),
.B2(n_10),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_62),
.C(n_61),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_4),
.C(n_5),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_70),
.B(n_3),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_63),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_73),
.C(n_4),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_71),
.C(n_6),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_74),
.Y(n_77)
);


endmodule