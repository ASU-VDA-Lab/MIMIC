module fake_jpeg_574_n_158 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_26),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_13),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_1),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_62),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_1),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_63),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_60),
.A2(n_53),
.B1(n_41),
.B2(n_52),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_49),
.B1(n_54),
.B2(n_61),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_51),
.B1(n_41),
.B2(n_54),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_70),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_60),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_65),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_78),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_51),
.B(n_63),
.C(n_42),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_79),
.A2(n_19),
.B1(n_37),
.B2(n_36),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_68),
.A2(n_49),
.B1(n_48),
.B2(n_45),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_83),
.B1(n_3),
.B2(n_4),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_47),
.B1(n_43),
.B2(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_48),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_89),
.Y(n_99)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_49),
.B1(n_45),
.B2(n_4),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_74),
.B1(n_65),
.B2(n_72),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_2),
.Y(n_89)
);

OAI32xp33_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_87),
.A3(n_76),
.B1(n_82),
.B2(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_27),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_70),
.C(n_74),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_101),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

NAND2x1_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_72),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_106),
.B(n_9),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_98),
.B(n_102),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_3),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_39),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_104),
.B(n_105),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_5),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_5),
.B(n_8),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_111),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_34),
.B(n_31),
.C(n_29),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_115),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_8),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_118),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_122),
.B(n_13),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_100),
.B1(n_103),
.B2(n_96),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_28),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_123),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_10),
.B(n_11),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_12),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_94),
.C(n_24),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_126),
.C(n_133),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_12),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_128),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_23),
.C(n_22),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_18),
.C(n_15),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_119),
.B1(n_120),
.B2(n_117),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_137),
.A2(n_132),
.B1(n_122),
.B2(n_127),
.Y(n_144)
);

XNOR2x1_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_111),
.Y(n_141)
);

OA21x2_ASAP7_75t_SL g146 ( 
.A1(n_141),
.A2(n_143),
.B(n_121),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_135),
.B(n_113),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_139),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_140),
.A2(n_132),
.B1(n_118),
.B2(n_130),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_143),
.C(n_141),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_136),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_149),
.C(n_150),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_144),
.B(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_145),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_152),
.B(n_146),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_153),
.A2(n_142),
.B(n_15),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_154),
.A2(n_14),
.B(n_16),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_14),
.B(n_16),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_17),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_17),
.Y(n_158)
);


endmodule