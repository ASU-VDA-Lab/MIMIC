module fake_jpeg_14057_n_232 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_42),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_50),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_46),
.B(n_31),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_23),
.B(n_21),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

NAND2x1_ASAP7_75t_SL g51 ( 
.A(n_17),
.B(n_0),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_0),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_56),
.Y(n_89)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_64),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_20),
.B1(n_26),
.B2(n_32),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_60),
.A2(n_76),
.B1(n_80),
.B2(n_83),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_71),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_36),
.A2(n_20),
.B1(n_26),
.B2(n_32),
.Y(n_76)
);

BUFx4f_ASAP7_75t_SL g77 ( 
.A(n_39),
.Y(n_77)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_81),
.Y(n_99)
);

AOI22x1_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_26),
.B1(n_27),
.B2(n_17),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_2),
.C(n_4),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_36),
.A2(n_20),
.B1(n_32),
.B2(n_38),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_41),
.B(n_31),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_92),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_42),
.A2(n_27),
.B1(n_22),
.B2(n_30),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_53),
.A2(n_22),
.B1(n_29),
.B2(n_24),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_88),
.B1(n_44),
.B2(n_3),
.Y(n_114)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_43),
.A2(n_30),
.B1(n_29),
.B2(n_24),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_23),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_2),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_68),
.B(n_19),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_95),
.B(n_118),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_19),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_56),
.Y(n_100)
);

OR2x2_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_52),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_57),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_107),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_80),
.B1(n_73),
.B2(n_76),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_1),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_62),
.B(n_12),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_108),
.B(n_109),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_88),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_2),
.B(n_3),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_114),
.B(n_63),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_73),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_4),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_67),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_120),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_77),
.B(n_11),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_5),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_6),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_122),
.A2(n_141),
.B1(n_119),
.B2(n_111),
.Y(n_160)
);

OAI32xp33_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_69),
.A3(n_60),
.B1(n_70),
.B2(n_67),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_130),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_95),
.B(n_77),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_134),
.C(n_135),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_129),
.A2(n_137),
.B(n_97),
.Y(n_165)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_146),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_11),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_133),
.B(n_145),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_91),
.C(n_72),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_66),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_84),
.B1(n_66),
.B2(n_72),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_SL g139 ( 
.A(n_103),
.B(n_6),
.C(n_7),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_SL g159 ( 
.A(n_139),
.B(n_101),
.C(n_120),
.Y(n_159)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_110),
.A2(n_84),
.B1(n_65),
.B2(n_91),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_118),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_99),
.B(n_7),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_7),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_103),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_164),
.C(n_124),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_112),
.B(n_96),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_150),
.B(n_161),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_101),
.B(n_98),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_144),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_162),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_149),
.B(n_139),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_122),
.B1(n_141),
.B2(n_137),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_102),
.B(n_115),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_108),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g163 ( 
.A(n_135),
.B(n_121),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_166),
.B(n_131),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_117),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_97),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_102),
.B(n_97),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_130),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_106),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_125),
.B1(n_143),
.B2(n_134),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_176),
.Y(n_189)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_174),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_171),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_182),
.C(n_185),
.Y(n_197)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_124),
.C(n_127),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_175),
.A2(n_155),
.B(n_159),
.Y(n_192)
);

NAND2x1_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_130),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_165),
.B(n_163),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_178),
.B(n_147),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_154),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_153),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_70),
.B1(n_75),
.B2(n_117),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_168),
.Y(n_196)
);

NOR3xp33_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_184),
.C(n_148),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_140),
.C(n_138),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_75),
.C(n_65),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_190),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_183),
.B(n_158),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_173),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_177),
.C(n_181),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_194),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_155),
.B(n_163),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_196),
.Y(n_201)
);

OA21x2_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_148),
.B(n_168),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_180),
.Y(n_202)
);

AO21x1_ASAP7_75t_L g214 ( 
.A1(n_202),
.A2(n_207),
.B(n_191),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_179),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_192),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_173),
.B1(n_170),
.B2(n_176),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_204),
.B(n_195),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_197),
.B(n_172),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_206),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_199),
.A2(n_198),
.B(n_189),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_212),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_197),
.C(n_182),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_210),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_185),
.C(n_189),
.Y(n_210)
);

AOI21x1_ASAP7_75t_SL g218 ( 
.A1(n_211),
.A2(n_214),
.B(n_201),
.Y(n_218)
);

INVx11_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_219),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_220),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_157),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_206),
.Y(n_220)
);

AOI21x1_ASAP7_75t_L g221 ( 
.A1(n_215),
.A2(n_177),
.B(n_207),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_221),
.A2(n_218),
.B(n_216),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_198),
.B1(n_196),
.B2(n_164),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_223),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_223),
.Y(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_227),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_217),
.C(n_220),
.Y(n_230)
);

OAI31xp33_ASAP7_75t_L g231 ( 
.A1(n_230),
.A2(n_229),
.A3(n_220),
.B(n_156),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_9),
.C(n_199),
.Y(n_232)
);


endmodule