module fake_jpeg_20493_n_120 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_17),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_1),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_60),
.Y(n_64)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_62),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_46),
.B(n_2),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_43),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_49),
.B1(n_42),
.B2(n_44),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_71),
.B1(n_76),
.B2(n_43),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_52),
.B1(n_49),
.B2(n_45),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVxp67_ASAP7_75t_SL g78 ( 
.A(n_72),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_85),
.Y(n_93)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_84),
.Y(n_97)
);

AO22x1_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_47),
.B1(n_53),
.B2(n_55),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_90),
.B1(n_3),
.B2(n_4),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_53),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_54),
.B1(n_48),
.B2(n_24),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_89),
.A2(n_22),
.B1(n_37),
.B2(n_36),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_95),
.B1(n_98),
.B2(n_100),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_82),
.A2(n_18),
.B1(n_35),
.B2(n_34),
.Y(n_95)
);

NAND2xp67_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_5),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_16),
.B(n_33),
.C(n_31),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_99),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_106),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_83),
.B(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_107),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_79),
.C(n_90),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_96),
.C(n_100),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_94),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_108),
.C(n_105),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_104),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_112),
.C(n_105),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_101),
.C(n_107),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_98),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_115),
.A2(n_99),
.B1(n_23),
.B2(n_26),
.Y(n_116)
);

OAI321xp33_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_13),
.A3(n_30),
.B1(n_29),
.B2(n_28),
.C(n_11),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

AOI321xp33_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_12),
.A3(n_27),
.B1(n_38),
.B2(n_9),
.C(n_6),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_6),
.C(n_7),
.Y(n_120)
);


endmodule