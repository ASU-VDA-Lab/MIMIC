module fake_jpeg_10298_n_46 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_46);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_32;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_12),
.A2(n_10),
.B1(n_17),
.B2(n_3),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_0),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_5),
.B(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVxp33_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_2),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_23),
.B1(n_19),
.B2(n_7),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_34),
.C(n_36),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_19),
.B1(n_6),
.B2(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_33),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_40),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_35),
.C(n_42),
.Y(n_45)
);

AOI321xp33_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_43),
.A3(n_37),
.B1(n_41),
.B2(n_13),
.C(n_16),
.Y(n_46)
);


endmodule