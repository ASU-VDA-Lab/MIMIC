module fake_jpeg_24192_n_277 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx8_ASAP7_75t_SL g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVxp33_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_32),
.B1(n_28),
.B2(n_16),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_16),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_22),
.B1(n_24),
.B2(n_30),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_49),
.B(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_55),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_32),
.B1(n_28),
.B2(n_22),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_58),
.B1(n_16),
.B2(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_20),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_22),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_60),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_16),
.B1(n_22),
.B2(n_24),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_31),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_34),
.B(n_17),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_17),
.B(n_23),
.C(n_27),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_66),
.B(n_30),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_82),
.Y(n_98)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_84),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_62),
.B1(n_64),
.B2(n_52),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_57),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_76),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_37),
.B(n_40),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_50),
.C(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_37),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_18),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_27),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_40),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_44),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_62),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_87),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_88),
.Y(n_99)
);

XNOR2x1_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_59),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_92),
.C(n_96),
.Y(n_126)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_59),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_62),
.B1(n_47),
.B2(n_46),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_80),
.B1(n_74),
.B2(n_86),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_73),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_106),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_107),
.B1(n_84),
.B2(n_54),
.Y(n_128)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_45),
.B1(n_52),
.B2(n_47),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_81),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_55),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_82),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_117),
.B1(n_124),
.B2(n_93),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_104),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_116),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_69),
.B1(n_45),
.B2(n_67),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_87),
.B(n_75),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_137),
.B(n_134),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_73),
.B(n_85),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_137),
.B(n_21),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_90),
.A2(n_45),
.B1(n_47),
.B2(n_81),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_106),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_128),
.A2(n_132),
.B1(n_101),
.B2(n_95),
.Y(n_141)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_135),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_61),
.C(n_49),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_134),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_84),
.B1(n_75),
.B2(n_54),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_59),
.C(n_82),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_96),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_111),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_92),
.A2(n_26),
.B(n_20),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_153),
.C(n_129),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_91),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_146),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_141),
.B1(n_147),
.B2(n_149),
.Y(n_173)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_154),
.B(n_125),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_94),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_98),
.B1(n_108),
.B2(n_83),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_115),
.B(n_109),
.Y(n_150)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_161),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_136),
.A2(n_126),
.B(n_135),
.C(n_115),
.D(n_113),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_98),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_121),
.B(n_78),
.Y(n_155)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_121),
.B(n_98),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_157),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_78),
.B1(n_21),
.B2(n_26),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_83),
.B1(n_103),
.B2(n_44),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_159),
.A2(n_112),
.B1(n_19),
.B2(n_17),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_128),
.A2(n_29),
.B1(n_19),
.B2(n_23),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_160),
.A2(n_164),
.B1(n_120),
.B2(n_29),
.Y(n_177)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_163),
.B(n_17),
.Y(n_180)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_162),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_175),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_168),
.B(n_186),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_126),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_171),
.C(n_181),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_118),
.B(n_114),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_129),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_7),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_156),
.Y(n_175)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_51),
.B(n_118),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_SL g207 ( 
.A(n_176),
.B(n_180),
.C(n_182),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_158),
.B1(n_159),
.B2(n_149),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_163),
.Y(n_181)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_23),
.A3(n_17),
.B1(n_0),
.B2(n_1),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_164),
.B1(n_172),
.B2(n_179),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_112),
.B(n_1),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_185),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_190),
.Y(n_211)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_196),
.B1(n_197),
.B2(n_202),
.Y(n_214)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_140),
.B1(n_145),
.B2(n_142),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_194),
.A2(n_206),
.B1(n_186),
.B2(n_182),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_151),
.B1(n_161),
.B2(n_145),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_184),
.A2(n_148),
.B1(n_139),
.B2(n_153),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_146),
.C(n_112),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_171),
.C(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_201),
.Y(n_212)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_166),
.A2(n_184),
.B1(n_172),
.B2(n_168),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_188),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_208),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_176),
.A2(n_186),
.B1(n_174),
.B2(n_180),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_169),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_7),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_207),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_210),
.A2(n_216),
.B1(n_226),
.B2(n_15),
.Y(n_239)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_207),
.B(n_203),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_217),
.B(n_221),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_219),
.C(n_204),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_181),
.C(n_178),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_223),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_192),
.B(n_176),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_205),
.B(n_199),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_225),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_7),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_0),
.B(n_1),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_224),
.A2(n_191),
.B(n_198),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_0),
.B(n_1),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_197),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_210),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_228),
.A2(n_239),
.B1(n_226),
.B2(n_216),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_196),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_231),
.B(n_232),
.Y(n_245)
);

BUFx12_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_233),
.A2(n_216),
.B(n_210),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_219),
.C(n_218),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_2),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_236),
.B(n_237),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_2),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_244),
.Y(n_256)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_242),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_229),
.C(n_232),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_223),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_2),
.C(n_3),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_230),
.C(n_5),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_249),
.B(n_4),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_252),
.C(n_253),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_232),
.C(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_245),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_4),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_247),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_246),
.Y(n_258)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_258),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_251),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_248),
.B1(n_240),
.B2(n_244),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_256),
.C(n_9),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_247),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_263),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_265),
.C(n_266),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_260),
.A2(n_256),
.B(n_9),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_267),
.A2(n_263),
.B(n_10),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_270),
.Y(n_273)
);

A2O1A1O1Ixp25_ASAP7_75t_L g271 ( 
.A1(n_268),
.A2(n_5),
.B(n_10),
.C(n_12),
.D(n_13),
.Y(n_271)
);

A2O1A1O1Ixp25_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_268),
.B(n_269),
.C(n_15),
.D(n_13),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_273),
.C(n_14),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_275),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_14),
.Y(n_277)
);


endmodule