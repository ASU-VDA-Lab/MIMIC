module real_aes_2332_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_769;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g539 ( .A(n_0), .B(n_160), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_1), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_2), .B(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g118 ( .A(n_3), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_4), .B(n_501), .Y(n_500) );
NAND2xp33_ASAP7_75t_SL g582 ( .A(n_5), .B(n_147), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_6), .B(n_127), .Y(n_151) );
INVx1_ASAP7_75t_L g575 ( .A(n_7), .Y(n_575) );
INVx1_ASAP7_75t_L g173 ( .A(n_8), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g791 ( .A(n_9), .Y(n_791) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_10), .Y(n_189) );
AND2x2_ASAP7_75t_L g498 ( .A(n_11), .B(n_204), .Y(n_498) );
INVx2_ASAP7_75t_L g126 ( .A(n_12), .Y(n_126) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_13), .Y(n_486) );
INVx1_ASAP7_75t_L g161 ( .A(n_14), .Y(n_161) );
AOI221x1_ASAP7_75t_L g578 ( .A1(n_15), .A2(n_178), .B1(n_503), .B2(n_579), .C(n_581), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_16), .B(n_501), .Y(n_562) );
INVx1_ASAP7_75t_L g489 ( .A(n_17), .Y(n_489) );
INVx1_ASAP7_75t_L g158 ( .A(n_18), .Y(n_158) );
INVx1_ASAP7_75t_SL g233 ( .A(n_19), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_20), .B(n_138), .Y(n_137) );
AOI33xp33_ASAP7_75t_L g210 ( .A1(n_21), .A2(n_49), .A3(n_115), .B1(n_133), .B2(n_211), .B3(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_22), .A2(n_503), .B(n_504), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_23), .B(n_160), .Y(n_505) );
AOI221xp5_ASAP7_75t_SL g549 ( .A1(n_24), .A2(n_39), .B1(n_501), .B2(n_503), .C(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g182 ( .A(n_25), .Y(n_182) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_26), .A2(n_88), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g128 ( .A(n_26), .B(n_88), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_27), .B(n_163), .Y(n_566) );
INVxp67_ASAP7_75t_L g577 ( .A(n_28), .Y(n_577) );
AND2x2_ASAP7_75t_L g524 ( .A(n_29), .B(n_203), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_30), .B(n_171), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_31), .A2(n_503), .B(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_32), .B(n_163), .Y(n_551) );
AND2x2_ASAP7_75t_L g121 ( .A(n_33), .B(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g132 ( .A(n_33), .Y(n_132) );
AND2x2_ASAP7_75t_L g147 ( .A(n_33), .B(n_118), .Y(n_147) );
OR2x6_ASAP7_75t_L g487 ( .A(n_34), .B(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_35), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_36), .B(n_171), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g111 ( .A1(n_37), .A2(n_112), .B1(n_124), .B2(n_127), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_38), .B(n_144), .Y(n_143) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_40), .A2(n_79), .B1(n_130), .B2(n_503), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_41), .B(n_138), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_42), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_43), .B(n_160), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_44), .B(n_149), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_45), .B(n_138), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_46), .Y(n_123) );
AND2x2_ASAP7_75t_L g542 ( .A(n_47), .B(n_203), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_48), .B(n_203), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_50), .B(n_138), .Y(n_201) );
INVx1_ASAP7_75t_L g116 ( .A(n_51), .Y(n_116) );
INVx1_ASAP7_75t_L g140 ( .A(n_51), .Y(n_140) );
AND2x2_ASAP7_75t_L g202 ( .A(n_52), .B(n_203), .Y(n_202) );
AOI221xp5_ASAP7_75t_L g170 ( .A1(n_53), .A2(n_71), .B1(n_130), .B2(n_171), .C(n_172), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_54), .B(n_171), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_55), .B(n_501), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_56), .B(n_124), .Y(n_191) );
AOI21xp5_ASAP7_75t_SL g221 ( .A1(n_57), .A2(n_130), .B(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g515 ( .A(n_58), .B(n_203), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_59), .B(n_163), .Y(n_540) );
INVx1_ASAP7_75t_L g154 ( .A(n_60), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_61), .B(n_160), .Y(n_513) );
AND2x2_ASAP7_75t_SL g567 ( .A(n_62), .B(n_204), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_63), .A2(n_503), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g200 ( .A(n_64), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_65), .B(n_163), .Y(n_506) );
AND2x2_ASAP7_75t_SL g531 ( .A(n_66), .B(n_149), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_67), .A2(n_130), .B(n_199), .Y(n_198) );
AOI222xp33_ASAP7_75t_L g99 ( .A1(n_68), .A2(n_100), .B1(n_784), .B2(n_795), .C1(n_814), .C2(n_818), .Y(n_99) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_68), .A2(n_86), .B1(n_478), .B2(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_68), .Y(n_800) );
INVx1_ASAP7_75t_L g122 ( .A(n_69), .Y(n_122) );
INVx1_ASAP7_75t_L g142 ( .A(n_69), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_70), .B(n_171), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_72), .Y(n_807) );
AND2x2_ASAP7_75t_L g235 ( .A(n_73), .B(n_178), .Y(n_235) );
INVx1_ASAP7_75t_L g155 ( .A(n_74), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_75), .A2(n_130), .B(n_232), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g129 ( .A1(n_76), .A2(n_130), .B(n_136), .C(n_148), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_77), .B(n_501), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_78), .A2(n_82), .B1(n_171), .B2(n_501), .Y(n_529) );
INVx1_ASAP7_75t_L g490 ( .A(n_80), .Y(n_490) );
AND2x2_ASAP7_75t_SL g219 ( .A(n_81), .B(n_178), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_83), .A2(n_130), .B1(n_208), .B2(n_209), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_84), .B(n_160), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_85), .B(n_160), .Y(n_552) );
NOR3xp33_ASAP7_75t_L g104 ( .A(n_86), .B(n_105), .C(n_332), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_86), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_87), .A2(n_503), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g223 ( .A(n_89), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_90), .B(n_163), .Y(n_512) );
AND2x2_ASAP7_75t_L g214 ( .A(n_91), .B(n_178), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_92), .A2(n_180), .B(n_181), .C(n_183), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_93), .B(n_501), .Y(n_541) );
INVxp67_ASAP7_75t_L g580 ( .A(n_94), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_95), .B(n_163), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_96), .A2(n_503), .B(n_564), .Y(n_563) );
BUFx2_ASAP7_75t_L g792 ( .A(n_97), .Y(n_792) );
BUFx2_ASAP7_75t_SL g822 ( .A(n_97), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_98), .B(n_138), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_776), .B(n_777), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OAI22xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_482), .B1(n_491), .B2(n_772), .Y(n_102) );
AO22x2_ASAP7_75t_L g778 ( .A1(n_103), .A2(n_483), .B1(n_491), .B2(n_773), .Y(n_778) );
AOI211x1_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_374), .B(n_475), .C(n_479), .Y(n_103) );
INVxp67_ASAP7_75t_L g477 ( .A(n_105), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_105), .B(n_419), .Y(n_804) );
NAND3xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_279), .C(n_312), .Y(n_105) );
AOI211xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_236), .B(n_245), .C(n_269), .Y(n_106) );
OAI21xp33_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_165), .B(n_215), .Y(n_107) );
OR2x2_ASAP7_75t_L g289 ( .A(n_108), .B(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g417 ( .A(n_108), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g401 ( .A(n_109), .B(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_SL g421 ( .A1(n_109), .A2(n_422), .B1(n_425), .B2(n_426), .Y(n_421) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_150), .Y(n_109) );
INVx1_ASAP7_75t_L g268 ( .A(n_110), .Y(n_268) );
AND2x4_ASAP7_75t_L g285 ( .A(n_110), .B(n_266), .Y(n_285) );
INVx2_ASAP7_75t_L g307 ( .A(n_110), .Y(n_307) );
AND2x2_ASAP7_75t_L g355 ( .A(n_110), .B(n_218), .Y(n_355) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_110), .Y(n_369) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_129), .Y(n_110) );
NOR3xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_119), .C(n_123), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g171 ( .A(n_114), .B(n_120), .Y(n_171) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
OR2x6_ASAP7_75t_L g145 ( .A(n_115), .B(n_134), .Y(n_145) );
INVxp33_ASAP7_75t_L g211 ( .A(n_115), .Y(n_211) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g135 ( .A(n_116), .B(n_118), .Y(n_135) );
AND2x4_ASAP7_75t_L g163 ( .A(n_116), .B(n_141), .Y(n_163) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x6_ASAP7_75t_L g503 ( .A(n_121), .B(n_135), .Y(n_503) );
INVx2_ASAP7_75t_L g134 ( .A(n_122), .Y(n_134) );
AND2x6_ASAP7_75t_L g160 ( .A(n_122), .B(n_139), .Y(n_160) );
INVx4_ASAP7_75t_L g178 ( .A(n_124), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_124), .B(n_188), .Y(n_187) );
AOI21x1_ASAP7_75t_L g535 ( .A1(n_124), .A2(n_536), .B(n_542), .Y(n_535) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx4f_ASAP7_75t_L g149 ( .A(n_125), .Y(n_149) );
AND2x4_ASAP7_75t_L g127 ( .A(n_126), .B(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_SL g204 ( .A(n_126), .B(n_128), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_127), .B(n_146), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_127), .A2(n_221), .B(n_225), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_127), .A2(n_500), .B(n_502), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_127), .B(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_127), .B(n_577), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_127), .B(n_580), .Y(n_579) );
NOR3xp33_ASAP7_75t_L g581 ( .A(n_127), .B(n_156), .C(n_582), .Y(n_581) );
INVxp67_ASAP7_75t_L g190 ( .A(n_130), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_130), .A2(n_171), .B1(n_574), .B2(n_576), .Y(n_573) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_135), .Y(n_130) );
NOR2x1p5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
INVx1_ASAP7_75t_L g212 ( .A(n_133), .Y(n_212) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_143), .B(n_146), .Y(n_136) );
INVx1_ASAP7_75t_L g156 ( .A(n_138), .Y(n_156) );
AND2x4_ASAP7_75t_L g501 ( .A(n_138), .B(n_147), .Y(n_501) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OAI22xp5_ASAP7_75t_L g153 ( .A1(n_145), .A2(n_154), .B1(n_155), .B2(n_156), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_SL g172 ( .A1(n_145), .A2(n_146), .B(n_173), .C(n_174), .Y(n_172) );
INVxp67_ASAP7_75t_L g180 ( .A(n_145), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_145), .A2(n_146), .B(n_200), .C(n_201), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_145), .A2(n_146), .B(n_223), .C(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_SL g232 ( .A1(n_145), .A2(n_146), .B(n_233), .C(n_234), .Y(n_232) );
INVx1_ASAP7_75t_L g208 ( .A(n_146), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_146), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_146), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_146), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_146), .A2(n_539), .B(n_540), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_146), .A2(n_551), .B(n_552), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_146), .A2(n_565), .B(n_566), .Y(n_564) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_148), .A2(n_206), .B(n_214), .Y(n_205) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_148), .A2(n_206), .B(n_214), .Y(n_250) );
AOI21x1_ASAP7_75t_L g527 ( .A1(n_148), .A2(n_528), .B(n_531), .Y(n_527) );
INVx2_ASAP7_75t_SL g148 ( .A(n_149), .Y(n_148) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_149), .A2(n_170), .B(n_175), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_149), .A2(n_562), .B(n_563), .Y(n_561) );
AND2x2_ASAP7_75t_L g226 ( .A(n_150), .B(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g255 ( .A(n_150), .Y(n_255) );
INVx3_ASAP7_75t_L g266 ( .A(n_150), .Y(n_266) );
AND2x4_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
OAI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_157), .B(n_164), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_156), .B(n_182), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B1(n_161), .B2(n_162), .Y(n_157) );
INVxp67_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVxp67_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_165), .A2(n_350), .B1(n_352), .B2(n_354), .Y(n_349) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_165), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_193), .Y(n_166) );
INVx3_ASAP7_75t_L g239 ( .A(n_167), .Y(n_239) );
AND2x2_ASAP7_75t_L g247 ( .A(n_167), .B(n_248), .Y(n_247) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_167), .Y(n_277) );
NAND2x1_ASAP7_75t_SL g366 ( .A(n_167), .B(n_238), .Y(n_366) );
AND2x4_ASAP7_75t_L g167 ( .A(n_168), .B(n_176), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g244 ( .A(n_169), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_169), .B(n_250), .Y(n_262) );
AND2x2_ASAP7_75t_L g275 ( .A(n_169), .B(n_176), .Y(n_275) );
AND2x4_ASAP7_75t_L g282 ( .A(n_169), .B(n_283), .Y(n_282) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_169), .Y(n_331) );
INVx1_ASAP7_75t_L g341 ( .A(n_169), .Y(n_341) );
INVxp67_ASAP7_75t_L g424 ( .A(n_169), .Y(n_424) );
INVx1_ASAP7_75t_L g192 ( .A(n_171), .Y(n_192) );
INVx1_ASAP7_75t_L g242 ( .A(n_176), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_176), .B(n_252), .Y(n_261) );
INVx2_ASAP7_75t_L g329 ( .A(n_176), .Y(n_329) );
INVx1_ASAP7_75t_L g372 ( .A(n_176), .Y(n_372) );
OR2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_186), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B1(n_184), .B2(n_185), .Y(n_177) );
INVx3_ASAP7_75t_L g185 ( .A(n_178), .Y(n_185) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_185), .A2(n_196), .B(n_202), .Y(n_195) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_185), .A2(n_196), .B(n_202), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_190), .B1(n_191), .B2(n_192), .Y(n_186) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g298 ( .A(n_193), .B(n_275), .Y(n_298) );
AND2x2_ASAP7_75t_L g447 ( .A(n_193), .B(n_371), .Y(n_447) );
AND2x2_ASAP7_75t_L g453 ( .A(n_193), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_193), .B(n_414), .Y(n_464) );
AND2x4_ASAP7_75t_L g193 ( .A(n_194), .B(n_205), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2x1_ASAP7_75t_L g243 ( .A(n_195), .B(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g390 ( .A(n_195), .B(n_329), .Y(n_390) );
AND2x2_ASAP7_75t_L g394 ( .A(n_195), .B(n_249), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_203), .Y(n_228) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_203), .A2(n_549), .B(n_553), .Y(n_548) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g238 ( .A(n_205), .Y(n_238) );
INVx2_ASAP7_75t_L g283 ( .A(n_205), .Y(n_283) );
AND2x2_ASAP7_75t_L g328 ( .A(n_205), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_207), .B(n_213), .Y(n_206) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_226), .Y(n_216) );
OR2x6_ASAP7_75t_L g396 ( .A(n_217), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g400 ( .A(n_217), .B(n_401), .Y(n_400) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx4_ASAP7_75t_L g259 ( .A(n_218), .Y(n_259) );
AND2x4_ASAP7_75t_L g267 ( .A(n_218), .B(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g302 ( .A(n_218), .B(n_227), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_218), .B(n_325), .Y(n_348) );
AND2x2_ASAP7_75t_L g364 ( .A(n_218), .B(n_255), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_218), .B(n_320), .Y(n_418) );
INVx2_ASAP7_75t_L g433 ( .A(n_218), .Y(n_433) );
OR2x6_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
AND2x2_ASAP7_75t_L g278 ( .A(n_226), .B(n_267), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_226), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_SL g382 ( .A(n_226), .B(n_305), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_226), .B(n_318), .Y(n_411) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_227), .Y(n_257) );
AND2x2_ASAP7_75t_L g265 ( .A(n_227), .B(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_227), .Y(n_288) );
INVx2_ASAP7_75t_L g291 ( .A(n_227), .Y(n_291) );
INVx1_ASAP7_75t_L g324 ( .A(n_227), .Y(n_324) );
INVx1_ASAP7_75t_L g402 ( .A(n_227), .Y(n_402) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_235), .Y(n_227) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_228), .A2(n_509), .B(n_515), .Y(n_508) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_228), .A2(n_518), .B(n_524), .Y(n_517) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_228), .A2(n_518), .B(n_524), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
NAND2xp33_ASAP7_75t_L g236 ( .A(n_237), .B(n_240), .Y(n_236) );
OR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_238), .B(n_241), .Y(n_314) );
AND4x1_ASAP7_75t_SL g404 ( .A(n_238), .B(n_379), .C(n_405), .D(n_407), .Y(n_404) );
OR2x2_ASAP7_75t_L g458 ( .A(n_238), .B(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g350 ( .A(n_239), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
AND2x2_ASAP7_75t_L g293 ( .A(n_242), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_242), .B(n_251), .Y(n_416) );
AND2x2_ASAP7_75t_L g362 ( .A(n_243), .B(n_328), .Y(n_362) );
OAI32xp33_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_253), .A3(n_258), .B1(n_260), .B2(n_263), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g413 ( .A(n_248), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g426 ( .A(n_248), .B(n_344), .Y(n_426) );
AND2x4_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
INVx1_ASAP7_75t_L g389 ( .A(n_249), .Y(n_389) );
AND2x2_ASAP7_75t_L g423 ( .A(n_249), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_250), .B(n_252), .Y(n_351) );
INVx3_ASAP7_75t_L g274 ( .A(n_251), .Y(n_274) );
NAND2x1p5_ASAP7_75t_L g339 ( .A(n_251), .B(n_340), .Y(n_339) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_252), .Y(n_311) );
AND2x2_ASAP7_75t_L g330 ( .A(n_252), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g358 ( .A(n_254), .Y(n_358) );
NAND2x1_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g304 ( .A(n_255), .Y(n_304) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_255), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_258), .B(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g296 ( .A(n_259), .B(n_264), .Y(n_296) );
AND2x4_ASAP7_75t_L g318 ( .A(n_259), .B(n_268), .Y(n_318) );
AND2x4_ASAP7_75t_SL g368 ( .A(n_259), .B(n_369), .Y(n_368) );
NOR2x1_ASAP7_75t_L g380 ( .A(n_259), .B(n_336), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_260), .A2(n_456), .B1(n_458), .B2(n_460), .Y(n_455) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx2_ASAP7_75t_SL g468 ( .A(n_261), .Y(n_468) );
INVx2_ASAP7_75t_L g294 ( .A(n_262), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_265), .B(n_271), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_265), .A2(n_467), .B1(n_470), .B2(n_473), .Y(n_469) );
INVx1_ASAP7_75t_L g325 ( .A(n_266), .Y(n_325) );
AND2x2_ASAP7_75t_L g398 ( .A(n_266), .B(n_307), .Y(n_398) );
INVx2_ASAP7_75t_L g271 ( .A(n_267), .Y(n_271) );
OAI21xp5_ASAP7_75t_SL g269 ( .A1(n_270), .A2(n_272), .B(n_276), .Y(n_269) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_273), .A2(n_428), .B1(n_431), .B2(n_432), .Y(n_427) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_274), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_274), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g443 ( .A(n_274), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
NOR3xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_295), .C(n_299), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_284), .B1(n_289), .B2(n_292), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g309 ( .A(n_282), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g370 ( .A(n_282), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g383 ( .A(n_282), .B(n_372), .Y(n_383) );
AND2x2_ASAP7_75t_L g431 ( .A(n_282), .B(n_390), .Y(n_431) );
AND2x2_ASAP7_75t_L g467 ( .A(n_282), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx4_ASAP7_75t_L g336 ( .A(n_285), .Y(n_336) );
AND2x2_ASAP7_75t_L g432 ( .A(n_285), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx2_ASAP7_75t_L g437 ( .A(n_288), .Y(n_437) );
AND2x2_ASAP7_75t_L g445 ( .A(n_288), .B(n_398), .Y(n_445) );
INVx1_ASAP7_75t_L g347 ( .A(n_290), .Y(n_347) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g320 ( .A(n_291), .Y(n_320) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_293), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_294), .B(n_443), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_303), .B(n_308), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_301), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
AOI21xp33_ASAP7_75t_SL g312 ( .A1(n_304), .A2(n_313), .B(n_315), .Y(n_312) );
AND2x2_ASAP7_75t_L g353 ( .A(n_304), .B(n_318), .Y(n_353) );
AND2x4_ASAP7_75t_L g322 ( .A(n_305), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_305), .B(n_402), .Y(n_410) );
INVx2_ASAP7_75t_SL g438 ( .A(n_305), .Y(n_438) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AOI21xp33_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_321), .B(n_326), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_318), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_318), .B(n_323), .Y(n_466) );
AND2x2_ASAP7_75t_L g363 ( .A(n_319), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g367 ( .A(n_319), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g406 ( .A(n_319), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_319), .B(n_336), .Y(n_425) );
INVx1_ASAP7_75t_L g454 ( .A(n_319), .Y(n_454) );
INVx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_SL g323 ( .A(n_324), .B(n_325), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_324), .B(n_398), .Y(n_430) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx1_ASAP7_75t_L g338 ( .A(n_328), .Y(n_338) );
AND2x2_ASAP7_75t_L g344 ( .A(n_329), .B(n_341), .Y(n_344) );
INVxp67_ASAP7_75t_L g480 ( .A(n_332), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_332), .B(n_375), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_359), .Y(n_332) );
NOR3xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_349), .C(n_356), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_337), .B1(n_342), .B2(n_345), .Y(n_334) );
INVx2_ASAP7_75t_L g373 ( .A(n_336), .Y(n_373) );
NAND2xp5_ASAP7_75t_R g391 ( .A(n_336), .B(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx3_ASAP7_75t_L g387 ( .A(n_340), .Y(n_387) );
BUFx3_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g439 ( .A(n_343), .Y(n_439) );
INVx2_ASAP7_75t_L g459 ( .A(n_344), .Y(n_459) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_346), .A2(n_463), .B1(n_465), .B2(n_467), .Y(n_462) );
NOR2x1_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
NOR3xp33_ASAP7_75t_L g356 ( .A(n_350), .B(n_355), .C(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI222xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_363), .B1(n_365), .B2(n_367), .C1(n_370), .C2(n_373), .Y(n_359) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_364), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_SL g392 ( .A(n_368), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_368), .B(n_437), .Y(n_460) );
INVx1_ASAP7_75t_L g414 ( .A(n_371), .Y(n_414) );
OA21x2_ASAP7_75t_L g449 ( .A1(n_371), .A2(n_450), .B(n_451), .Y(n_449) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g393 ( .A(n_372), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g407 ( .A(n_372), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_419), .Y(n_374) );
INVxp67_ASAP7_75t_L g481 ( .A(n_375), .Y(n_481) );
NAND3xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_384), .C(n_403), .Y(n_375) );
NOR2x1_ASAP7_75t_L g376 ( .A(n_377), .B(n_381), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_391), .B1(n_393), .B2(n_395), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx2_ASAP7_75t_L g452 ( .A(n_387), .Y(n_452) );
NAND2x1p5_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
AND2x2_ASAP7_75t_L g422 ( .A(n_390), .B(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_399), .Y(n_395) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_399), .A2(n_441), .B1(n_444), .B2(n_446), .Y(n_440) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g470 ( .A(n_402), .B(n_471), .Y(n_470) );
NOR3xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_408), .C(n_415), .Y(n_403) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g457 ( .A(n_406), .B(n_432), .Y(n_457) );
AOI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_411), .B(n_412), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVxp67_ASAP7_75t_L g476 ( .A(n_419), .Y(n_476) );
NAND4xp75_ASAP7_75t_L g419 ( .A(n_420), .B(n_434), .C(n_448), .D(n_461), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_427), .Y(n_420) );
NAND2x1p5_ASAP7_75t_L g474 ( .A(n_423), .B(n_468), .Y(n_474) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g472 ( .A(n_433), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_439), .B(n_440), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_438), .B(n_452), .Y(n_451) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_453), .B(n_455), .Y(n_448) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_469), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B(n_478), .Y(n_475) );
AOI21xp5_ASAP7_75t_SL g479 ( .A1(n_478), .A2(n_480), .B(n_481), .Y(n_479) );
INVx4_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
INVx3_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_485), .Y(n_484) );
AND2x6_ASAP7_75t_SL g485 ( .A(n_486), .B(n_487), .Y(n_485) );
OR2x6_ASAP7_75t_SL g774 ( .A(n_486), .B(n_775), .Y(n_774) );
OR2x2_ASAP7_75t_L g783 ( .A(n_486), .B(n_487), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_486), .B(n_775), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g775 ( .A(n_487), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
INVx3_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_702), .Y(n_492) );
NOR4xp25_ASAP7_75t_SL g493 ( .A(n_494), .B(n_595), .C(n_639), .D(n_666), .Y(n_493) );
OAI221xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_558), .B1(n_568), .B2(n_583), .C(n_585), .Y(n_494) );
AOI32xp33_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_525), .A3(n_532), .B1(n_543), .B2(n_554), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_496), .B(n_738), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_496), .A2(n_708), .B1(n_766), .B2(n_769), .Y(n_765) );
AND2x4_ASAP7_75t_SL g496 ( .A(n_497), .B(n_507), .Y(n_496) );
INVx5_ASAP7_75t_L g557 ( .A(n_497), .Y(n_557) );
OR2x2_ASAP7_75t_L g584 ( .A(n_497), .B(n_556), .Y(n_584) );
AND2x4_ASAP7_75t_L g586 ( .A(n_497), .B(n_517), .Y(n_586) );
INVx2_ASAP7_75t_L g601 ( .A(n_497), .Y(n_601) );
OR2x2_ASAP7_75t_L g613 ( .A(n_497), .B(n_526), .Y(n_613) );
AND2x2_ASAP7_75t_L g620 ( .A(n_497), .B(n_516), .Y(n_620) );
AND2x2_ASAP7_75t_SL g662 ( .A(n_497), .B(n_545), .Y(n_662) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_497), .Y(n_719) );
OR2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
INVx3_ASAP7_75t_SL g614 ( .A(n_507), .Y(n_614) );
AND2x2_ASAP7_75t_L g633 ( .A(n_507), .B(n_557), .Y(n_633) );
AOI32xp33_ASAP7_75t_L g748 ( .A1(n_507), .A2(n_619), .A3(n_649), .B1(n_679), .B2(n_714), .Y(n_748) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_516), .Y(n_507) );
AND2x2_ASAP7_75t_L g588 ( .A(n_508), .B(n_526), .Y(n_588) );
OR2x2_ASAP7_75t_L g604 ( .A(n_508), .B(n_517), .Y(n_604) );
INVx1_ASAP7_75t_L g627 ( .A(n_508), .Y(n_627) );
INVx2_ASAP7_75t_L g643 ( .A(n_508), .Y(n_643) );
AND2x2_ASAP7_75t_L g680 ( .A(n_508), .B(n_545), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_508), .B(n_517), .Y(n_699) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_508), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_514), .Y(n_509) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g735 ( .A(n_517), .B(n_526), .Y(n_735) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_517), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .Y(n_518) );
OR2x2_ASAP7_75t_L g583 ( .A(n_525), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g589 ( .A(n_525), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g602 ( .A(n_525), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g764 ( .A(n_525), .B(n_633), .Y(n_764) );
BUFx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g693 ( .A(n_526), .B(n_643), .Y(n_693) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_527), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_532), .B(n_660), .Y(n_762) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_533), .B(n_710), .Y(n_709) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g547 ( .A(n_534), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g569 ( .A(n_534), .Y(n_569) );
AND2x2_ASAP7_75t_L g593 ( .A(n_534), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_534), .B(n_571), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_534), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g651 ( .A(n_534), .Y(n_651) );
OR2x2_ASAP7_75t_L g670 ( .A(n_534), .B(n_597), .Y(n_670) );
INVx1_ASAP7_75t_L g677 ( .A(n_534), .Y(n_677) );
NOR2xp33_ASAP7_75t_R g729 ( .A(n_534), .B(n_560), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_534), .B(n_572), .Y(n_733) );
INVx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_541), .Y(n_536) );
AOI32xp33_ASAP7_75t_L g756 ( .A1(n_543), .A2(n_592), .A3(n_757), .B1(n_758), .B2(n_759), .Y(n_756) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
INVx2_ASAP7_75t_L g623 ( .A(n_545), .Y(n_623) );
AND2x4_ASAP7_75t_L g642 ( .A(n_545), .B(n_643), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_545), .B(n_614), .Y(n_671) );
OR2x2_ASAP7_75t_L g725 ( .A(n_545), .B(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g683 ( .A(n_546), .B(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g741 ( .A(n_546), .B(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_547), .B(n_560), .Y(n_707) );
AND2x2_ASAP7_75t_L g744 ( .A(n_547), .B(n_710), .Y(n_744) );
INVx2_ASAP7_75t_L g594 ( .A(n_548), .Y(n_594) );
INVx2_ASAP7_75t_L g597 ( .A(n_548), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_548), .B(n_560), .Y(n_617) );
INVx1_ASAP7_75t_L g648 ( .A(n_548), .Y(n_648) );
OR2x2_ASAP7_75t_L g674 ( .A(n_548), .B(n_560), .Y(n_674) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_548), .Y(n_726) );
BUFx3_ASAP7_75t_L g755 ( .A(n_548), .Y(n_755) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g624 ( .A(n_555), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_555), .B(n_642), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_555), .B(n_713), .Y(n_712) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_556), .B(n_627), .Y(n_626) );
OAI21xp33_ASAP7_75t_L g656 ( .A1(n_556), .A2(n_623), .B(n_641), .Y(n_656) );
OAI32xp33_ASAP7_75t_L g678 ( .A1(n_557), .A2(n_679), .A3(n_681), .B1(n_683), .B2(n_685), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_557), .B(n_642), .Y(n_751) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g684 ( .A(n_559), .Y(n_684) );
NOR2x1p5_ASAP7_75t_L g754 ( .A(n_559), .B(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x4_ASAP7_75t_L g570 ( .A(n_560), .B(n_571), .Y(n_570) );
AND2x4_ASAP7_75t_SL g592 ( .A(n_560), .B(n_572), .Y(n_592) );
OR2x2_ASAP7_75t_L g596 ( .A(n_560), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g631 ( .A(n_560), .Y(n_631) );
AND2x2_ASAP7_75t_L g649 ( .A(n_560), .B(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g660 ( .A(n_560), .B(n_572), .Y(n_660) );
OR2x2_ASAP7_75t_L g722 ( .A(n_560), .B(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g739 ( .A(n_560), .B(n_670), .Y(n_739) );
INVx1_ASAP7_75t_L g771 ( .A(n_560), .Y(n_771) );
OR2x6_ASAP7_75t_L g560 ( .A(n_561), .B(n_567), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_569), .B(n_648), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_570), .B(n_682), .Y(n_681) );
AOI222xp33_ASAP7_75t_L g686 ( .A1(n_570), .A2(n_687), .B1(n_692), .B2(n_694), .C1(n_697), .C2(n_700), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_570), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g714 ( .A(n_570), .B(n_593), .Y(n_714) );
AND2x2_ASAP7_75t_L g676 ( .A(n_571), .B(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g691 ( .A(n_571), .B(n_596), .Y(n_691) );
INVx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_572), .B(n_597), .Y(n_629) );
AND2x4_ASAP7_75t_L g650 ( .A(n_572), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g710 ( .A(n_572), .B(n_631), .Y(n_710) );
AND2x4_ASAP7_75t_L g572 ( .A(n_573), .B(n_578), .Y(n_572) );
INVx1_ASAP7_75t_SL g590 ( .A(n_584), .Y(n_590) );
NAND2xp33_ASAP7_75t_SL g759 ( .A(n_584), .B(n_614), .Y(n_759) );
A2O1A1Ixp33_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B(n_589), .C(n_591), .Y(n_585) );
INVx2_ASAP7_75t_SL g636 ( .A(n_586), .Y(n_636) );
AND2x2_ASAP7_75t_L g640 ( .A(n_587), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_588), .B(n_636), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g661 ( .A1(n_588), .A2(n_626), .B(n_662), .C(n_663), .Y(n_661) );
AND2x2_ASAP7_75t_L g738 ( .A(n_588), .B(n_719), .Y(n_738) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
AND2x4_ASAP7_75t_L g637 ( .A(n_592), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_SL g742 ( .A(n_592), .Y(n_742) );
OAI211xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_598), .B(n_605), .C(n_632), .Y(n_595) );
INVx2_ASAP7_75t_L g607 ( .A(n_596), .Y(n_607) );
OR2x2_ASAP7_75t_L g654 ( .A(n_596), .B(n_655), .Y(n_654) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_597), .Y(n_638) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_600), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g692 ( .A(n_600), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_600), .B(n_680), .Y(n_746) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AOI222xp33_ASAP7_75t_L g704 ( .A1(n_602), .A2(n_705), .B1(n_706), .B2(n_708), .C1(n_711), .C2(n_714), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_603), .A2(n_668), .B1(n_671), .B2(n_672), .C(n_678), .Y(n_667) );
AND2x2_ASAP7_75t_L g705 ( .A(n_603), .B(n_662), .Y(n_705) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp33_ASAP7_75t_SL g618 ( .A(n_604), .B(n_619), .Y(n_618) );
AOI221x1_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_610), .B1(n_615), .B2(n_618), .C(n_621), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
AND2x2_ASAP7_75t_L g758 ( .A(n_608), .B(n_696), .Y(n_758) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g616 ( .A(n_609), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
OAI32xp33_ASAP7_75t_L g724 ( .A1(n_614), .A2(n_655), .A3(n_725), .B1(n_727), .B2(n_731), .Y(n_724) );
OAI21xp33_ASAP7_75t_SL g743 ( .A1(n_615), .A2(n_744), .B(n_745), .Y(n_743) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AOI21xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_625), .B(n_628), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
OR2x2_ASAP7_75t_L g625 ( .A(n_623), .B(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g698 ( .A(n_623), .B(n_699), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_627), .A2(n_653), .B1(n_656), .B2(n_657), .C(n_661), .Y(n_652) );
INVx1_ASAP7_75t_L g728 ( .A(n_627), .Y(n_728) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_627), .Y(n_734) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
OAI21xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B(n_637), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_636), .B(n_701), .Y(n_700) );
OAI21xp5_ASAP7_75t_SL g639 ( .A1(n_640), .A2(n_644), .B(n_652), .Y(n_639) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_643), .Y(n_713) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_649), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_646), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVxp67_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g665 ( .A(n_648), .Y(n_665) );
INVx1_ASAP7_75t_L g655 ( .A(n_650), .Y(n_655) );
AND2x2_ASAP7_75t_SL g664 ( .A(n_650), .B(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_650), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_650), .B(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g669 ( .A(n_660), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_665), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_667), .B(n_686), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g682 ( .A(n_670), .Y(n_682) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx1_ASAP7_75t_SL g696 ( .A(n_674), .Y(n_696) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_676), .B(n_754), .Y(n_753) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_677), .Y(n_690) );
BUFx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_688), .B(n_691), .Y(n_687) );
INVxp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g701 ( .A(n_693), .Y(n_701) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g720 ( .A(n_699), .Y(n_720) );
NOR4xp25_ASAP7_75t_L g702 ( .A(n_703), .B(n_736), .C(n_747), .D(n_760), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_715), .Y(n_703) );
O2A1O1Ixp33_ASAP7_75t_L g715 ( .A1(n_705), .A2(n_716), .B(n_721), .C(n_724), .Y(n_715) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_SL g717 ( .A(n_718), .B(n_720), .Y(n_717) );
OAI211xp5_ASAP7_75t_L g727 ( .A1(n_718), .A2(n_728), .B(n_729), .C(n_730), .Y(n_727) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
OAI21xp33_ASAP7_75t_SL g731 ( .A1(n_732), .A2(n_734), .B(n_735), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_SL g766 ( .A(n_735), .B(n_767), .Y(n_766) );
OAI221xp5_ASAP7_75t_SL g736 ( .A1(n_737), .A2(n_739), .B1(n_740), .B2(n_741), .C(n_743), .Y(n_736) );
INVx1_ASAP7_75t_SL g740 ( .A(n_738), .Y(n_740) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND3xp33_ASAP7_75t_SL g747 ( .A(n_748), .B(n_749), .C(n_756), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_752), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
OAI21xp33_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_763), .B(n_765), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVxp33_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_773), .Y(n_772) );
CKINVDCx11_ASAP7_75t_R g773 ( .A(n_774), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g777 ( .A1(n_776), .A2(n_778), .B(n_779), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
INVx1_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_793), .Y(n_786) );
INVxp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g788 ( .A(n_789), .B(n_792), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
OR2x2_ASAP7_75t_SL g817 ( .A(n_790), .B(n_792), .Y(n_817) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_790), .A2(n_820), .B(n_823), .Y(n_819) );
BUFx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
OR2x2_ASAP7_75t_L g806 ( .A(n_794), .B(n_807), .Y(n_806) );
BUFx2_ASAP7_75t_R g813 ( .A(n_794), .Y(n_813) );
BUFx2_ASAP7_75t_L g824 ( .A(n_794), .Y(n_824) );
INVxp67_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
OAI21x1_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_808), .B(n_811), .Y(n_796) );
OAI21xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_801), .B(n_806), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
NOR2x1_ASAP7_75t_L g808 ( .A(n_799), .B(n_809), .Y(n_808) );
INVxp67_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
BUFx2_ASAP7_75t_L g810 ( .A(n_803), .Y(n_810) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_806), .B(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_SL g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_SL g814 ( .A(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_SL g818 ( .A(n_819), .Y(n_818) );
CKINVDCx11_ASAP7_75t_R g820 ( .A(n_821), .Y(n_820) );
CKINVDCx8_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
endmodule