module fake_jpeg_25700_n_310 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_22),
.B(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_40),
.Y(n_48)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_44),
.B(n_32),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_52),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_17),
.B1(n_25),
.B2(n_18),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_51),
.B1(n_31),
.B2(n_39),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_50),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_17),
.B1(n_25),
.B2(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_37),
.B1(n_39),
.B2(n_17),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_61),
.A2(n_87),
.B1(n_40),
.B2(n_38),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_58),
.A2(n_18),
.B1(n_31),
.B2(n_30),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_65),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_64),
.B(n_74),
.Y(n_123)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_76),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_43),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_69),
.A2(n_78),
.B(n_65),
.Y(n_95)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_19),
.B1(n_16),
.B2(n_40),
.Y(n_103)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_93),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_58),
.A2(n_30),
.B1(n_28),
.B2(n_21),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_84),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_39),
.B1(n_20),
.B2(n_23),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_48),
.B1(n_41),
.B2(n_19),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_43),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_41),
.B1(n_42),
.B2(n_40),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_48),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_91),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_57),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_21),
.Y(n_92)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_95),
.B(n_61),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_117),
.B1(n_118),
.B2(n_78),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_34),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_81),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_75),
.A2(n_16),
.B1(n_33),
.B2(n_23),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_99),
.A2(n_110),
.B1(n_122),
.B2(n_73),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_103),
.A2(n_112),
.B1(n_87),
.B2(n_86),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_20),
.B1(n_23),
.B2(n_26),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_67),
.A2(n_40),
.B1(n_38),
.B2(n_36),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_82),
.A2(n_40),
.B1(n_38),
.B2(n_36),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_78),
.A2(n_23),
.B1(n_20),
.B2(n_40),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_71),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_126),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_146),
.B1(n_116),
.B2(n_89),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_101),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_130),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_149),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_69),
.B1(n_63),
.B2(n_66),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_147),
.B1(n_112),
.B2(n_96),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_135),
.Y(n_163)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_69),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_97),
.B1(n_116),
.B2(n_79),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_91),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_140),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_101),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_139),
.A2(n_142),
.B(n_145),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_64),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_108),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_141),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_95),
.B(n_36),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_76),
.Y(n_143)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_34),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_118),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_111),
.A2(n_0),
.B(n_1),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_59),
.B1(n_70),
.B2(n_74),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_83),
.Y(n_148)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_120),
.C(n_100),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_104),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_150),
.A2(n_26),
.B(n_24),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_88),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_151),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_153),
.B1(n_160),
.B2(n_170),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_144),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_140),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_157),
.B(n_165),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_158),
.A2(n_172),
.B1(n_177),
.B2(n_180),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_129),
.A2(n_114),
.B1(n_107),
.B2(n_105),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_141),
.A2(n_121),
.B1(n_114),
.B2(n_102),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_105),
.B(n_107),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_169),
.A2(n_182),
.B(n_0),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_139),
.A2(n_109),
.B1(n_115),
.B2(n_104),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_109),
.B1(n_115),
.B2(n_102),
.Y(n_172)
);

AO22x1_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_102),
.B1(n_68),
.B2(n_60),
.Y(n_173)
);

AO22x2_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_128),
.B1(n_130),
.B2(n_150),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_26),
.B1(n_24),
.B2(n_34),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_178),
.B1(n_152),
.B2(n_181),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_26),
.B1(n_24),
.B2(n_8),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_135),
.A2(n_26),
.B1(n_24),
.B2(n_8),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_127),
.Y(n_193)
);

XNOR2x1_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_149),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_188),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_162),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_205),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_143),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_191),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_174),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_189),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_126),
.Y(n_190)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_131),
.Y(n_191)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_196),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_193),
.A2(n_195),
.B(n_197),
.Y(n_224)
);

XOR2x1_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_138),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_168),
.B(n_159),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_198),
.A2(n_210),
.B(n_1),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_133),
.C(n_137),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_200),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_148),
.C(n_124),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_206),
.B1(n_177),
.B2(n_180),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_134),
.C(n_7),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_203),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_6),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_15),
.Y(n_204)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_164),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_160),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_5),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_209),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_167),
.B(n_14),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_154),
.B(n_5),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_211),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_170),
.B1(n_179),
.B2(n_166),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_213),
.A2(n_214),
.B1(n_221),
.B2(n_227),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_208),
.A2(n_166),
.B1(n_158),
.B2(n_167),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_184),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_208),
.A2(n_172),
.B1(n_171),
.B2(n_178),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_198),
.Y(n_226)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_185),
.A2(n_173),
.B1(n_155),
.B2(n_161),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_173),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_182),
.B1(n_7),
.B2(n_9),
.Y(n_231)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_198),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_192),
.Y(n_234)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_218),
.B(n_200),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_246),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_239),
.A2(n_230),
.B(n_226),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_199),
.C(n_188),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_244),
.C(n_248),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_191),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_251),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_183),
.C(n_195),
.Y(n_244)
);

NOR2x1_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_197),
.Y(n_245)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_197),
.C(n_203),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_207),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_252),
.B1(n_222),
.B2(n_228),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_197),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_216),
.C(n_224),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_259),
.C(n_260),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_224),
.C(n_221),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_213),
.C(n_214),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_262),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_239),
.B1(n_238),
.B2(n_245),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_266),
.B1(n_243),
.B2(n_3),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_226),
.B1(n_233),
.B2(n_229),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_240),
.A2(n_222),
.B(n_9),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_12),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_9),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_236),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_279),
.Y(n_289)
);

NAND2xp33_ASAP7_75t_SL g287 ( 
.A(n_270),
.B(n_280),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_237),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_272),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_278),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_276),
.B(n_266),
.Y(n_283)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_261),
.A2(n_11),
.B1(n_12),
.B2(n_4),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_263),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_254),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_282),
.C(n_268),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_253),
.C(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_286),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_259),
.C(n_253),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_292),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_274),
.B(n_277),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_291),
.A2(n_287),
.B(n_269),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_260),
.C(n_276),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_295),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_254),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_265),
.B(n_262),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_295),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_302),
.C(n_297),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_264),
.B(n_3),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_304),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g306 ( 
.A(n_305),
.B(n_298),
.CI(n_300),
.CON(n_306),
.SN(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_296),
.C(n_2),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_306),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_2),
.C(n_4),
.Y(n_309)
);

AO21x1_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_2),
.B(n_4),
.Y(n_310)
);


endmodule