module real_aes_2298_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_500;
wire n_307;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AO22x2_ASAP7_75t_L g115 ( .A1(n_0), .A2(n_56), .B1(n_112), .B2(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_1), .B(n_229), .Y(n_305) );
AOI22xp33_ASAP7_75t_SL g524 ( .A1(n_1), .A2(n_101), .B1(n_102), .B2(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_1), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_2), .B(n_255), .Y(n_267) );
XOR2xp5_ASAP7_75t_L g532 ( .A(n_3), .B(n_102), .Y(n_532) );
INVx1_ASAP7_75t_L g90 ( .A(n_4), .Y(n_90) );
AO22x2_ASAP7_75t_L g111 ( .A1(n_5), .A2(n_17), .B1(n_112), .B2(n_113), .Y(n_111) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_6), .A2(n_21), .B1(n_184), .B2(n_187), .Y(n_183) );
AND2x2_ASAP7_75t_L g258 ( .A(n_7), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g269 ( .A(n_8), .B(n_270), .Y(n_269) );
AOI22xp33_ASAP7_75t_SL g143 ( .A1(n_9), .A2(n_38), .B1(n_144), .B2(n_146), .Y(n_143) );
INVx2_ASAP7_75t_L g218 ( .A(n_10), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_11), .B(n_255), .Y(n_324) );
INVx1_ASAP7_75t_L g98 ( .A(n_12), .Y(n_98) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_12), .B(n_229), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_13), .A2(n_32), .B1(n_149), .B2(n_153), .Y(n_148) );
OAI22xp5_ASAP7_75t_SL g96 ( .A1(n_14), .A2(n_97), .B1(n_98), .B2(n_99), .Y(n_96) );
INVx1_ASAP7_75t_L g99 ( .A(n_14), .Y(n_99) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_14), .A2(n_71), .B1(n_222), .B2(n_229), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_15), .A2(n_68), .B1(n_198), .B2(n_199), .Y(n_197) );
INVx1_ASAP7_75t_L g199 ( .A(n_15), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_16), .A2(n_19), .B1(n_175), .B2(n_178), .Y(n_174) );
OAI221xp5_ASAP7_75t_L g82 ( .A1(n_17), .A2(n_56), .B1(n_60), .B2(n_83), .C(n_85), .Y(n_82) );
OR2x2_ASAP7_75t_L g219 ( .A(n_18), .B(n_70), .Y(n_219) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_18), .A2(n_70), .B(n_218), .Y(n_248) );
INVx3_ASAP7_75t_L g112 ( .A(n_20), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_22), .A2(n_192), .B1(n_202), .B2(n_203), .Y(n_191) );
INVx1_ASAP7_75t_L g202 ( .A(n_22), .Y(n_202) );
AO21x2_ASAP7_75t_L g319 ( .A1(n_23), .A2(n_259), .B(n_320), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_24), .A2(n_237), .B(n_265), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_25), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_26), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_27), .B(n_255), .Y(n_304) );
INVx1_ASAP7_75t_SL g121 ( .A(n_28), .Y(n_121) );
INVx1_ASAP7_75t_L g92 ( .A(n_29), .Y(n_92) );
AND2x2_ASAP7_75t_L g227 ( .A(n_29), .B(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g235 ( .A(n_29), .B(n_90), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_30), .B(n_229), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_31), .B(n_255), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_33), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_34), .B(n_229), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_35), .A2(n_237), .B(n_251), .Y(n_250) );
AO22x2_ASAP7_75t_L g124 ( .A1(n_36), .A2(n_60), .B1(n_112), .B2(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_37), .B(n_253), .Y(n_281) );
AOI22xp33_ASAP7_75t_SL g131 ( .A1(n_39), .A2(n_66), .B1(n_132), .B2(n_137), .Y(n_131) );
AOI22xp33_ASAP7_75t_SL g105 ( .A1(n_40), .A2(n_50), .B1(n_106), .B2(n_126), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_41), .B(n_229), .Y(n_321) );
INVx1_ASAP7_75t_L g225 ( .A(n_42), .Y(n_225) );
INVx1_ASAP7_75t_L g232 ( .A(n_42), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_43), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g289 ( .A(n_44), .B(n_216), .Y(n_289) );
INVx1_ASAP7_75t_L g122 ( .A(n_45), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_46), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_47), .B(n_253), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_48), .B(n_229), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_49), .B(n_229), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_51), .A2(n_237), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g541 ( .A(n_51), .Y(n_541) );
AND2x2_ASAP7_75t_L g315 ( .A(n_52), .B(n_217), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_53), .B(n_253), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_54), .B(n_253), .Y(n_325) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_55), .A2(n_72), .B1(n_237), .B2(n_239), .Y(n_236) );
INVxp33_ASAP7_75t_L g87 ( .A(n_56), .Y(n_87) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_57), .B(n_255), .Y(n_312) );
INVx1_ASAP7_75t_L g228 ( .A(n_58), .Y(n_228) );
INVx1_ASAP7_75t_L g234 ( .A(n_58), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_59), .B(n_253), .Y(n_266) );
INVxp67_ASAP7_75t_L g86 ( .A(n_60), .Y(n_86) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_61), .A2(n_237), .B(n_293), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_62), .A2(n_237), .B(n_279), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_63), .A2(n_237), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g306 ( .A(n_64), .B(n_217), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_65), .B(n_216), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_67), .A2(n_196), .B1(n_197), .B2(n_200), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_67), .Y(n_196) );
INVx1_ASAP7_75t_L g198 ( .A(n_68), .Y(n_198) );
AND2x2_ASAP7_75t_L g282 ( .A(n_69), .B(n_270), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_73), .A2(n_237), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_74), .B(n_255), .Y(n_280) );
INVxp67_ASAP7_75t_L g194 ( .A(n_75), .Y(n_194) );
BUFx2_ASAP7_75t_L g314 ( .A(n_76), .Y(n_314) );
BUFx2_ASAP7_75t_SL g84 ( .A(n_77), .Y(n_84) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_93), .B1(n_204), .B2(n_521), .C(n_523), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
AND3x1_ASAP7_75t_SL g81 ( .A(n_82), .B(n_88), .C(n_91), .Y(n_81) );
INVxp67_ASAP7_75t_L g531 ( .A(n_82), .Y(n_531) );
CKINVDCx8_ASAP7_75t_R g83 ( .A(n_84), .Y(n_83) );
NOR2xp33_ASAP7_75t_L g85 ( .A(n_86), .B(n_87), .Y(n_85) );
CKINVDCx16_ASAP7_75t_R g529 ( .A(n_88), .Y(n_529) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_88), .A2(n_538), .B(n_540), .Y(n_537) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x2_ASAP7_75t_L g223 ( .A(n_89), .B(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_SL g535 ( .A(n_89), .B(n_91), .Y(n_535) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
AND2x2_ASAP7_75t_L g238 ( .A(n_90), .B(n_225), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_91), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
NOR2x1p5_ASAP7_75t_L g240 ( .A(n_92), .B(n_241), .Y(n_240) );
XOR2xp5_ASAP7_75t_L g93 ( .A(n_94), .B(n_191), .Y(n_93) );
AOI22xp5_ASAP7_75t_L g94 ( .A1(n_95), .A2(n_96), .B1(n_100), .B2(n_101), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_96), .Y(n_95) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x4_ASAP7_75t_L g102 ( .A(n_103), .B(n_156), .Y(n_102) );
NOR2x1_ASAP7_75t_L g103 ( .A(n_104), .B(n_142), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_105), .B(n_131), .Y(n_104) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx8_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_117), .Y(n_108) );
AND2x2_ASAP7_75t_L g145 ( .A(n_109), .B(n_136), .Y(n_145) );
AND2x4_ASAP7_75t_L g151 ( .A(n_109), .B(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g165 ( .A(n_109), .B(n_166), .Y(n_165) );
AND2x4_ASAP7_75t_L g109 ( .A(n_110), .B(n_114), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g130 ( .A(n_111), .Y(n_130) );
AND2x2_ASAP7_75t_L g141 ( .A(n_111), .B(n_115), .Y(n_141) );
AND2x4_ASAP7_75t_L g147 ( .A(n_111), .B(n_114), .Y(n_147) );
INVx2_ASAP7_75t_L g113 ( .A(n_112), .Y(n_113) );
INVx1_ASAP7_75t_L g116 ( .A(n_112), .Y(n_116) );
OAI22x1_ASAP7_75t_L g119 ( .A1(n_112), .A2(n_120), .B1(n_121), .B2(n_122), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_112), .Y(n_120) );
INVx1_ASAP7_75t_L g125 ( .A(n_112), .Y(n_125) );
INVxp67_ASAP7_75t_L g190 ( .A(n_114), .Y(n_190) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g129 ( .A(n_115), .B(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g128 ( .A(n_117), .B(n_129), .Y(n_128) );
AND2x4_ASAP7_75t_L g146 ( .A(n_117), .B(n_147), .Y(n_146) );
AND2x4_ASAP7_75t_L g155 ( .A(n_117), .B(n_141), .Y(n_155) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_123), .Y(n_117) );
AND2x2_ASAP7_75t_L g136 ( .A(n_118), .B(n_124), .Y(n_136) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g152 ( .A(n_119), .B(n_123), .Y(n_152) );
AND2x2_ASAP7_75t_L g166 ( .A(n_119), .B(n_124), .Y(n_166) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_119), .Y(n_172) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx2_ASAP7_75t_L g140 ( .A(n_124), .Y(n_140) );
INVx2_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
INVx8_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g135 ( .A(n_129), .B(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g177 ( .A(n_129), .B(n_152), .Y(n_177) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_130), .Y(n_182) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x4_ASAP7_75t_L g186 ( .A(n_136), .B(n_147), .Y(n_186) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx5_ASAP7_75t_SL g138 ( .A(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_L g171 ( .A(n_141), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_148), .Y(n_142) );
BUFx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g161 ( .A(n_147), .B(n_152), .Y(n_161) );
INVx1_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
INVx6_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NOR2x1_ASAP7_75t_L g156 ( .A(n_157), .B(n_173), .Y(n_156) );
OAI222xp33_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_162), .B1(n_163), .B2(n_167), .C1(n_168), .C2(n_169), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx6f_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx6_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x4_ASAP7_75t_L g180 ( .A(n_166), .B(n_181), .Y(n_180) );
AND2x4_ASAP7_75t_L g189 ( .A(n_166), .B(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx12f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_183), .Y(n_173) );
BUFx6f_ASAP7_75t_SL g175 ( .A(n_176), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
BUFx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx6_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
CKINVDCx16_ASAP7_75t_R g203 ( .A(n_192), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B1(n_195), .B2(n_201), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_195), .Y(n_201) );
INVx1_ASAP7_75t_L g200 ( .A(n_197), .Y(n_200) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_458), .Y(n_205) );
NAND3xp33_ASAP7_75t_L g206 ( .A(n_207), .B(n_374), .C(n_411), .Y(n_206) );
NOR3xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_342), .C(n_357), .Y(n_207) );
OAI221xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_286), .B1(n_316), .B2(n_328), .C(n_329), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_211), .B(n_271), .Y(n_210) );
OAI22xp33_ASAP7_75t_SL g402 ( .A1(n_211), .A2(n_366), .B1(n_403), .B2(n_406), .Y(n_402) );
OR2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_243), .Y(n_211) );
OAI21xp33_ASAP7_75t_SL g412 ( .A1(n_212), .A2(n_413), .B(n_419), .Y(n_412) );
OR2x2_ASAP7_75t_L g441 ( .A(n_212), .B(n_273), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_212), .B(n_361), .Y(n_442) );
INVx2_ASAP7_75t_L g473 ( .A(n_212), .Y(n_473) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_213), .B(n_333), .Y(n_454) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g328 ( .A(n_214), .B(n_246), .Y(n_328) );
BUFx3_ASAP7_75t_L g354 ( .A(n_214), .Y(n_354) );
AND2x2_ASAP7_75t_L g490 ( .A(n_214), .B(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g513 ( .A(n_214), .B(n_274), .Y(n_513) );
AND2x4_ASAP7_75t_L g214 ( .A(n_215), .B(n_220), .Y(n_214) );
AND2x4_ASAP7_75t_L g285 ( .A(n_215), .B(n_220), .Y(n_285) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_216), .A2(n_221), .B(n_236), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_216), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_216), .A2(n_277), .B(n_278), .Y(n_276) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_SL g217 ( .A(n_218), .B(n_219), .Y(n_217) );
AND2x4_ASAP7_75t_L g296 ( .A(n_218), .B(n_219), .Y(n_296) );
AND2x4_ASAP7_75t_L g222 ( .A(n_223), .B(n_226), .Y(n_222) );
INVx1_ASAP7_75t_L g540 ( .A(n_223), .Y(n_540) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x4_ASAP7_75t_L g255 ( .A(n_225), .B(n_233), .Y(n_255) );
INVx1_ASAP7_75t_L g539 ( .A(n_226), .Y(n_539) );
BUFx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x6_ASAP7_75t_L g237 ( .A(n_227), .B(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g242 ( .A(n_228), .Y(n_242) );
AND2x6_ASAP7_75t_L g253 ( .A(n_228), .B(n_231), .Y(n_253) );
AND2x4_ASAP7_75t_L g229 ( .A(n_230), .B(n_235), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx5_ASAP7_75t_L g256 ( .A(n_235), .Y(n_256) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_237), .Y(n_522) );
AND2x4_ASAP7_75t_L g239 ( .A(n_238), .B(n_240), .Y(n_239) );
INVx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_244), .B(n_274), .Y(n_433) );
INVx1_ASAP7_75t_L g470 ( .A(n_244), .Y(n_470) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_260), .Y(n_244) );
AND2x2_ASAP7_75t_L g284 ( .A(n_245), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g491 ( .A(n_245), .Y(n_491) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g334 ( .A(n_246), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_246), .B(n_260), .Y(n_335) );
AND2x2_ASAP7_75t_L g356 ( .A(n_246), .B(n_275), .Y(n_356) );
AND2x2_ASAP7_75t_L g438 ( .A(n_246), .B(n_261), .Y(n_438) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_249), .B(n_258), .Y(n_246) );
INVx4_ASAP7_75t_L g259 ( .A(n_247), .Y(n_259) );
INVx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
BUFx4f_ASAP7_75t_L g270 ( .A(n_248), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_257), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_254), .B(n_256), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_253), .B(n_314), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_256), .A2(n_266), .B(n_267), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_256), .A2(n_280), .B(n_281), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_256), .A2(n_294), .B(n_295), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_256), .A2(n_303), .B(n_304), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_256), .A2(n_312), .B(n_313), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_256), .A2(n_324), .B(n_325), .Y(n_323) );
INVx3_ASAP7_75t_L g299 ( .A(n_259), .Y(n_299) );
AND2x4_ASAP7_75t_SL g331 ( .A(n_260), .B(n_275), .Y(n_331) );
INVx1_ASAP7_75t_L g362 ( .A(n_260), .Y(n_362) );
INVx2_ASAP7_75t_L g370 ( .A(n_260), .Y(n_370) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_260), .Y(n_394) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_261), .Y(n_283) );
AOI21x1_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_263), .B(n_269), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_268), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_270), .A2(n_309), .B(n_310), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_284), .Y(n_271) );
AND2x2_ASAP7_75t_L g509 ( .A(n_272), .B(n_372), .Y(n_509) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_283), .Y(n_273) );
NAND2x1p5_ASAP7_75t_L g368 ( .A(n_274), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g420 ( .A(n_274), .B(n_335), .Y(n_420) );
AND2x2_ASAP7_75t_L g437 ( .A(n_274), .B(n_438), .Y(n_437) );
INVx4_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g361 ( .A(n_275), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g377 ( .A(n_275), .Y(n_377) );
AND2x2_ASAP7_75t_L g421 ( .A(n_275), .B(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g428 ( .A(n_275), .B(n_429), .Y(n_428) );
NOR2x1_ASAP7_75t_L g443 ( .A(n_275), .B(n_334), .Y(n_443) );
BUFx2_ASAP7_75t_L g453 ( .A(n_275), .Y(n_453) );
AND2x2_ASAP7_75t_L g478 ( .A(n_275), .B(n_438), .Y(n_478) );
AND2x2_ASAP7_75t_L g499 ( .A(n_275), .B(n_500), .Y(n_499) );
OR2x6_ASAP7_75t_L g275 ( .A(n_276), .B(n_282), .Y(n_275) );
INVx1_ASAP7_75t_L g430 ( .A(n_283), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_284), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g460 ( .A(n_284), .B(n_331), .Y(n_460) );
INVx3_ASAP7_75t_L g367 ( .A(n_285), .Y(n_367) );
AND2x2_ASAP7_75t_L g500 ( .A(n_285), .B(n_422), .Y(n_500) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_287), .A2(n_330), .B1(n_335), .B2(n_336), .Y(n_329) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_297), .Y(n_287) );
INVx4_ASAP7_75t_L g327 ( .A(n_288), .Y(n_327) );
INVx2_ASAP7_75t_L g364 ( .A(n_288), .Y(n_364) );
NAND2x1_ASAP7_75t_L g390 ( .A(n_288), .B(n_307), .Y(n_390) );
OR2x2_ASAP7_75t_L g405 ( .A(n_288), .B(n_340), .Y(n_405) );
OR2x2_ASAP7_75t_SL g432 ( .A(n_288), .B(n_404), .Y(n_432) );
AND2x2_ASAP7_75t_L g445 ( .A(n_288), .B(n_319), .Y(n_445) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_288), .Y(n_466) );
OR2x6_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_292), .B(n_296), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_296), .A2(n_321), .B(n_322), .Y(n_320) );
INVx2_ASAP7_75t_L g345 ( .A(n_297), .Y(n_345) );
AND2x2_ASAP7_75t_L g477 ( .A(n_297), .B(n_451), .Y(n_477) );
NOR2x1_ASAP7_75t_SL g297 ( .A(n_298), .B(n_307), .Y(n_297) );
AND2x2_ASAP7_75t_L g318 ( .A(n_298), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g494 ( .A(n_298), .B(n_417), .Y(n_494) );
AO21x1_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_300), .B(n_306), .Y(n_298) );
AO21x2_ASAP7_75t_L g341 ( .A1(n_299), .A2(n_300), .B(n_306), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_305), .Y(n_300) );
OR2x2_ASAP7_75t_L g326 ( .A(n_307), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g337 ( .A(n_307), .B(n_327), .Y(n_337) );
AND2x2_ASAP7_75t_L g383 ( .A(n_307), .B(n_340), .Y(n_383) );
OR2x2_ASAP7_75t_L g404 ( .A(n_307), .B(n_319), .Y(n_404) );
INVx2_ASAP7_75t_SL g410 ( .A(n_307), .Y(n_410) );
AND2x2_ASAP7_75t_L g416 ( .A(n_307), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g426 ( .A(n_307), .B(n_409), .Y(n_426) );
BUFx2_ASAP7_75t_L g448 ( .A(n_307), .Y(n_448) );
OR2x6_ASAP7_75t_L g307 ( .A(n_308), .B(n_315), .Y(n_307) );
INVx2_ASAP7_75t_L g495 ( .A(n_316), .Y(n_495) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_326), .Y(n_316) );
OR2x2_ASAP7_75t_L g520 ( .A(n_317), .B(n_364), .Y(n_520) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_318), .B(n_327), .Y(n_386) );
AND2x2_ASAP7_75t_L g457 ( .A(n_318), .B(n_337), .Y(n_457) );
INVx1_ASAP7_75t_L g339 ( .A(n_319), .Y(n_339) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_319), .Y(n_348) );
INVx1_ASAP7_75t_L g381 ( .A(n_319), .Y(n_381) );
INVx2_ASAP7_75t_L g417 ( .A(n_319), .Y(n_417) );
NOR2xp67_ASAP7_75t_L g347 ( .A(n_327), .B(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_L g407 ( .A(n_327), .Y(n_407) );
INVx2_ASAP7_75t_SL g483 ( .A(n_328), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_330), .A2(n_385), .B1(n_387), .B2(n_391), .Y(n_384) );
AND2x2_ASAP7_75t_SL g330 ( .A(n_331), .B(n_332), .Y(n_330) );
AND2x2_ASAP7_75t_L g511 ( .A(n_331), .B(n_367), .Y(n_511) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_333), .B(n_377), .Y(n_456) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g422 ( .A(n_334), .B(n_370), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_335), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g365 ( .A(n_336), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g479 ( .A1(n_336), .A2(n_480), .B1(n_484), .B2(n_486), .C(n_488), .Y(n_479) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
AND2x2_ASAP7_75t_L g349 ( .A(n_337), .B(n_350), .Y(n_349) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_337), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_337), .B(n_380), .Y(n_435) );
INVx1_ASAP7_75t_SL g431 ( .A(n_338), .Y(n_431) );
AOI221xp5_ASAP7_75t_SL g459 ( .A1(n_338), .A2(n_349), .B1(n_460), .B2(n_461), .C(n_464), .Y(n_459) );
AOI322xp5_ASAP7_75t_L g492 ( .A1(n_338), .A2(n_410), .A3(n_437), .B1(n_493), .B2(n_495), .C1(n_496), .C2(n_499), .Y(n_492) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
BUFx2_ASAP7_75t_L g359 ( .A(n_339), .Y(n_359) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_340), .Y(n_351) );
INVx2_ASAP7_75t_L g409 ( .A(n_340), .Y(n_409) );
AND2x2_ASAP7_75t_L g450 ( .A(n_340), .B(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OA21x2_ASAP7_75t_SL g342 ( .A1(n_343), .A2(n_349), .B(n_352), .Y(n_342) );
AOI211xp5_ASAP7_75t_L g512 ( .A1(n_343), .A2(n_513), .B(n_514), .C(n_518), .Y(n_512) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
OR2x2_ASAP7_75t_L g401 ( .A(n_345), .B(n_363), .Y(n_401) );
OR2x2_ASAP7_75t_L g485 ( .A(n_345), .B(n_380), .Y(n_485) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g425 ( .A(n_347), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g503 ( .A(n_350), .Y(n_503) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g389 ( .A(n_351), .Y(n_389) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
OR2x2_ASAP7_75t_L g358 ( .A(n_354), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g393 ( .A(n_356), .B(n_394), .Y(n_393) );
OAI322xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .A3(n_363), .B1(n_365), .B2(n_366), .C1(n_371), .C2(n_373), .Y(n_357) );
INVx1_ASAP7_75t_L g399 ( .A(n_358), .Y(n_399) );
OR2x2_ASAP7_75t_L g371 ( .A(n_360), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_360), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g382 ( .A(n_364), .B(n_383), .Y(n_382) );
OAI32xp33_ASAP7_75t_L g427 ( .A1(n_364), .A2(n_428), .A3(n_431), .B1(n_432), .B2(n_433), .Y(n_427) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx2_ASAP7_75t_L g372 ( .A(n_367), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_367), .B(n_430), .Y(n_429) );
NOR2x1_ASAP7_75t_L g469 ( .A(n_367), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g493 ( .A(n_367), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g414 ( .A(n_368), .Y(n_414) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_372), .B(n_438), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_395), .Y(n_374) );
OAI21xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B(n_384), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_SL g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g444 ( .A(n_383), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_386), .A2(n_406), .B1(n_508), .B2(n_510), .Y(n_507) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g434 ( .A1(n_388), .A2(n_435), .B(n_436), .C(n_439), .Y(n_434) );
OR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx3_ASAP7_75t_L g516 ( .A(n_390), .Y(n_516) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g397 ( .A(n_394), .Y(n_397) );
AO21x1_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_398), .B(n_402), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g462 ( .A(n_397), .Y(n_462) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_403), .B(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g418 ( .A(n_405), .Y(n_418) );
OR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g475 ( .A(n_408), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
NOR3xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_434), .C(n_446), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
OAI21xp5_ASAP7_75t_SL g476 ( .A1(n_415), .A2(n_477), .B(n_478), .Y(n_476) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
INVx1_ASAP7_75t_L g451 ( .A(n_417), .Y(n_451) );
O2A1O1Ixp5_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_421), .B(n_423), .C(n_427), .Y(n_419) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_429), .Y(n_519) );
INVx2_ASAP7_75t_L g504 ( .A(n_432), .Y(n_504) );
AOI21xp33_ASAP7_75t_L g518 ( .A1(n_433), .A2(n_519), .B(n_520), .Y(n_518) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g498 ( .A(n_438), .Y(n_498) );
OAI31xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_442), .A3(n_443), .B(n_444), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g517 ( .A(n_445), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_452), .B(n_455), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
BUFx2_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g467 ( .A(n_450), .Y(n_467) );
AOI21xp33_ASAP7_75t_SL g514 ( .A1(n_452), .A2(n_515), .B(n_517), .Y(n_514) );
OR2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVx2_ASAP7_75t_L g482 ( .A(n_453), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_453), .B(n_473), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_453), .B(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g463 ( .A(n_454), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
NAND5xp2_ASAP7_75t_L g458 ( .A(n_459), .B(n_479), .C(n_492), .D(n_501), .E(n_512), .Y(n_458) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
OAI221xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_468), .B1(n_471), .B2(n_474), .C(n_476), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVxp67_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVxp67_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_505), .B(n_507), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
INVx1_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
INVxp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OAI222xp33_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_526), .B1(n_532), .B2(n_533), .C1(n_536), .C2(n_541), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
INVxp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
endmodule