module fake_jpeg_11130_n_603 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_603);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_603;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_3),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_SL g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_12),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_60),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_62),
.Y(n_189)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_24),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_64),
.B(n_77),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_65),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_66),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_67),
.Y(n_179)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_71),
.Y(n_159)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_72),
.Y(n_163)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_73),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_74),
.Y(n_195)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_75),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_20),
.B(n_18),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_24),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_79),
.B(n_81),
.Y(n_151)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_24),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_83),
.Y(n_181)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_85),
.Y(n_168)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_86),
.Y(n_171)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_87),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_88),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_20),
.B(n_16),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_89),
.B(n_91),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_90),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_24),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_92),
.Y(n_190)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_94),
.Y(n_194)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_95),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_96),
.Y(n_208)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_101),
.Y(n_196)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_102),
.Y(n_198)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_47),
.B(n_16),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_106),
.B(n_111),
.Y(n_187)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_47),
.B(n_49),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_49),
.B(n_0),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_115),
.B(n_117),
.Y(n_200)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_27),
.Y(n_116)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_26),
.B(n_59),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_30),
.Y(n_118)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_32),
.Y(n_119)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_32),
.Y(n_120)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_120),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_24),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_121),
.B(n_124),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

BUFx4f_ASAP7_75t_SL g128 ( 
.A(n_122),
.Y(n_128)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_42),
.Y(n_123)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_26),
.B(n_0),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_41),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g191 ( 
.A(n_126),
.Y(n_191)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_127),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_68),
.B(n_37),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_133),
.B(n_192),
.Y(n_227)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_62),
.B(n_36),
.Y(n_138)
);

NAND2xp33_ASAP7_75t_SL g219 ( 
.A(n_138),
.B(n_207),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_36),
.C(n_51),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_140),
.B(n_156),
.C(n_180),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_142),
.Y(n_221)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

BUFx2_ASAP7_75t_SL g230 ( 
.A(n_146),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_149),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_94),
.B(n_36),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_157),
.B(n_184),
.Y(n_235)
);

BUFx4f_ASAP7_75t_SL g165 ( 
.A(n_76),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_165),
.Y(n_258)
);

OR2x2_ASAP7_75t_SL g166 ( 
.A(n_86),
.B(n_41),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_166),
.B(n_35),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_113),
.B(n_44),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_167),
.B(n_0),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_72),
.A2(n_36),
.B1(n_35),
.B2(n_41),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_177),
.A2(n_73),
.B1(n_108),
.B2(n_114),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_116),
.B(n_102),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_82),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_93),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_186),
.B(n_204),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_71),
.B(n_31),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_98),
.B(n_55),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_205),
.Y(n_232)
);

BUFx4f_ASAP7_75t_SL g197 ( 
.A(n_95),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_197),
.Y(n_261)
);

NAND2x2_ASAP7_75t_L g201 ( 
.A(n_60),
.B(n_34),
.Y(n_201)
);

OA22x2_ASAP7_75t_L g238 ( 
.A1(n_201),
.A2(n_105),
.B1(n_100),
.B2(n_88),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_103),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_112),
.B(n_31),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_83),
.B(n_51),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_61),
.A2(n_57),
.B1(n_52),
.B2(n_25),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_210),
.A2(n_57),
.B1(n_52),
.B2(n_25),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_213),
.Y(n_302)
);

INVx11_ASAP7_75t_L g214 ( 
.A(n_147),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_214),
.Y(n_334)
);

CKINVDCx12_ASAP7_75t_R g215 ( 
.A(n_132),
.Y(n_215)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_215),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_216),
.Y(n_293)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_217),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_90),
.B1(n_66),
.B2(n_74),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_218),
.A2(n_233),
.B1(n_257),
.B2(n_272),
.Y(n_289)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_220),
.Y(n_305)
);

CKINVDCx12_ASAP7_75t_R g222 ( 
.A(n_154),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_222),
.Y(n_292)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_144),
.Y(n_223)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_223),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_224),
.Y(n_301)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_160),
.Y(n_225)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_225),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_228),
.A2(n_263),
.B1(n_264),
.B2(n_274),
.Y(n_328)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_153),
.Y(n_229)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_229),
.Y(n_314)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_202),
.B(n_172),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_231),
.B(n_266),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_131),
.A2(n_130),
.B1(n_145),
.B2(n_173),
.Y(n_233)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_234),
.Y(n_339)
);

O2A1O1Ixp33_ASAP7_75t_SL g236 ( 
.A1(n_207),
.A2(n_60),
.B(n_67),
.C(n_99),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_236),
.B(n_250),
.Y(n_317)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_237),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_238),
.B(n_240),
.Y(n_286)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_136),
.Y(n_239)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_239),
.Y(n_327)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_168),
.Y(n_241)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_241),
.Y(n_330)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_136),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_242),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_174),
.B(n_44),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_244),
.B(n_270),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_181),
.Y(n_246)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_246),
.Y(n_340)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_151),
.Y(n_247)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_247),
.Y(n_311)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_151),
.Y(n_248)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_248),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_249),
.B(n_265),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_142),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_170),
.Y(n_251)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_251),
.Y(n_294)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_175),
.Y(n_252)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_252),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_200),
.B(n_58),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_253),
.B(n_267),
.Y(n_287)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_141),
.Y(n_254)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_254),
.Y(n_296)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_169),
.Y(n_255)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_255),
.Y(n_306)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_185),
.Y(n_256)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_256),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_201),
.A2(n_65),
.B1(n_120),
.B2(n_119),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_200),
.A2(n_29),
.B(n_37),
.C(n_59),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_259),
.B(n_273),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_164),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_260),
.B(n_262),
.Y(n_320)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_143),
.A2(n_67),
.B1(n_35),
.B2(n_57),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_189),
.A2(n_25),
.B1(n_125),
.B2(n_55),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_191),
.Y(n_265)
);

AND2x2_ASAP7_75t_SL g266 ( 
.A(n_134),
.B(n_137),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_187),
.B(n_58),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_196),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_268),
.B(n_269),
.Y(n_321)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_182),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_150),
.B(n_50),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_187),
.B(n_50),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_271),
.B(n_277),
.Y(n_313)
);

OAI22xp33_ASAP7_75t_L g272 ( 
.A1(n_210),
.A2(n_46),
.B1(n_40),
.B2(n_38),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_178),
.A2(n_46),
.B(n_40),
.C(n_38),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_164),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_149),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_275),
.B(n_276),
.Y(n_325)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_129),
.Y(n_276)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_148),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_278),
.B(n_279),
.Y(n_329)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_135),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_191),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_280),
.B(n_281),
.Y(n_337)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_206),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_171),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_282),
.B(n_284),
.Y(n_338)
);

AND2x2_ASAP7_75t_SL g283 ( 
.A(n_178),
.B(n_2),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_283),
.B(n_128),
.C(n_4),
.Y(n_341)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_183),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_164),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_285),
.A2(n_209),
.B1(n_161),
.B2(n_179),
.Y(n_315)
);

AO22x1_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_177),
.B1(n_212),
.B2(n_167),
.Y(n_290)
);

OA22x2_ASAP7_75t_SL g381 ( 
.A1(n_290),
.A2(n_190),
.B1(n_5),
.B2(n_6),
.Y(n_381)
);

OR2x6_ASAP7_75t_L g300 ( 
.A(n_219),
.B(n_146),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_300),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_226),
.B(n_150),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_307),
.B(n_260),
.C(n_128),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_240),
.A2(n_199),
.B1(n_198),
.B2(n_159),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_308),
.A2(n_315),
.B1(n_324),
.B2(n_326),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_235),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_309),
.B(n_332),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_232),
.B(n_162),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_333),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_238),
.A2(n_156),
.B1(n_180),
.B2(n_211),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_316),
.A2(n_335),
.B1(n_280),
.B2(n_265),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_283),
.A2(n_165),
.B(n_197),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_323),
.A2(n_246),
.B(n_208),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_264),
.A2(n_159),
.B1(n_203),
.B2(n_195),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_228),
.A2(n_211),
.B1(n_203),
.B2(n_195),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_243),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_227),
.B(n_273),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_238),
.A2(n_158),
.B1(n_152),
.B2(n_139),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_231),
.B(n_158),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_336),
.B(n_341),
.Y(n_358)
);

INVx8_ASAP7_75t_L g342 ( 
.A(n_303),
.Y(n_342)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_342),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_317),
.A2(n_257),
.B1(n_218),
.B2(n_263),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_343),
.A2(n_347),
.B1(n_354),
.B2(n_360),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_303),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_344),
.Y(n_385)
);

BUFx12f_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_345),
.B(n_359),
.Y(n_387)
);

NAND2x1_ASAP7_75t_L g346 ( 
.A(n_300),
.B(n_236),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_346),
.A2(n_376),
.B(n_379),
.Y(n_409)
);

OAI22xp33_ASAP7_75t_L g347 ( 
.A1(n_328),
.A2(n_224),
.B1(n_216),
.B2(n_213),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_333),
.B(n_259),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_348),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_286),
.B(n_266),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_349),
.B(n_361),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_296),
.A2(n_252),
.B1(n_258),
.B2(n_278),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_350),
.A2(n_381),
.B1(n_334),
.B2(n_340),
.Y(n_420)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_331),
.Y(n_351)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_351),
.Y(n_388)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_331),
.Y(n_353)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

INVx5_ASAP7_75t_L g355 ( 
.A(n_339),
.Y(n_355)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_355),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_312),
.B(n_220),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_368),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_319),
.B(n_245),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_299),
.A2(n_274),
.B1(n_285),
.B2(n_239),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_286),
.B(n_323),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_286),
.A2(n_242),
.B1(n_152),
.B2(n_254),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_363),
.A2(n_362),
.B1(n_302),
.B2(n_295),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_311),
.B(n_221),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_364),
.B(n_365),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_318),
.B(n_237),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_325),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_366),
.B(n_370),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_290),
.A2(n_217),
.B1(n_261),
.B2(n_258),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_367),
.A2(n_373),
.B1(n_376),
.B2(n_370),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_299),
.B(n_261),
.Y(n_368)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_339),
.Y(n_369)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_300),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_378),
.C(n_382),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_304),
.B(n_3),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_372),
.B(n_383),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_300),
.A2(n_230),
.B1(n_161),
.B2(n_209),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_292),
.B(n_251),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_374),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_337),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_375),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_288),
.B(n_208),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_306),
.Y(n_377)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_377),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_307),
.B(n_214),
.C(n_234),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_304),
.B(n_190),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_287),
.B(n_313),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_300),
.A2(n_4),
.B(n_5),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_384),
.A2(n_346),
.B(n_379),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_352),
.A2(n_290),
.B1(n_289),
.B2(n_288),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_389),
.A2(n_392),
.B1(n_404),
.B2(n_405),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_357),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_394),
.B(n_402),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_397),
.B(n_373),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_356),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_352),
.A2(n_288),
.B1(n_341),
.B2(n_295),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_362),
.A2(n_327),
.B1(n_296),
.B2(n_329),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_380),
.A2(n_368),
.B1(n_363),
.B2(n_381),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_406),
.B(n_417),
.Y(n_427)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_351),
.Y(n_407)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_407),
.Y(n_421)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_353),
.Y(n_411)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_411),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_380),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_412),
.B(n_345),
.Y(n_431)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_377),
.Y(n_414)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_414),
.Y(n_440)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_355),
.Y(n_416)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_416),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_381),
.A2(n_327),
.B1(n_302),
.B2(n_301),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_418),
.Y(n_444)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_369),
.Y(n_419)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_419),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_420),
.A2(n_345),
.B1(n_334),
.B2(n_347),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_390),
.A2(n_381),
.B1(n_348),
.B2(n_384),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_422),
.A2(n_426),
.B1(n_428),
.B2(n_429),
.Y(n_469)
);

INVx13_ASAP7_75t_L g423 ( 
.A(n_412),
.Y(n_423)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_423),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_396),
.B(n_378),
.C(n_382),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_424),
.B(n_415),
.C(n_406),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_390),
.A2(n_358),
.B1(n_343),
.B2(n_371),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_402),
.A2(n_361),
.B1(n_346),
.B2(n_349),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_386),
.B(n_401),
.Y(n_430)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_430),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_431),
.B(n_436),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_386),
.B(n_366),
.Y(n_433)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_433),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_434),
.A2(n_395),
.B1(n_399),
.B2(n_400),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_394),
.B(n_372),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_442),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_393),
.B(n_338),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_397),
.A2(n_361),
.B1(n_349),
.B2(n_376),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_438),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_389),
.A2(n_342),
.B1(n_344),
.B2(n_293),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_387),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_449),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_401),
.B(n_321),
.Y(n_441)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_441),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_387),
.B(n_345),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_418),
.A2(n_340),
.B(n_294),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_445),
.A2(n_414),
.B(n_403),
.Y(n_464)
);

CKINVDCx10_ASAP7_75t_R g446 ( 
.A(n_400),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_446),
.Y(n_478)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_388),
.Y(n_448)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_448),
.Y(n_470)
);

OAI21xp33_ASAP7_75t_SL g449 ( 
.A1(n_409),
.A2(n_294),
.B(n_322),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_409),
.A2(n_320),
.B(n_322),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_450),
.A2(n_398),
.B(n_413),
.Y(n_454)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_388),
.Y(n_451)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_451),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_396),
.A2(n_301),
.B1(n_293),
.B2(n_330),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_452),
.B(n_404),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_454),
.A2(n_423),
.B1(n_391),
.B2(n_407),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_431),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_482),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_439),
.Y(n_461)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_461),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_464),
.A2(n_450),
.B(n_445),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_465),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_433),
.B(n_403),
.Y(n_466)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_466),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_424),
.B(n_413),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_468),
.B(n_483),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_SL g471 ( 
.A1(n_444),
.A2(n_393),
.B1(n_416),
.B2(n_419),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_471),
.A2(n_458),
.B1(n_478),
.B2(n_434),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_472),
.A2(n_429),
.B1(n_449),
.B2(n_438),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_473),
.B(n_437),
.C(n_452),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_435),
.B(n_410),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_474),
.B(n_475),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_425),
.B(n_398),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_425),
.B(n_415),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_476),
.B(n_480),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_430),
.B(n_411),
.Y(n_477)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_477),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_436),
.B(n_330),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_421),
.Y(n_481)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_481),
.Y(n_506)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_421),
.Y(n_482)
);

NOR4xp25_ASAP7_75t_L g483 ( 
.A(n_441),
.B(n_405),
.C(n_392),
.D(n_417),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_485),
.A2(n_505),
.B1(n_472),
.B2(n_464),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_432),
.Y(n_487)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_487),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_462),
.B(n_432),
.Y(n_488)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_488),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_457),
.A2(n_469),
.B1(n_453),
.B2(n_462),
.Y(n_490)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_490),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_426),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_492),
.B(n_502),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_508),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_463),
.B(n_446),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_497),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_467),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_498),
.B(n_501),
.C(n_478),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_469),
.A2(n_453),
.B1(n_427),
.B2(n_442),
.Y(n_499)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_499),
.Y(n_519)
);

XNOR2x1_ASAP7_75t_L g524 ( 
.A(n_500),
.B(n_510),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_468),
.B(n_428),
.C(n_427),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_454),
.B(n_422),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_465),
.B(n_429),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_503),
.B(n_459),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_456),
.A2(n_459),
.B1(n_460),
.B2(n_483),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_463),
.A2(n_451),
.B1(n_448),
.B2(n_440),
.Y(n_507)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_507),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_456),
.A2(n_429),
.B1(n_440),
.B2(n_443),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_516),
.A2(n_500),
.B1(n_493),
.B2(n_508),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_486),
.B(n_460),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_517),
.B(n_531),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_489),
.B(n_467),
.Y(n_518)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_518),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_521),
.B(n_523),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_492),
.B(n_477),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_525),
.B(n_528),
.C(n_529),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_505),
.B(n_461),
.Y(n_526)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_526),
.Y(n_550)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_484),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_527),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_498),
.B(n_461),
.C(n_455),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_501),
.B(n_455),
.C(n_447),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_487),
.B(n_481),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_530),
.Y(n_537)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_484),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_502),
.B(n_482),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_532),
.B(n_504),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_519),
.A2(n_510),
.B1(n_494),
.B2(n_495),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_535),
.A2(n_470),
.B1(n_479),
.B2(n_443),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_529),
.B(n_503),
.C(n_509),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_536),
.B(n_541),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_539),
.A2(n_514),
.B1(n_512),
.B2(n_524),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_511),
.A2(n_495),
.B(n_494),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_540),
.A2(n_545),
.B(n_506),
.Y(n_564)
);

INVxp33_ASAP7_75t_L g541 ( 
.A(n_513),
.Y(n_541)
);

AOI21xp33_ASAP7_75t_L g543 ( 
.A1(n_511),
.A2(n_488),
.B(n_491),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_543),
.B(n_549),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_544),
.B(n_532),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_516),
.A2(n_515),
.B(n_522),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_525),
.B(n_509),
.C(n_491),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_547),
.B(n_548),
.C(n_536),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_528),
.B(n_504),
.C(n_447),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_523),
.B(n_408),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_551),
.B(n_560),
.Y(n_570)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_538),
.Y(n_552)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_552),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_SL g553 ( 
.A(n_547),
.B(n_520),
.Y(n_553)
);

NOR2xp67_ASAP7_75t_SL g568 ( 
.A(n_553),
.B(n_556),
.Y(n_568)
);

FAx1_ASAP7_75t_SL g555 ( 
.A(n_540),
.B(n_521),
.CI(n_530),
.CON(n_555),
.SN(n_555)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_555),
.B(n_558),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_SL g556 ( 
.A(n_542),
.B(n_520),
.Y(n_556)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_557),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_533),
.B(n_548),
.C(n_542),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_541),
.B(n_408),
.Y(n_559)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_559),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_534),
.A2(n_506),
.B1(n_524),
.B2(n_479),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_562),
.B(n_565),
.C(n_537),
.Y(n_571)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_546),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_563),
.A2(n_564),
.B(n_537),
.Y(n_567)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_567),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_558),
.B(n_533),
.C(n_545),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_569),
.B(n_572),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_571),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_551),
.B(n_550),
.C(n_535),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_561),
.B(n_399),
.C(n_395),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_574),
.B(n_576),
.C(n_565),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_553),
.B(n_470),
.C(n_391),
.Y(n_576)
);

OAI322xp33_ASAP7_75t_L g578 ( 
.A1(n_566),
.A2(n_554),
.A3(n_557),
.B1(n_555),
.B2(n_556),
.C1(n_564),
.C2(n_560),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_578),
.A2(n_582),
.B1(n_310),
.B2(n_297),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_577),
.B(n_555),
.Y(n_579)
);

AO21x1_ASAP7_75t_L g592 ( 
.A1(n_579),
.A2(n_314),
.B(n_298),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_581),
.B(n_310),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_575),
.A2(n_423),
.B1(n_385),
.B2(n_305),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_573),
.A2(n_569),
.B1(n_576),
.B2(n_570),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_583),
.B(n_584),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_570),
.B(n_385),
.C(n_306),
.Y(n_584)
);

AOI322xp5_ASAP7_75t_L g588 ( 
.A1(n_585),
.A2(n_568),
.A3(n_385),
.B1(n_314),
.B2(n_298),
.C1(n_291),
.C2(n_305),
.Y(n_588)
);

AOI21xp33_ASAP7_75t_L g593 ( 
.A1(n_588),
.A2(n_591),
.B(n_579),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_589),
.B(n_590),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_580),
.B(n_297),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_592),
.B(n_584),
.C(n_586),
.Y(n_595)
);

O2A1O1Ixp33_ASAP7_75t_L g598 ( 
.A1(n_593),
.A2(n_595),
.B(n_596),
.C(n_6),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_591),
.B(n_586),
.Y(n_596)
);

AOI322xp5_ASAP7_75t_L g597 ( 
.A1(n_594),
.A2(n_582),
.A3(n_587),
.B1(n_581),
.B2(n_10),
.C1(n_6),
.C2(n_14),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_597),
.B(n_598),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_SL g600 ( 
.A1(n_599),
.A2(n_6),
.B(n_8),
.Y(n_600)
);

O2A1O1Ixp33_ASAP7_75t_L g601 ( 
.A1(n_600),
.A2(n_8),
.B(n_9),
.C(n_11),
.Y(n_601)
);

O2A1O1Ixp33_ASAP7_75t_SL g602 ( 
.A1(n_601),
.A2(n_8),
.B(n_9),
.C(n_14),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_602),
.A2(n_14),
.B(n_384),
.Y(n_603)
);


endmodule