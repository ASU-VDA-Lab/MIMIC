module fake_ibex_1432_n_1561 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_247, n_274, n_55, n_130, n_275, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_267, n_268, n_8, n_118, n_224, n_273, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_264, n_124, n_37, n_256, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_263, n_27, n_165, n_242, n_278, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_262, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_14, n_0, n_239, n_94, n_134, n_12, n_266, n_42, n_77, n_112, n_257, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_258, n_80, n_172, n_215, n_250, n_279, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_261, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_281, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_260, n_99, n_280, n_269, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_270, n_230, n_96, n_185, n_271, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_265, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_259, n_132, n_174, n_276, n_277, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_272, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1561);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_247;
input n_274;
input n_55;
input n_130;
input n_275;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_267;
input n_268;
input n_8;
input n_118;
input n_224;
input n_273;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_264;
input n_124;
input n_37;
input n_256;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_263;
input n_27;
input n_165;
input n_242;
input n_278;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_262;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_266;
input n_42;
input n_77;
input n_112;
input n_257;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_258;
input n_80;
input n_172;
input n_215;
input n_250;
input n_279;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_261;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_281;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_260;
input n_99;
input n_280;
input n_269;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_270;
input n_230;
input n_96;
input n_185;
input n_271;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_265;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_259;
input n_132;
input n_174;
input n_276;
input n_277;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_272;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1561;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_1509;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_1506;
wire n_881;
wire n_734;
wire n_1558;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_1434;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1531;
wire n_1332;
wire n_482;
wire n_282;
wire n_1424;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1521;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1477;
wire n_1364;
wire n_1540;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1522;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_1545;
wire n_351;
wire n_456;
wire n_1471;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1470;
wire n_444;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_650;
wire n_409;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_291;
wire n_318;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_303;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1560;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1497;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_1458;
wire n_1460;
wire n_326;
wire n_1340;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_1538;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_300;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_480;
wire n_1057;
wire n_354;
wire n_1473;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1501;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_1513;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_284;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_387;
wire n_688;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1369;
wire n_1297;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_335;
wire n_1499;
wire n_1500;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_305;
wire n_566;
wire n_581;
wire n_416;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_537;
wire n_1113;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1559;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_84),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_3),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_270),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_210),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_278),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_78),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_105),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_152),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_136),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_1),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_15),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_204),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_249),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_238),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_252),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_21),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_267),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_164),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_160),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_49),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_273),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_272),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_16),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_100),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_122),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_181),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_143),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_170),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_90),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_183),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_201),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_151),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_159),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_108),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_167),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_250),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_179),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_202),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_123),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_206),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_156),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_222),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_203),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_142),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_41),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_128),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_53),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_274),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_26),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_105),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_262),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_243),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_71),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_32),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_114),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_217),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_245),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_161),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_197),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_244),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_166),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_42),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_113),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_255),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_173),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_54),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_195),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_263),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_62),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_168),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_264),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_52),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_118),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_246),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_81),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_256),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_3),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_171),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_220),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_23),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_2),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_241),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_239),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_182),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_231),
.B(n_49),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_72),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_94),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_124),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_135),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_91),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_118),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_200),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_240),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_247),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_17),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_225),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_169),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_251),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_184),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_198),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_261),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_218),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_237),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_212),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_139),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_269),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_83),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_122),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_125),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_101),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_32),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_59),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_119),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_157),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_103),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_130),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_50),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_276),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_74),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_90),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_77),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_258),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_10),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_29),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_129),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_148),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_109),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_248),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_257),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_209),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_95),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_208),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_277),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_38),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_266),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_213),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_205),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_136),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_39),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_26),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_253),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_279),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_180),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_95),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_77),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_275),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_199),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_196),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_46),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_42),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_28),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_216),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_130),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_18),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_29),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_107),
.Y(n_437)
);

BUFx10_ASAP7_75t_L g438 ( 
.A(n_74),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_271),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_176),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_28),
.Y(n_441)
);

NOR2xp67_ASAP7_75t_L g442 ( 
.A(n_174),
.B(n_132),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_35),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_162),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_91),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_227),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_65),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_137),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_140),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_21),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_12),
.Y(n_451)
);

BUFx10_ASAP7_75t_L g452 ( 
.A(n_215),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_207),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_43),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_265),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_175),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_99),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_146),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_172),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_79),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_224),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_281),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_75),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_35),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_133),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_165),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_11),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_81),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_185),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_223),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_163),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_101),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_5),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_117),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_228),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_325),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_340),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_340),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_340),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_299),
.B(n_141),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_335),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_402),
.A2(n_4),
.B1(n_0),
.B2(n_2),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_319),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_319),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_438),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_407),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_335),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_322),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_407),
.Y(n_489)
);

OA21x2_ASAP7_75t_L g490 ( 
.A1(n_322),
.A2(n_145),
.B(n_144),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_335),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_376),
.A2(n_5),
.B1(n_0),
.B2(n_4),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_357),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_283),
.B(n_6),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_332),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_422),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_325),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_327),
.B(n_6),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_438),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_438),
.Y(n_500)
);

BUFx12f_ASAP7_75t_L g501 ( 
.A(n_452),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_297),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_449),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_433),
.B(n_7),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_408),
.B(n_7),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_297),
.Y(n_506)
);

OAI22x1_ASAP7_75t_SL g507 ( 
.A1(n_431),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_301),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_365),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_365),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_297),
.Y(n_511)
);

BUFx12f_ASAP7_75t_L g512 ( 
.A(n_452),
.Y(n_512)
);

INVx6_ASAP7_75t_L g513 ( 
.A(n_452),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_344),
.B(n_8),
.Y(n_514)
);

XNOR2x2_ASAP7_75t_L g515 ( 
.A(n_291),
.B(n_9),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_457),
.B(n_433),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_344),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_297),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_425),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_425),
.B(n_426),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_426),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_412),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_282),
.B(n_11),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_370),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_412),
.B(n_12),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_370),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_443),
.B(n_13),
.Y(n_527)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_337),
.Y(n_528)
);

INVxp33_ASAP7_75t_SL g529 ( 
.A(n_305),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_395),
.A2(n_444),
.B(n_399),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_290),
.B(n_13),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_360),
.B(n_14),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_360),
.B(n_14),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_395),
.B(n_16),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_304),
.Y(n_535)
);

OAI22x1_ASAP7_75t_R g536 ( 
.A1(n_431),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_305),
.A2(n_22),
.B1(n_19),
.B2(n_20),
.Y(n_537)
);

OAI22x1_ASAP7_75t_L g538 ( 
.A1(n_306),
.A2(n_23),
.B1(n_20),
.B2(n_22),
.Y(n_538)
);

AND2x6_ASAP7_75t_L g539 ( 
.A(n_409),
.B(n_147),
.Y(n_539)
);

OAI22x1_ASAP7_75t_L g540 ( 
.A1(n_306),
.A2(n_27),
.B1(n_24),
.B2(n_25),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_310),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_310),
.A2(n_31),
.B1(n_27),
.B2(n_30),
.Y(n_542)
);

CKINVDCx8_ASAP7_75t_R g543 ( 
.A(n_320),
.Y(n_543)
);

BUFx12f_ASAP7_75t_L g544 ( 
.A(n_296),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_370),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_320),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_284),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_460),
.B(n_30),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_329),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_288),
.B(n_31),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_292),
.B(n_33),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_315),
.Y(n_552)
);

INVx5_ASAP7_75t_L g553 ( 
.A(n_409),
.Y(n_553)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_399),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_396),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_444),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_460),
.B(n_33),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_396),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_285),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_289),
.Y(n_560)
);

BUFx12f_ASAP7_75t_L g561 ( 
.A(n_296),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_295),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_331),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_463),
.A2(n_37),
.B1(n_34),
.B2(n_36),
.Y(n_564)
);

CKINVDCx16_ASAP7_75t_R g565 ( 
.A(n_448),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_463),
.A2(n_39),
.B1(n_36),
.B2(n_38),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_329),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_530),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_483),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_514),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_499),
.B(n_300),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_503),
.B(n_465),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_513),
.B(n_294),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_513),
.Y(n_574)
);

CKINVDCx6p67_ASAP7_75t_R g575 ( 
.A(n_544),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_529),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_514),
.Y(n_577)
);

NOR2x1p5_ASAP7_75t_L g578 ( 
.A(n_501),
.B(n_465),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_499),
.B(n_300),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_513),
.B(n_342),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_500),
.B(n_302),
.Y(n_581)
);

BUFx6f_ASAP7_75t_SL g582 ( 
.A(n_514),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_500),
.B(n_302),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_487),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_541),
.B(n_467),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_485),
.B(n_303),
.Y(n_586)
);

BUFx6f_ASAP7_75t_SL g587 ( 
.A(n_532),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_529),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_547),
.B(n_298),
.Y(n_589)
);

NAND3xp33_ASAP7_75t_L g590 ( 
.A(n_496),
.B(n_473),
.C(n_472),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_477),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_520),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_547),
.B(n_501),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_512),
.B(n_303),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_483),
.Y(n_595)
);

AND2x2_ASAP7_75t_SL g596 ( 
.A(n_480),
.B(n_366),
.Y(n_596)
);

BUFx6f_ASAP7_75t_SL g597 ( 
.A(n_532),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_512),
.B(n_307),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_484),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_477),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_516),
.B(n_307),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_487),
.B(n_541),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_476),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_484),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_478),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_488),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_546),
.B(n_472),
.Y(n_607)
);

NOR2x1_ASAP7_75t_L g608 ( 
.A(n_508),
.B(n_309),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_520),
.Y(n_609)
);

BUFx10_ASAP7_75t_L g610 ( 
.A(n_495),
.Y(n_610)
);

NAND2x1_ASAP7_75t_L g611 ( 
.A(n_532),
.B(n_533),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_SL g612 ( 
.A(n_523),
.B(n_363),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_478),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_520),
.B(n_308),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_493),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_479),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_546),
.B(n_473),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_543),
.B(n_308),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_479),
.Y(n_619)
);

NAND3xp33_ASAP7_75t_L g620 ( 
.A(n_504),
.B(n_474),
.C(n_326),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_479),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_533),
.B(n_311),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_479),
.Y(n_623)
);

INVxp33_ASAP7_75t_L g624 ( 
.A(n_548),
.Y(n_624)
);

INVx6_ASAP7_75t_L g625 ( 
.A(n_554),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_493),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_525),
.Y(n_627)
);

BUFx6f_ASAP7_75t_SL g628 ( 
.A(n_533),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_517),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_494),
.B(n_474),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_544),
.B(n_312),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_486),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_486),
.Y(n_633)
);

BUFx10_ASAP7_75t_L g634 ( 
.A(n_504),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_561),
.B(n_312),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_521),
.B(n_313),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_535),
.B(n_314),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_481),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_498),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_491),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_489),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_561),
.B(n_314),
.Y(n_642)
);

INVxp33_ASAP7_75t_L g643 ( 
.A(n_557),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_489),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_531),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_490),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_502),
.Y(n_647)
);

CKINVDCx6p67_ASAP7_75t_R g648 ( 
.A(n_565),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_502),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_552),
.B(n_316),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_531),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_502),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_506),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_505),
.B(n_362),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_497),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_506),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_528),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_506),
.Y(n_658)
);

NOR2x1p5_ASAP7_75t_L g659 ( 
.A(n_549),
.B(n_336),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_563),
.B(n_318),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_509),
.Y(n_661)
);

AOI21x1_ASAP7_75t_L g662 ( 
.A1(n_534),
.A2(n_321),
.B(n_317),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_559),
.B(n_560),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_511),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_511),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_522),
.B(n_519),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_518),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_518),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_559),
.B(n_318),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_518),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_510),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_527),
.B(n_372),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_490),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_510),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_518),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_560),
.B(n_323),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_556),
.Y(n_677)
);

AO21x2_ASAP7_75t_L g678 ( 
.A1(n_534),
.A2(n_551),
.B(n_550),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_562),
.B(n_323),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_562),
.B(n_522),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_549),
.Y(n_681)
);

AND3x2_ASAP7_75t_L g682 ( 
.A(n_536),
.B(n_417),
.C(n_353),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_524),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_556),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_528),
.B(n_324),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_524),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_554),
.B(n_324),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_524),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_539),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_526),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_526),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_555),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_526),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_567),
.B(n_405),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_526),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_555),
.Y(n_696)
);

BUFx10_ASAP7_75t_L g697 ( 
.A(n_539),
.Y(n_697)
);

CKINVDCx6p67_ASAP7_75t_R g698 ( 
.A(n_538),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_567),
.Y(n_699)
);

INVx8_ASAP7_75t_L g700 ( 
.A(n_553),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_553),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_545),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_515),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_639),
.B(n_380),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_602),
.B(n_287),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_614),
.B(n_459),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_636),
.B(n_637),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_571),
.B(n_462),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_650),
.B(n_470),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_579),
.B(n_470),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_696),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_592),
.Y(n_712)
);

NAND3xp33_ASAP7_75t_L g713 ( 
.A(n_590),
.B(n_542),
.C(n_537),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_585),
.B(n_482),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_581),
.B(n_475),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_602),
.A2(n_364),
.B1(n_373),
.B2(n_363),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_576),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_650),
.B(n_475),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_660),
.B(n_286),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_592),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_660),
.B(n_293),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_611),
.A2(n_354),
.B(n_358),
.C(n_350),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_588),
.B(n_328),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_585),
.Y(n_724)
);

NOR2x1p5_ASAP7_75t_L g725 ( 
.A(n_575),
.B(n_507),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_617),
.Y(n_726)
);

NOR2xp67_ASAP7_75t_L g727 ( 
.A(n_572),
.B(n_540),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_617),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_655),
.B(n_341),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_630),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_609),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_648),
.Y(n_732)
);

AO221x1_ASAP7_75t_L g733 ( 
.A1(n_703),
.A2(n_566),
.B1(n_564),
.B2(n_381),
.C(n_386),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_584),
.A2(n_373),
.B1(n_381),
.B2(n_364),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_609),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_630),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_681),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_666),
.Y(n_738)
);

OR2x6_ASAP7_75t_L g739 ( 
.A(n_578),
.B(n_361),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_661),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_587),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_669),
.B(n_348),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_583),
.B(n_601),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_666),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_620),
.B(n_333),
.Y(n_745)
);

INVx8_ASAP7_75t_L g746 ( 
.A(n_582),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_676),
.B(n_679),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_593),
.B(n_492),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_645),
.B(n_338),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_629),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_651),
.B(n_339),
.Y(n_751)
);

NOR2x1_ASAP7_75t_L g752 ( 
.A(n_594),
.B(n_598),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_661),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_607),
.B(n_375),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_672),
.B(n_334),
.C(n_330),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_589),
.B(n_377),
.Y(n_756)
);

INVx8_ASAP7_75t_L g757 ( 
.A(n_582),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_698),
.A2(n_386),
.B1(n_454),
.B2(n_448),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_573),
.B(n_384),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_624),
.B(n_343),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_580),
.B(n_385),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_684),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_689),
.Y(n_763)
);

INVxp33_ASAP7_75t_L g764 ( 
.A(n_694),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_627),
.B(n_685),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_622),
.B(n_403),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_684),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_569),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_570),
.A2(n_368),
.B1(n_389),
.B2(n_367),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_603),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_634),
.B(n_410),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_634),
.B(n_411),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_634),
.B(n_413),
.Y(n_773)
);

INVxp33_ASAP7_75t_L g774 ( 
.A(n_694),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_624),
.B(n_643),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_569),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_643),
.B(n_416),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_703),
.A2(n_394),
.B(n_398),
.C(n_391),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_570),
.B(n_418),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_595),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_577),
.B(n_423),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_672),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_577),
.B(n_424),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_577),
.A2(n_400),
.B1(n_406),
.B2(n_401),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_654),
.B(n_347),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_699),
.B(n_356),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_608),
.B(n_427),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_611),
.B(n_428),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_603),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_595),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_638),
.B(n_640),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_574),
.B(n_439),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_574),
.B(n_440),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_599),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_599),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_678),
.B(n_446),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_604),
.Y(n_797)
);

NOR3xp33_ASAP7_75t_L g798 ( 
.A(n_612),
.B(n_371),
.C(n_369),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_678),
.B(n_453),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_678),
.B(n_458),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_604),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_625),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_586),
.B(n_345),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_680),
.B(n_388),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_606),
.Y(n_805)
);

AOI22x1_ASAP7_75t_L g806 ( 
.A1(n_568),
.A2(n_349),
.B1(n_351),
.B2(n_346),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_615),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_596),
.A2(n_582),
.B1(n_597),
.B2(n_587),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_587),
.B(n_352),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_596),
.A2(n_392),
.B1(n_393),
.B2(n_390),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_626),
.B(n_397),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_597),
.A2(n_419),
.B1(n_421),
.B2(n_404),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_697),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_610),
.B(n_434),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_597),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_697),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_SL g817 ( 
.A1(n_682),
.A2(n_464),
.B1(n_468),
.B2(n_454),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_671),
.B(n_450),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_628),
.A2(n_451),
.B1(n_415),
.B2(n_420),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_674),
.B(n_355),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_659),
.B(n_430),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_674),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_677),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_628),
.A2(n_435),
.B1(n_437),
.B2(n_432),
.Y(n_824)
);

NAND2xp33_ASAP7_75t_SL g825 ( 
.A(n_631),
.B(n_464),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_687),
.B(n_359),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_648),
.Y(n_827)
);

NAND2x1p5_ASAP7_75t_L g828 ( 
.A(n_635),
.B(n_441),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_663),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_610),
.B(n_468),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_701),
.Y(n_831)
);

O2A1O1Ixp5_ASAP7_75t_L g832 ( 
.A1(n_662),
.A2(n_378),
.B(n_379),
.C(n_374),
.Y(n_832)
);

NAND3xp33_ASAP7_75t_SL g833 ( 
.A(n_642),
.B(n_383),
.C(n_382),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_662),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_692),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_657),
.Y(n_836)
);

BUFx12f_ASAP7_75t_SL g837 ( 
.A(n_575),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_618),
.B(n_387),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_657),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_646),
.B(n_414),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_698),
.A2(n_447),
.B1(n_445),
.B2(n_436),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_646),
.B(n_429),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_700),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_673),
.B(n_442),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_647),
.A2(n_456),
.B1(n_461),
.B2(n_455),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_649),
.B(n_466),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_649),
.B(n_469),
.Y(n_847)
);

BUFx5_ASAP7_75t_L g848 ( 
.A(n_641),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_641),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_652),
.B(n_471),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_720),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_717),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_713),
.A2(n_436),
.B1(n_558),
.B2(n_545),
.Y(n_853)
);

A2O1A1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_840),
.A2(n_436),
.B(n_558),
.C(n_545),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_717),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_707),
.B(n_40),
.Y(n_856)
);

NOR2x2_ASAP7_75t_L g857 ( 
.A(n_739),
.B(n_41),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_724),
.B(n_43),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_737),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_724),
.B(n_44),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_764),
.B(n_44),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_747),
.B(n_728),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_704),
.B(n_45),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_704),
.B(n_45),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_732),
.B(n_46),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_730),
.B(n_47),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_774),
.B(n_47),
.Y(n_867)
);

A2O1A1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_840),
.A2(n_656),
.B(n_658),
.C(n_653),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_832),
.A2(n_834),
.B(n_842),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_765),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_837),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_796),
.A2(n_800),
.B(n_799),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_709),
.B(n_48),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_842),
.A2(n_600),
.B(n_591),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_736),
.B(n_50),
.Y(n_875)
);

INVx1_ASAP7_75t_SL g876 ( 
.A(n_723),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_738),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_791),
.A2(n_613),
.B(n_605),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_827),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_808),
.B(n_641),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_786),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_779),
.A2(n_613),
.B(n_605),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_718),
.B(n_51),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_SL g884 ( 
.A(n_746),
.B(n_664),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_778),
.A2(n_667),
.B(n_668),
.C(n_665),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_785),
.B(n_51),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_781),
.A2(n_619),
.B(n_616),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_726),
.B(n_775),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_783),
.A2(n_623),
.B(n_621),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_744),
.B(n_722),
.Y(n_890)
);

NOR2xp67_ASAP7_75t_L g891 ( 
.A(n_755),
.B(n_734),
.Y(n_891)
);

O2A1O1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_778),
.A2(n_668),
.B(n_670),
.C(n_667),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_830),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_746),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_769),
.B(n_784),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_705),
.B(n_748),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_746),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_745),
.A2(n_633),
.B(n_632),
.Y(n_898)
);

BUFx4f_ASAP7_75t_L g899 ( 
.A(n_757),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_714),
.B(n_55),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_716),
.B(n_55),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_757),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_757),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_741),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_749),
.A2(n_675),
.B(n_686),
.C(n_683),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_749),
.B(n_56),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_742),
.A2(n_690),
.B(n_688),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_741),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_788),
.A2(n_691),
.B(n_690),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_760),
.B(n_57),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_751),
.B(n_57),
.Y(n_911)
);

AND2x6_ASAP7_75t_L g912 ( 
.A(n_816),
.B(n_693),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_751),
.B(n_58),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_841),
.A2(n_702),
.B1(n_695),
.B2(n_644),
.Y(n_914)
);

AO21x1_ASAP7_75t_L g915 ( 
.A1(n_844),
.A2(n_58),
.B(n_59),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_752),
.B(n_60),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_798),
.A2(n_721),
.B(n_719),
.C(n_811),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_815),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_814),
.B(n_798),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_743),
.B(n_60),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_768),
.A2(n_150),
.B(n_149),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_776),
.A2(n_154),
.B(n_153),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_780),
.B(n_61),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_733),
.A2(n_727),
.B1(n_806),
.B2(n_731),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_SL g925 ( 
.A(n_758),
.B(n_62),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_SL g926 ( 
.A1(n_758),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_825),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_812),
.B(n_67),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_790),
.B(n_68),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_835),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_821),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_794),
.A2(n_158),
.B(n_155),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_712),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_933)
);

BUFx8_ASAP7_75t_SL g934 ( 
.A(n_739),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_795),
.B(n_69),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_797),
.B(n_70),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_821),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_843),
.Y(n_938)
);

AND2x2_ASAP7_75t_SL g939 ( 
.A(n_841),
.B(n_72),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_821),
.B(n_777),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_810),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_801),
.A2(n_73),
.B1(n_76),
.B2(n_78),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_739),
.B(n_79),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_750),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_763),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_819),
.B(n_80),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_824),
.B(n_80),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_706),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_818),
.B(n_85),
.Y(n_949)
);

BUFx8_ASAP7_75t_L g950 ( 
.A(n_831),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_803),
.B(n_85),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_803),
.B(n_86),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_805),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_953)
);

NOR2x1p5_ASAP7_75t_SL g954 ( 
.A(n_848),
.B(n_177),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_817),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_754),
.B(n_87),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_SL g957 ( 
.A(n_771),
.B(n_89),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_SL g958 ( 
.A1(n_725),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_807),
.B(n_92),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_772),
.B(n_773),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_735),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_809),
.B(n_93),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_816),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_822),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_828),
.Y(n_965)
);

AO21x1_ASAP7_75t_L g966 ( 
.A1(n_844),
.A2(n_96),
.B(n_97),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_823),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_706),
.B(n_828),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_838),
.B(n_97),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_729),
.Y(n_970)
);

NOR2xp67_ASAP7_75t_L g971 ( 
.A(n_833),
.B(n_98),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_708),
.B(n_98),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_820),
.A2(n_211),
.B(n_268),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_766),
.B(n_99),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_708),
.B(n_100),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_710),
.B(n_102),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_710),
.B(n_102),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_792),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_715),
.B(n_104),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_829),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_816),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_804),
.B(n_809),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_770),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_839),
.B(n_106),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_845),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_756),
.B(n_110),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_759),
.B(n_111),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_826),
.B(n_112),
.Y(n_988)
);

AO21x1_ASAP7_75t_L g989 ( 
.A1(n_846),
.A2(n_847),
.B(n_850),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_761),
.A2(n_113),
.B(n_114),
.C(n_115),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_740),
.A2(n_214),
.B(n_260),
.Y(n_991)
);

AO21x1_ASAP7_75t_L g992 ( 
.A1(n_753),
.A2(n_115),
.B(n_116),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_762),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_767),
.A2(n_219),
.B(n_259),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_787),
.B(n_120),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_789),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_793),
.B(n_121),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_813),
.B(n_124),
.Y(n_998)
);

INVx4_ASAP7_75t_L g999 ( 
.A(n_836),
.Y(n_999)
);

NOR2xp67_ASAP7_75t_L g1000 ( 
.A(n_711),
.B(n_126),
.Y(n_1000)
);

BUFx4f_ASAP7_75t_L g1001 ( 
.A(n_802),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_934),
.Y(n_1002)
);

NAND2x1p5_ASAP7_75t_L g1003 ( 
.A(n_899),
.B(n_813),
.Y(n_1003)
);

INVx5_ASAP7_75t_L g1004 ( 
.A(n_902),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_862),
.B(n_127),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_917),
.A2(n_849),
.B(n_128),
.C(n_131),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_859),
.B(n_127),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_890),
.A2(n_870),
.B(n_862),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_960),
.A2(n_221),
.B(n_254),
.Y(n_1009)
);

AOI21xp33_ASAP7_75t_L g1010 ( 
.A1(n_982),
.A2(n_134),
.B(n_135),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_871),
.Y(n_1011)
);

NOR2x1_ASAP7_75t_L g1012 ( 
.A(n_879),
.B(n_134),
.Y(n_1012)
);

AOI21xp33_ASAP7_75t_L g1013 ( 
.A1(n_896),
.A2(n_940),
.B(n_968),
.Y(n_1013)
);

AND2x6_ASAP7_75t_L g1014 ( 
.A(n_984),
.B(n_138),
.Y(n_1014)
);

AO31x2_ASAP7_75t_L g1015 ( 
.A1(n_989),
.A2(n_138),
.A3(n_178),
.B(n_186),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_868),
.A2(n_187),
.B(n_188),
.Y(n_1016)
);

BUFx2_ASAP7_75t_R g1017 ( 
.A(n_955),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_852),
.B(n_189),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_855),
.B(n_190),
.Y(n_1019)
);

AO31x2_ASAP7_75t_L g1020 ( 
.A1(n_992),
.A2(n_191),
.A3(n_192),
.B(n_193),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_885),
.A2(n_194),
.B(n_226),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_891),
.B(n_229),
.Y(n_1022)
);

OA22x2_ASAP7_75t_L g1023 ( 
.A1(n_919),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_876),
.B(n_234),
.Y(n_1024)
);

AO21x2_ASAP7_75t_L g1025 ( 
.A1(n_921),
.A2(n_235),
.B(n_236),
.Y(n_1025)
);

NOR2x1_ASAP7_75t_SL g1026 ( 
.A(n_965),
.B(n_242),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_944),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_894),
.B(n_280),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_877),
.B(n_888),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_904),
.B(n_908),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_893),
.B(n_943),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_950),
.Y(n_1032)
);

CKINVDCx9p33_ASAP7_75t_R g1033 ( 
.A(n_928),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_907),
.A2(n_874),
.B(n_909),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_892),
.A2(n_967),
.B(n_898),
.Y(n_1035)
);

AOI211x1_ASAP7_75t_L g1036 ( 
.A1(n_915),
.A2(n_966),
.B(n_856),
.C(n_864),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_882),
.A2(n_889),
.B(n_887),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_875),
.B(n_970),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_SL g1039 ( 
.A1(n_922),
.A2(n_932),
.B(n_973),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_950),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_931),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_979),
.A2(n_995),
.B(n_987),
.C(n_974),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_863),
.A2(n_864),
.B(n_997),
.C(n_886),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_894),
.B(n_897),
.Y(n_1044)
);

AO31x2_ASAP7_75t_L g1045 ( 
.A1(n_854),
.A2(n_905),
.A3(n_923),
.B(n_929),
.Y(n_1045)
);

AOI221x1_ASAP7_75t_L g1046 ( 
.A1(n_973),
.A2(n_932),
.B1(n_922),
.B2(n_991),
.C(n_994),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_963),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_956),
.A2(n_986),
.B(n_878),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_939),
.B(n_918),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_910),
.B(n_858),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_963),
.Y(n_1051)
);

O2A1O1Ixp5_ASAP7_75t_L g1052 ( 
.A1(n_962),
.A2(n_976),
.B(n_977),
.C(n_972),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_929),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_935),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_936),
.A2(n_959),
.B(n_964),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_920),
.A2(n_906),
.B(n_913),
.C(n_911),
.Y(n_1056)
);

AND2x6_ASAP7_75t_SL g1057 ( 
.A(n_946),
.B(n_916),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_866),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_951),
.A2(n_952),
.B(n_975),
.C(n_988),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_866),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_897),
.B(n_903),
.Y(n_1061)
);

AOI21xp33_ASAP7_75t_L g1062 ( 
.A1(n_858),
.A2(n_860),
.B(n_978),
.Y(n_1062)
);

O2A1O1Ixp5_ASAP7_75t_L g1063 ( 
.A1(n_998),
.A2(n_949),
.B(n_873),
.C(n_883),
.Y(n_1063)
);

NAND2x1p5_ASAP7_75t_L g1064 ( 
.A(n_903),
.B(n_926),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_901),
.B(n_937),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_860),
.B(n_969),
.Y(n_1066)
);

INVx3_ASAP7_75t_SL g1067 ( 
.A(n_857),
.Y(n_1067)
);

AOI221xp5_ASAP7_75t_L g1068 ( 
.A1(n_861),
.A2(n_867),
.B1(n_925),
.B2(n_947),
.C(n_985),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_958),
.Y(n_1069)
);

INVx5_ASAP7_75t_L g1070 ( 
.A(n_912),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_980),
.B(n_916),
.Y(n_1071)
);

OR2x6_ASAP7_75t_L g1072 ( 
.A(n_865),
.B(n_953),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_999),
.B(n_961),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_969),
.B(n_924),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_945),
.Y(n_1075)
);

BUFx5_ASAP7_75t_L g1076 ( 
.A(n_912),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_941),
.B(n_999),
.Y(n_1077)
);

INVx5_ASAP7_75t_L g1078 ( 
.A(n_912),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_983),
.B(n_851),
.Y(n_1079)
);

AO31x2_ASAP7_75t_L g1080 ( 
.A1(n_914),
.A2(n_942),
.A3(n_953),
.B(n_985),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_SL g1081 ( 
.A(n_884),
.B(n_981),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_993),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_945),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_948),
.A2(n_927),
.B1(n_996),
.B2(n_933),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_1001),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_971),
.B(n_957),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1000),
.B(n_1001),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_912),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_954),
.A2(n_872),
.B(n_869),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_862),
.B(n_782),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_872),
.A2(n_869),
.B(n_832),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_862),
.B(n_782),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_872),
.A2(n_869),
.B(n_832),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_862),
.Y(n_1094)
);

INVxp67_ASAP7_75t_SL g1095 ( 
.A(n_859),
.Y(n_1095)
);

AOI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_982),
.A2(n_699),
.B(n_681),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_896),
.A2(n_939),
.B1(n_900),
.B2(n_925),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_862),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_881),
.B(n_764),
.Y(n_1099)
);

NOR2x1_ASAP7_75t_SL g1100 ( 
.A(n_859),
.B(n_862),
.Y(n_1100)
);

NAND2x1p5_ASAP7_75t_L g1101 ( 
.A(n_899),
.B(n_902),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_917),
.A2(n_982),
.B(n_979),
.C(n_885),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_934),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_872),
.A2(n_869),
.B(n_832),
.Y(n_1104)
);

NAND2x1_ASAP7_75t_L g1105 ( 
.A(n_912),
.B(n_938),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_SL g1106 ( 
.A1(n_921),
.A2(n_932),
.B(n_922),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_862),
.B(n_782),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_899),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_989),
.A2(n_872),
.A3(n_992),
.B(n_840),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_917),
.A2(n_982),
.B(n_979),
.C(n_885),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_859),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_862),
.B(n_782),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_934),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_862),
.B(n_782),
.Y(n_1114)
);

OAI21xp33_ASAP7_75t_SL g1115 ( 
.A1(n_939),
.A2(n_929),
.B(n_923),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_SL g1116 ( 
.A1(n_921),
.A2(n_932),
.B(n_922),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_881),
.B(n_764),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_862),
.B(n_782),
.Y(n_1118)
);

NAND2x1p5_ASAP7_75t_L g1119 ( 
.A(n_899),
.B(n_902),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_899),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_862),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_896),
.A2(n_939),
.B1(n_900),
.B2(n_925),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_862),
.B(n_782),
.Y(n_1123)
);

AO21x2_ASAP7_75t_L g1124 ( 
.A1(n_869),
.A2(n_872),
.B(n_921),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_862),
.B(n_782),
.Y(n_1125)
);

AOI21xp33_ASAP7_75t_L g1126 ( 
.A1(n_982),
.A2(n_699),
.B(n_681),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_939),
.A2(n_862),
.B1(n_895),
.B2(n_984),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_881),
.B(n_764),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_989),
.A2(n_872),
.A3(n_992),
.B(n_840),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_859),
.B(n_862),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_862),
.B(n_782),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_859),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_862),
.B(n_782),
.Y(n_1133)
);

AOI21xp33_ASAP7_75t_L g1134 ( 
.A1(n_982),
.A2(n_699),
.B(n_681),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_SL g1135 ( 
.A(n_925),
.B(n_588),
.C(n_576),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_862),
.B(n_782),
.Y(n_1136)
);

NAND2x1p5_ASAP7_75t_L g1137 ( 
.A(n_899),
.B(n_902),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_862),
.B(n_782),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_862),
.B(n_782),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_862),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_862),
.B(n_782),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_938),
.Y(n_1142)
);

INVxp67_ASAP7_75t_SL g1143 ( 
.A(n_859),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_862),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_SL g1145 ( 
.A(n_859),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_862),
.B(n_782),
.Y(n_1146)
);

NAND3xp33_ASAP7_75t_L g1147 ( 
.A(n_853),
.B(n_990),
.C(n_979),
.Y(n_1147)
);

AOI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_982),
.A2(n_699),
.B(n_681),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_930),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_859),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_938),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_862),
.Y(n_1152)
);

NAND3xp33_ASAP7_75t_L g1153 ( 
.A(n_853),
.B(n_990),
.C(n_979),
.Y(n_1153)
);

AO21x1_ASAP7_75t_L g1154 ( 
.A1(n_921),
.A2(n_932),
.B(n_922),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_859),
.Y(n_1155)
);

OAI22x1_ASAP7_75t_L g1156 ( 
.A1(n_859),
.A2(n_716),
.B1(n_734),
.B2(n_549),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_930),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_899),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_896),
.A2(n_939),
.B1(n_900),
.B2(n_925),
.Y(n_1159)
);

OR2x6_ASAP7_75t_L g1160 ( 
.A(n_859),
.B(n_746),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_862),
.B(n_782),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_862),
.B(n_782),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_939),
.A2(n_862),
.B1(n_895),
.B2(n_984),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_862),
.B(n_782),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_862),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_862),
.B(n_782),
.Y(n_1166)
);

O2A1O1Ixp5_ASAP7_75t_L g1167 ( 
.A1(n_880),
.A2(n_989),
.B(n_979),
.C(n_962),
.Y(n_1167)
);

NOR2x1_ASAP7_75t_R g1168 ( 
.A(n_1002),
.B(n_1113),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1094),
.B(n_1098),
.Y(n_1169)
);

NAND3xp33_ASAP7_75t_L g1170 ( 
.A(n_1036),
.B(n_1042),
.C(n_1043),
.Y(n_1170)
);

AO21x2_ASAP7_75t_L g1171 ( 
.A1(n_1106),
.A2(n_1116),
.B(n_1089),
.Y(n_1171)
);

NAND2x1p5_ASAP7_75t_L g1172 ( 
.A(n_1108),
.B(n_1070),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1111),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1130),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1039),
.A2(n_1059),
.B(n_1056),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1108),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_1105),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1004),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1013),
.B(n_1121),
.Y(n_1179)
);

OR2x6_ASAP7_75t_L g1180 ( 
.A(n_1160),
.B(n_1101),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1037),
.A2(n_1048),
.B(n_1154),
.Y(n_1181)
);

BUFx12f_ASAP7_75t_L g1182 ( 
.A(n_1032),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1034),
.A2(n_1046),
.B(n_1091),
.Y(n_1183)
);

OR2x6_ASAP7_75t_L g1184 ( 
.A(n_1160),
.B(n_1119),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_1090),
.B(n_1092),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1091),
.A2(n_1104),
.B(n_1093),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1127),
.A2(n_1163),
.B1(n_1122),
.B2(n_1159),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_1004),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1140),
.B(n_1144),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1147),
.A2(n_1153),
.B(n_1066),
.Y(n_1190)
);

AO21x1_ASAP7_75t_L g1191 ( 
.A1(n_1127),
.A2(n_1163),
.B(n_1021),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1152),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_1155),
.Y(n_1193)
);

NAND3xp33_ASAP7_75t_L g1194 ( 
.A(n_1036),
.B(n_1006),
.C(n_1068),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1097),
.A2(n_1122),
.B1(n_1159),
.B2(n_1165),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_SL g1196 ( 
.A1(n_1100),
.A2(n_1026),
.B(n_1055),
.Y(n_1196)
);

CKINVDCx16_ASAP7_75t_R g1197 ( 
.A(n_1103),
.Y(n_1197)
);

NAND2x1p5_ASAP7_75t_L g1198 ( 
.A(n_1070),
.B(n_1078),
.Y(n_1198)
);

INVx3_ASAP7_75t_SL g1199 ( 
.A(n_1160),
.Y(n_1199)
);

NOR2xp67_ASAP7_75t_L g1200 ( 
.A(n_1004),
.B(n_1040),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1107),
.B(n_1114),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1049),
.A2(n_1135),
.B1(n_1097),
.B2(n_1014),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1084),
.A2(n_1167),
.B(n_1052),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1112),
.B(n_1133),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_1118),
.B(n_1123),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1014),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_1030),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1014),
.A2(n_1053),
.B1(n_1054),
.B2(n_1072),
.Y(n_1208)
);

CKINVDCx11_ASAP7_75t_R g1209 ( 
.A(n_1067),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1115),
.B(n_1023),
.Y(n_1210)
);

AO21x2_ASAP7_75t_L g1211 ( 
.A1(n_1124),
.A2(n_1035),
.B(n_1055),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1070),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1050),
.A2(n_1166),
.B1(n_1125),
.B2(n_1131),
.Y(n_1213)
);

BUFx8_ASAP7_75t_L g1214 ( 
.A(n_1145),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1115),
.A2(n_1010),
.B(n_1074),
.C(n_1161),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1027),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_SL g1217 ( 
.A1(n_1008),
.A2(n_1016),
.B(n_1088),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1082),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1141),
.B(n_1164),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_1132),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_SL g1221 ( 
.A(n_1017),
.B(n_1137),
.Y(n_1221)
);

OA21x2_ASAP7_75t_L g1222 ( 
.A1(n_1016),
.A2(n_1063),
.B(n_1022),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1149),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1157),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1014),
.A2(n_1072),
.B1(n_1058),
.B2(n_1060),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1007),
.Y(n_1226)
);

BUFx2_ASAP7_75t_R g1227 ( 
.A(n_1069),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1072),
.A2(n_1065),
.B1(n_1007),
.B2(n_1062),
.Y(n_1228)
);

INVxp67_ASAP7_75t_SL g1229 ( 
.A(n_1047),
.Y(n_1229)
);

AOI22x1_ASAP7_75t_L g1230 ( 
.A1(n_1009),
.A2(n_1064),
.B1(n_1151),
.B2(n_1142),
.Y(n_1230)
);

AOI221xp5_ASAP7_75t_L g1231 ( 
.A1(n_1162),
.A2(n_1136),
.B1(n_1139),
.B2(n_1138),
.C(n_1146),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1029),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_SL g1233 ( 
.A1(n_1086),
.A2(n_1005),
.B(n_1077),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1150),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1038),
.Y(n_1235)
);

BUFx8_ASAP7_75t_L g1236 ( 
.A(n_1145),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1087),
.A2(n_1019),
.B(n_1018),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_1051),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1057),
.B(n_1096),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1011),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1031),
.B(n_1071),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1003),
.A2(n_1085),
.B(n_1073),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1071),
.Y(n_1243)
);

AOI22x1_ASAP7_75t_L g1244 ( 
.A1(n_1028),
.A2(n_1075),
.B1(n_1083),
.B2(n_1024),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1085),
.A2(n_1076),
.B(n_1012),
.Y(n_1245)
);

NAND3xp33_ASAP7_75t_L g1246 ( 
.A(n_1126),
.B(n_1148),
.C(n_1134),
.Y(n_1246)
);

AOI22x1_ASAP7_75t_L g1247 ( 
.A1(n_1028),
.A2(n_1083),
.B1(n_1075),
.B2(n_1156),
.Y(n_1247)
);

NOR2xp67_ASAP7_75t_L g1248 ( 
.A(n_1120),
.B(n_1158),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1109),
.A2(n_1129),
.A3(n_1015),
.B(n_1020),
.Y(n_1249)
);

AO21x2_ASAP7_75t_L g1250 ( 
.A1(n_1025),
.A2(n_1015),
.B(n_1109),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1099),
.B(n_1128),
.Y(n_1251)
);

OA21x2_ASAP7_75t_L g1252 ( 
.A1(n_1015),
.A2(n_1129),
.B(n_1109),
.Y(n_1252)
);

AO21x2_ASAP7_75t_L g1253 ( 
.A1(n_1025),
.A2(n_1045),
.B(n_1020),
.Y(n_1253)
);

INVx4_ASAP7_75t_SL g1254 ( 
.A(n_1080),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1044),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1081),
.A2(n_1143),
.B(n_1095),
.Y(n_1256)
);

NAND2x1p5_ASAP7_75t_L g1257 ( 
.A(n_1061),
.B(n_1041),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1080),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1079),
.B(n_1080),
.Y(n_1259)
);

INVx8_ASAP7_75t_L g1260 ( 
.A(n_1057),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1033),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1117),
.Y(n_1262)
);

AO21x2_ASAP7_75t_L g1263 ( 
.A1(n_1106),
.A2(n_1116),
.B(n_1089),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1112),
.B(n_1133),
.Y(n_1264)
);

NAND3xp33_ASAP7_75t_L g1265 ( 
.A(n_1036),
.B(n_1042),
.C(n_1043),
.Y(n_1265)
);

BUFx2_ASAP7_75t_SL g1266 ( 
.A(n_1103),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1108),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1043),
.A2(n_1110),
.B(n_1102),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1043),
.A2(n_1110),
.B(n_1102),
.Y(n_1269)
);

INVx3_ASAP7_75t_SL g1270 ( 
.A(n_1002),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1108),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1004),
.Y(n_1272)
);

AO21x2_ASAP7_75t_L g1273 ( 
.A1(n_1106),
.A2(n_1116),
.B(n_1089),
.Y(n_1273)
);

CKINVDCx8_ASAP7_75t_R g1274 ( 
.A(n_1032),
.Y(n_1274)
);

NAND3xp33_ASAP7_75t_L g1275 ( 
.A(n_1036),
.B(n_1042),
.C(n_1043),
.Y(n_1275)
);

AO21x2_ASAP7_75t_L g1276 ( 
.A1(n_1106),
.A2(n_1116),
.B(n_1089),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1013),
.B(n_724),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_1127),
.Y(n_1278)
);

BUFx4f_ASAP7_75t_SL g1279 ( 
.A(n_1103),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_SL g1280 ( 
.A1(n_1100),
.A2(n_1163),
.B(n_1127),
.Y(n_1280)
);

OAI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1246),
.A2(n_1213),
.B(n_1190),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1260),
.A2(n_1239),
.B1(n_1206),
.B2(n_1187),
.Y(n_1282)
);

BUFx10_ASAP7_75t_L g1283 ( 
.A(n_1180),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1218),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1216),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1229),
.Y(n_1286)
);

INVx4_ASAP7_75t_SL g1287 ( 
.A(n_1199),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1258),
.Y(n_1288)
);

NAND2x1p5_ASAP7_75t_L g1289 ( 
.A(n_1169),
.B(n_1189),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1259),
.Y(n_1290)
);

BUFx8_ASAP7_75t_L g1291 ( 
.A(n_1182),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1198),
.Y(n_1292)
);

BUFx12f_ASAP7_75t_L g1293 ( 
.A(n_1209),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1204),
.B(n_1232),
.Y(n_1294)
);

AO21x1_ASAP7_75t_SL g1295 ( 
.A1(n_1208),
.A2(n_1225),
.B(n_1202),
.Y(n_1295)
);

AOI21xp33_ASAP7_75t_L g1296 ( 
.A1(n_1215),
.A2(n_1233),
.B(n_1170),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1219),
.B(n_1264),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1185),
.B(n_1201),
.Y(n_1298)
);

CKINVDCx6p67_ASAP7_75t_R g1299 ( 
.A(n_1270),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1198),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1214),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1205),
.B(n_1231),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1208),
.B(n_1225),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1192),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1192),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1229),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1238),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1223),
.Y(n_1308)
);

BUFx2_ASAP7_75t_SL g1309 ( 
.A(n_1200),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1224),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1178),
.Y(n_1311)
);

OA21x2_ASAP7_75t_L g1312 ( 
.A1(n_1181),
.A2(n_1183),
.B(n_1175),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1235),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1169),
.B(n_1189),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_SL g1315 ( 
.A1(n_1260),
.A2(n_1239),
.B1(n_1280),
.B2(n_1195),
.Y(n_1315)
);

BUFx10_ASAP7_75t_L g1316 ( 
.A(n_1180),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1211),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_1180),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1211),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1231),
.B(n_1179),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1212),
.B(n_1177),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1188),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1179),
.B(n_1268),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1254),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1254),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1254),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1188),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1269),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1265),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1275),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1215),
.A2(n_1277),
.B(n_1203),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1210),
.Y(n_1332)
);

OR2x6_ASAP7_75t_L g1333 ( 
.A(n_1260),
.B(n_1184),
.Y(n_1333)
);

INVx1_ASAP7_75t_SL g1334 ( 
.A(n_1240),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_SL g1335 ( 
.A(n_1221),
.B(n_1227),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1172),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1222),
.A2(n_1217),
.B(n_1191),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1226),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1173),
.Y(n_1339)
);

AO21x2_ASAP7_75t_L g1340 ( 
.A1(n_1186),
.A2(n_1250),
.B(n_1253),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1241),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1277),
.A2(n_1228),
.B1(n_1202),
.B2(n_1262),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1288),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1288),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1328),
.B(n_1186),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1289),
.A2(n_1278),
.B1(n_1228),
.B2(n_1194),
.Y(n_1346)
);

INVx4_ASAP7_75t_L g1347 ( 
.A(n_1289),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1290),
.B(n_1171),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1324),
.B(n_1263),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_SL g1350 ( 
.A1(n_1309),
.A2(n_1266),
.B1(n_1197),
.B2(n_1261),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1286),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1306),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1323),
.B(n_1252),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1302),
.A2(n_1244),
.B1(n_1247),
.B2(n_1199),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1306),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1311),
.Y(n_1356)
);

BUFx2_ASAP7_75t_SL g1357 ( 
.A(n_1336),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1323),
.B(n_1273),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1340),
.B(n_1276),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1340),
.B(n_1276),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1314),
.A2(n_1196),
.B1(n_1262),
.B2(n_1230),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1307),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1320),
.B(n_1249),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1311),
.Y(n_1364)
);

INVx1_ASAP7_75t_SL g1365 ( 
.A(n_1322),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1312),
.B(n_1331),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1303),
.A2(n_1207),
.B1(n_1234),
.B2(n_1243),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1317),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1304),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1305),
.Y(n_1370)
);

INVx8_ASAP7_75t_L g1371 ( 
.A(n_1357),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1358),
.B(n_1325),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1358),
.B(n_1326),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1343),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1351),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1358),
.B(n_1326),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1366),
.B(n_1348),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1369),
.B(n_1313),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1343),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1344),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1352),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1366),
.B(n_1319),
.Y(n_1382)
);

NOR2xp67_ASAP7_75t_L g1383 ( 
.A(n_1354),
.B(n_1332),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1353),
.B(n_1329),
.Y(n_1384)
);

INVxp67_ASAP7_75t_SL g1385 ( 
.A(n_1351),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1366),
.B(n_1330),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1348),
.B(n_1330),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1348),
.B(n_1332),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1369),
.B(n_1285),
.Y(n_1389)
);

AND2x4_ASAP7_75t_SL g1390 ( 
.A(n_1347),
.B(n_1314),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1350),
.B(n_1274),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1370),
.B(n_1281),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1346),
.A2(n_1295),
.B1(n_1282),
.B2(n_1315),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1353),
.B(n_1294),
.Y(n_1394)
);

NOR2xp67_ASAP7_75t_L g1395 ( 
.A(n_1354),
.B(n_1337),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1368),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1370),
.B(n_1284),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1353),
.B(n_1298),
.Y(n_1398)
);

NOR2xp67_ASAP7_75t_L g1399 ( 
.A(n_1355),
.B(n_1336),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1355),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1362),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1350),
.B(n_1182),
.Y(n_1402)
);

AND2x4_ASAP7_75t_SL g1403 ( 
.A(n_1347),
.B(n_1314),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1391),
.B(n_1335),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1381),
.Y(n_1405)
);

NOR3x1_ASAP7_75t_L g1406 ( 
.A(n_1402),
.B(n_1318),
.C(n_1291),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1377),
.B(n_1359),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1374),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1396),
.Y(n_1409)
);

NOR3xp33_ASAP7_75t_SL g1410 ( 
.A(n_1392),
.B(n_1301),
.C(n_1346),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1389),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1374),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1377),
.B(n_1359),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1372),
.B(n_1349),
.Y(n_1414)
);

NOR3xp33_ASAP7_75t_L g1415 ( 
.A(n_1397),
.B(n_1296),
.C(n_1334),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1379),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1398),
.B(n_1345),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1398),
.B(n_1345),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1379),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1383),
.B(n_1365),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1378),
.Y(n_1421)
);

NOR2x1p5_ASAP7_75t_L g1422 ( 
.A(n_1385),
.B(n_1299),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1394),
.B(n_1363),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1394),
.B(n_1363),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1380),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1380),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1386),
.B(n_1359),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1386),
.B(n_1360),
.Y(n_1428)
);

NOR2xp67_ASAP7_75t_SL g1429 ( 
.A(n_1371),
.B(n_1309),
.Y(n_1429)
);

AND2x4_ASAP7_75t_SL g1430 ( 
.A(n_1375),
.B(n_1347),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1408),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1408),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1417),
.B(n_1384),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1407),
.B(n_1372),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1412),
.Y(n_1435)
);

OR2x6_ASAP7_75t_L g1436 ( 
.A(n_1422),
.B(n_1371),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1417),
.B(n_1384),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1412),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1414),
.B(n_1399),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1416),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1407),
.B(n_1373),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1416),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1413),
.B(n_1373),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1413),
.B(n_1376),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1419),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1419),
.Y(n_1446)
);

NAND5xp2_ASAP7_75t_SL g1447 ( 
.A(n_1415),
.B(n_1393),
.C(n_1301),
.D(n_1342),
.E(n_1367),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1427),
.B(n_1376),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1430),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1426),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1409),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1414),
.B(n_1399),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1418),
.B(n_1382),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1409),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1451),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1436),
.A2(n_1410),
.B1(n_1383),
.B2(n_1423),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1448),
.B(n_1427),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1434),
.B(n_1428),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1436),
.A2(n_1404),
.B(n_1395),
.Y(n_1459)
);

AOI211x1_ASAP7_75t_L g1460 ( 
.A1(n_1434),
.A2(n_1429),
.B(n_1421),
.C(n_1411),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1436),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1436),
.A2(n_1395),
.B(n_1420),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1453),
.B(n_1418),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1441),
.B(n_1428),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1441),
.B(n_1405),
.Y(n_1465)
);

AOI322xp5_ASAP7_75t_L g1466 ( 
.A1(n_1443),
.A2(n_1444),
.A3(n_1448),
.B1(n_1449),
.B2(n_1452),
.C1(n_1439),
.C2(n_1414),
.Y(n_1466)
);

OAI21xp33_ASAP7_75t_SL g1467 ( 
.A1(n_1443),
.A2(n_1424),
.B(n_1423),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1435),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1439),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1451),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1444),
.B(n_1424),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1433),
.Y(n_1472)
);

OAI21xp33_ASAP7_75t_SL g1473 ( 
.A1(n_1453),
.A2(n_1365),
.B(n_1400),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1435),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1433),
.B(n_1405),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1439),
.A2(n_1387),
.B1(n_1388),
.B2(n_1339),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1456),
.A2(n_1430),
.B(n_1452),
.Y(n_1477)
);

OAI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1467),
.A2(n_1473),
.B1(n_1466),
.B2(n_1461),
.C(n_1459),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1458),
.B(n_1437),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1463),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1461),
.A2(n_1447),
.B(n_1452),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1462),
.A2(n_1429),
.B(n_1361),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1476),
.A2(n_1472),
.B1(n_1465),
.B2(n_1469),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1475),
.A2(n_1447),
.B(n_1371),
.Y(n_1484)
);

INVx2_ASAP7_75t_SL g1485 ( 
.A(n_1475),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1463),
.Y(n_1486)
);

OAI21xp33_ASAP7_75t_L g1487 ( 
.A1(n_1469),
.A2(n_1437),
.B(n_1440),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1468),
.Y(n_1488)
);

A2O1A1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1478),
.A2(n_1469),
.B(n_1465),
.C(n_1458),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1480),
.B(n_1464),
.Y(n_1490)
);

AOI221x1_ASAP7_75t_L g1491 ( 
.A1(n_1481),
.A2(n_1474),
.B1(n_1468),
.B2(n_1471),
.C(n_1455),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1486),
.Y(n_1492)
);

OAI211xp5_ASAP7_75t_L g1493 ( 
.A1(n_1477),
.A2(n_1460),
.B(n_1209),
.C(n_1371),
.Y(n_1493)
);

AOI222xp33_ASAP7_75t_L g1494 ( 
.A1(n_1482),
.A2(n_1464),
.B1(n_1474),
.B2(n_1293),
.C1(n_1457),
.C2(n_1291),
.Y(n_1494)
);

OAI221xp5_ASAP7_75t_L g1495 ( 
.A1(n_1482),
.A2(n_1361),
.B1(n_1455),
.B2(n_1470),
.C(n_1432),
.Y(n_1495)
);

NOR3xp33_ASAP7_75t_L g1496 ( 
.A(n_1484),
.B(n_1168),
.C(n_1193),
.Y(n_1496)
);

AOI221xp5_ASAP7_75t_L g1497 ( 
.A1(n_1487),
.A2(n_1470),
.B1(n_1438),
.B2(n_1450),
.C(n_1446),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1485),
.A2(n_1483),
.B(n_1479),
.Y(n_1498)
);

NAND2x1p5_ASAP7_75t_L g1499 ( 
.A(n_1488),
.B(n_1356),
.Y(n_1499)
);

OAI211xp5_ASAP7_75t_L g1500 ( 
.A1(n_1477),
.A2(n_1371),
.B(n_1406),
.C(n_1291),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_SL g1501 ( 
.A1(n_1478),
.A2(n_1293),
.B1(n_1279),
.B2(n_1270),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1478),
.A2(n_1347),
.B1(n_1381),
.B2(n_1299),
.Y(n_1502)
);

AOI221xp5_ASAP7_75t_L g1503 ( 
.A1(n_1478),
.A2(n_1431),
.B1(n_1445),
.B2(n_1442),
.C(n_1440),
.Y(n_1503)
);

OAI211xp5_ASAP7_75t_L g1504 ( 
.A1(n_1489),
.A2(n_1227),
.B(n_1236),
.C(n_1214),
.Y(n_1504)
);

NOR3xp33_ASAP7_75t_L g1505 ( 
.A(n_1501),
.B(n_1220),
.C(n_1251),
.Y(n_1505)
);

NAND4xp25_ASAP7_75t_L g1506 ( 
.A(n_1494),
.B(n_1297),
.C(n_1248),
.D(n_1272),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1500),
.A2(n_1333),
.B(n_1184),
.Y(n_1507)
);

NOR3xp33_ASAP7_75t_SL g1508 ( 
.A(n_1502),
.B(n_1279),
.C(n_1236),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1493),
.B(n_1442),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_SL g1510 ( 
.A1(n_1503),
.A2(n_1403),
.B(n_1390),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1492),
.B(n_1425),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1498),
.B(n_1490),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1499),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1497),
.B(n_1401),
.Y(n_1514)
);

OAI211xp5_ASAP7_75t_SL g1515 ( 
.A1(n_1495),
.A2(n_1318),
.B(n_1341),
.C(n_1267),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1512),
.B(n_1491),
.Y(n_1516)
);

NOR2xp67_ASAP7_75t_L g1517 ( 
.A(n_1504),
.B(n_1496),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1509),
.B(n_1499),
.Y(n_1518)
);

NOR4xp75_ASAP7_75t_L g1519 ( 
.A(n_1514),
.B(n_1176),
.C(n_1271),
.D(n_1267),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1511),
.B(n_1454),
.Y(n_1520)
);

OAI211xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1510),
.A2(n_1271),
.B(n_1176),
.C(n_1336),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1505),
.Y(n_1522)
);

NAND4xp25_ASAP7_75t_L g1523 ( 
.A(n_1507),
.B(n_1272),
.C(n_1364),
.D(n_1356),
.Y(n_1523)
);

AO22x2_ASAP7_75t_L g1524 ( 
.A1(n_1513),
.A2(n_1287),
.B1(n_1357),
.B2(n_1338),
.Y(n_1524)
);

NOR2xp67_ASAP7_75t_L g1525 ( 
.A(n_1506),
.B(n_1454),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1508),
.B(n_1387),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1517),
.B(n_1515),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1526),
.Y(n_1528)
);

AO22x2_ASAP7_75t_L g1529 ( 
.A1(n_1522),
.A2(n_1287),
.B1(n_1310),
.B2(n_1308),
.Y(n_1529)
);

NOR3x1_ASAP7_75t_L g1530 ( 
.A(n_1516),
.B(n_1245),
.C(n_1333),
.Y(n_1530)
);

NOR3xp33_ASAP7_75t_SL g1531 ( 
.A(n_1521),
.B(n_1523),
.C(n_1518),
.Y(n_1531)
);

NOR3xp33_ASAP7_75t_L g1532 ( 
.A(n_1525),
.B(n_1212),
.C(n_1242),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1520),
.B(n_1426),
.Y(n_1533)
);

NOR2x1_ASAP7_75t_L g1534 ( 
.A(n_1519),
.B(n_1184),
.Y(n_1534)
);

NAND3xp33_ASAP7_75t_SL g1535 ( 
.A(n_1524),
.B(n_1172),
.C(n_1257),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1524),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1526),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1517),
.A2(n_1237),
.B(n_1256),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1528),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1537),
.B(n_1363),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1527),
.A2(n_1333),
.B1(n_1287),
.B2(n_1316),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1529),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1531),
.A2(n_1333),
.B1(n_1287),
.B2(n_1316),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1530),
.B(n_1388),
.Y(n_1544)
);

XNOR2xp5_ASAP7_75t_L g1545 ( 
.A(n_1543),
.B(n_1534),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1542),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1539),
.A2(n_1536),
.B1(n_1529),
.B2(n_1533),
.Y(n_1547)
);

NOR2x1_ASAP7_75t_L g1548 ( 
.A(n_1540),
.B(n_1535),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1544),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1546),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1548),
.Y(n_1551)
);

XNOR2x2_ASAP7_75t_L g1552 ( 
.A(n_1551),
.B(n_1547),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1550),
.A2(n_1545),
.B(n_1549),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1552),
.Y(n_1554)
);

AOI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1553),
.A2(n_1541),
.B1(n_1532),
.B2(n_1538),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1554),
.A2(n_1257),
.B(n_1322),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1555),
.A2(n_1283),
.B1(n_1316),
.B2(n_1327),
.Y(n_1557)
);

AO221x1_ASAP7_75t_L g1558 ( 
.A1(n_1557),
.A2(n_1292),
.B1(n_1300),
.B2(n_1255),
.C(n_1174),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1558),
.A2(n_1556),
.B(n_1327),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1559),
.B(n_1356),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1560),
.A2(n_1364),
.B1(n_1283),
.B2(n_1321),
.Y(n_1561)
);


endmodule