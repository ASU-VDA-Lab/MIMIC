module fake_jpeg_7547_n_258 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_17),
.Y(n_50)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_16),
.B1(n_28),
.B2(n_23),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_43),
.A2(n_48),
.B1(n_49),
.B2(n_57),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_56),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_34),
.A2(n_16),
.B1(n_28),
.B2(n_23),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_30),
.B1(n_21),
.B2(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_50),
.B(n_65),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_24),
.B1(n_15),
.B2(n_27),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_63),
.B1(n_37),
.B2(n_19),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_0),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_60),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_35),
.A2(n_30),
.B1(n_18),
.B2(n_21),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_33),
.B(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_29),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_35),
.A2(n_27),
.B1(n_26),
.B2(n_15),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_26),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_73),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx2_ASAP7_75t_SL g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_64),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_60),
.B(n_38),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_78),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_81),
.B1(n_64),
.B2(n_46),
.Y(n_91)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_62),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_38),
.B1(n_29),
.B2(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_54),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_25),
.B1(n_22),
.B2(n_8),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_85),
.B1(n_65),
.B2(n_58),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_25),
.B1(n_22),
.B2(n_8),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_74),
.B1(n_72),
.B2(n_69),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_102),
.B1(n_81),
.B2(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_94),
.B(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_53),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_62),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_99),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_82),
.C(n_73),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_106),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_71),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_105),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_45),
.B1(n_58),
.B2(n_53),
.Y(n_102)
);

AO21x1_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_66),
.B(n_86),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_54),
.B(n_52),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_56),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_83),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_109),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_58),
.B1(n_45),
.B2(n_47),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_80),
.B1(n_78),
.B2(n_61),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_120),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_111),
.A2(n_91),
.B1(n_89),
.B2(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_112),
.B(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_122),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_84),
.B1(n_45),
.B2(n_69),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_115),
.B1(n_92),
.B2(n_102),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_119),
.B(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_66),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

INVxp67_ASAP7_75t_SL g122 ( 
.A(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_106),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_99),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_98),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_107),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_74),
.B1(n_80),
.B2(n_25),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_129),
.A2(n_87),
.B(n_101),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_68),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_131),
.B(n_132),
.Y(n_152)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_146),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_136),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_149),
.B1(n_154),
.B2(n_155),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_141),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_89),
.Y(n_140)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_117),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_123),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_150),
.Y(n_169)
);

BUFx24_ASAP7_75t_SL g143 ( 
.A(n_124),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_106),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_110),
.C(n_120),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_108),
.B1(n_94),
.B2(n_97),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_111),
.A2(n_87),
.B1(n_107),
.B2(n_95),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_166),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_168),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_167),
.C(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_130),
.C(n_119),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_133),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_130),
.C(n_119),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_172),
.B(n_130),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_174),
.Y(n_193)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_128),
.B1(n_115),
.B2(n_114),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_175),
.A2(n_147),
.B1(n_135),
.B2(n_128),
.Y(n_181)
);

BUFx12f_ASAP7_75t_SL g176 ( 
.A(n_134),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_124),
.B(n_132),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_178),
.B(n_192),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_146),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_194),
.Y(n_200)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_190),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_176),
.A2(n_149),
.B1(n_155),
.B2(n_154),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_183),
.A2(n_185),
.B1(n_191),
.B2(n_177),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_171),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_188),
.C(n_189),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_153),
.B1(n_138),
.B2(n_114),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_129),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_142),
.C(n_121),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_114),
.B1(n_141),
.B2(n_136),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_140),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_172),
.C(n_170),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_196),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_113),
.C(n_126),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_169),
.C(n_175),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_186),
.B1(n_22),
.B2(n_9),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_195),
.A2(n_160),
.B1(n_158),
.B2(n_114),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_212),
.B1(n_59),
.B2(n_1),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_157),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_22),
.C(n_68),
.Y(n_220)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_180),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_207),
.Y(n_213)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_159),
.Y(n_210)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_113),
.Y(n_211)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_189),
.A2(n_127),
.B1(n_55),
.B2(n_44),
.Y(n_212)
);

AO22x2_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_188),
.B1(n_179),
.B2(n_186),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_214),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_202),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_68),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_218),
.B(n_224),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_221),
.C(n_225),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_59),
.C(n_22),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_199),
.B1(n_201),
.B2(n_10),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_6),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_8),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_219),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_229),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_203),
.B1(n_202),
.B2(n_198),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_5),
.B1(n_12),
.B2(n_11),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_225),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_200),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_220),
.B(n_214),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_201),
.C(n_200),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_227),
.C(n_232),
.Y(n_242)
);

NOR4xp25_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_5),
.C(n_12),
.D(n_11),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_10),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_232),
.A2(n_213),
.B1(n_214),
.B2(n_216),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_239),
.B1(n_0),
.B2(n_1),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_240),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_215),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_241),
.B(n_4),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_233),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_4),
.Y(n_248)
);

AOI322xp5_ASAP7_75t_L g250 ( 
.A1(n_244),
.A2(n_247),
.A3(n_237),
.B1(n_236),
.B2(n_238),
.C1(n_9),
.C2(n_14),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_245),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_4),
.C(n_12),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_248),
.C(n_0),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_252),
.C(n_253),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_249),
.A2(n_14),
.B1(n_1),
.B2(n_2),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_245),
.C(n_2),
.Y(n_255)
);

AOI21x1_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_3),
.B(n_254),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_3),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_3),
.Y(n_258)
);


endmodule