module real_jpeg_18019_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_579),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_0),
.B(n_580),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_1),
.A2(n_27),
.B1(n_32),
.B2(n_35),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_1),
.A2(n_35),
.B1(n_222),
.B2(n_226),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_1),
.A2(n_35),
.B1(n_279),
.B2(n_284),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_1),
.A2(n_35),
.B1(n_356),
.B2(n_361),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_2),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_2),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_3),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_3),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_3),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_3),
.Y(n_129)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_3),
.Y(n_414)
);

BUFx5_ASAP7_75t_L g419 ( 
.A(n_3),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_4),
.A2(n_182),
.B1(n_185),
.B2(n_187),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_4),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_4),
.A2(n_187),
.B1(n_243),
.B2(n_246),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_4),
.A2(n_133),
.B1(n_187),
.B2(n_443),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_4),
.A2(n_187),
.B1(n_452),
.B2(n_456),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_5),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_54)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_5),
.A2(n_60),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_5),
.A2(n_60),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_5),
.A2(n_60),
.B1(n_303),
.B2(n_305),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_6),
.A2(n_27),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_6),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_6),
.A2(n_178),
.B1(n_328),
.B2(n_330),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_6),
.A2(n_178),
.B1(n_430),
.B2(n_431),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_6),
.A2(n_178),
.B1(n_471),
.B2(n_474),
.Y(n_470)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_7),
.A2(n_57),
.A3(n_199),
.B1(n_203),
.B2(n_207),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_7),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_7),
.A2(n_206),
.B1(n_251),
.B2(n_253),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_7),
.B(n_45),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_7),
.B(n_92),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_7),
.B(n_346),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_7),
.B(n_111),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_SL g500 ( 
.A1(n_7),
.A2(n_206),
.B1(n_243),
.B2(n_501),
.Y(n_500)
);

OAI32xp33_ASAP7_75t_L g505 ( 
.A1(n_7),
.A2(n_506),
.A3(n_509),
.B1(n_513),
.B2(n_518),
.Y(n_505)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_8),
.Y(n_220)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_8),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_8),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g347 ( 
.A(n_8),
.Y(n_347)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_9),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_10),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_10),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_10),
.Y(n_122)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_10),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_10),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_10),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_10),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_10),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_11),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_11),
.A2(n_33),
.B1(n_72),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_11),
.A2(n_72),
.B1(n_259),
.B2(n_261),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_11),
.A2(n_72),
.B1(n_271),
.B2(n_275),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_12),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_190)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_12),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_12),
.A2(n_194),
.B1(n_254),
.B2(n_315),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_12),
.A2(n_194),
.B1(n_436),
.B2(n_437),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_SL g495 ( 
.A1(n_12),
.A2(n_194),
.B1(n_496),
.B2(n_498),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_13),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_13),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_13),
.A2(n_105),
.B1(n_133),
.B2(n_138),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_13),
.A2(n_105),
.B1(n_296),
.B2(n_298),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_13),
.A2(n_105),
.B1(n_368),
.B2(n_370),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_14),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_16),
.Y(n_113)
);

BUFx4f_ASAP7_75t_L g117 ( 
.A(n_16),
.Y(n_117)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_16),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_16),
.Y(n_410)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g184 ( 
.A(n_17),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_165),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_163),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_156),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_22),
.B(n_156),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_143),
.C(n_148),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_24),
.A2(n_143),
.B1(n_558),
.B2(n_559),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_24),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_65),
.Y(n_24)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_25),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_36),
.B1(n_54),
.B2(n_64),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_26),
.A2(n_64),
.B(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_38),
.B1(n_40),
.B2(n_42),
.Y(n_37)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_29),
.Y(n_254)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_30),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_33),
.Y(n_146)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_36),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_36),
.A2(n_54),
.B(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_36),
.A2(n_64),
.B1(n_177),
.B2(n_250),
.Y(n_249)
);

OAI22x1_ASAP7_75t_SL g313 ( 
.A1(n_36),
.A2(n_64),
.B1(n_181),
.B2(n_314),
.Y(n_313)
);

OAI21x1_ASAP7_75t_SL g365 ( 
.A1(n_36),
.A2(n_314),
.B(n_366),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_36),
.A2(n_158),
.B(n_392),
.Y(n_391)
);

OR2x6_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_45),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_41),
.Y(n_210)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_45),
.B(n_145),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_45),
.A2(n_147),
.B1(n_176),
.B2(n_180),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_45),
.B(n_367),
.Y(n_366)
);

AO22x2_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_47),
.Y(n_196)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_47),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_48),
.Y(n_360)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_51),
.Y(n_329)
);

INVx6_ASAP7_75t_L g520 ( 
.A(n_51),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_62),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_63),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g252 ( 
.A(n_63),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_110),
.B2(n_142),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_66),
.B(n_142),
.C(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AO21x1_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_76),
.B(n_99),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_69),
.B(n_92),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_69),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_75),
.Y(n_193)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_75),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_76),
.A2(n_150),
.B(n_154),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_76),
.A2(n_92),
.B(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_76),
.A2(n_99),
.B(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_76),
.A2(n_92),
.B1(n_150),
.B2(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_77),
.A2(n_100),
.B1(n_190),
.B2(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_77),
.A2(n_101),
.B(n_155),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_77),
.A2(n_100),
.B1(n_242),
.B2(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_77),
.A2(n_100),
.B1(n_354),
.B2(n_355),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_77),
.A2(n_100),
.B1(n_327),
.B2(n_500),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_92),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_83),
.B1(n_86),
.B2(n_91),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_84),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_89),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

AO22x2_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_95),
.Y(n_430)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_96),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_96),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_96),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_97),
.Y(n_405)
);

NOR2xp67_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

INVxp33_ASAP7_75t_SL g160 ( 
.A(n_101),
.Y(n_160)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_102),
.Y(n_503)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_104),
.Y(n_205)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_104),
.Y(n_245)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_143),
.C(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_110),
.B(n_149),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_119),
.B(n_131),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_111),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_111),
.B(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_111),
.A2(n_119),
.B1(n_425),
.B2(n_429),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_111),
.A2(n_119),
.B1(n_429),
.B2(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_112),
.A2(n_256),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_112),
.B(n_132),
.Y(n_386)
);

OAI22xp33_ASAP7_75t_L g493 ( 
.A1(n_112),
.A2(n_256),
.B1(n_494),
.B2(n_495),
.Y(n_493)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_118),
.Y(n_112)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_113),
.Y(n_218)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_113),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_113),
.Y(n_436)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_113),
.Y(n_473)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_113),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_116),
.Y(n_480)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_117),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_117),
.Y(n_297)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_117),
.Y(n_455)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_119),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_119),
.B(n_258),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_119),
.A2(n_386),
.B(n_535),
.Y(n_534)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_123),
.B1(n_126),
.B2(n_130),
.Y(n_120)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_132),
.A2(n_256),
.B(n_257),
.Y(n_255)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_137),
.Y(n_263)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_137),
.Y(n_512)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_143),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_143),
.A2(n_559),
.B1(n_563),
.B2(n_564),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_148),
.B(n_557),
.Y(n_556)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_SL g330 ( 
.A(n_153),
.Y(n_330)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g582 ( 
.A(n_156),
.Y(n_582)
);

FAx1_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_159),
.CI(n_161),
.CON(n_156),
.SN(n_156)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_554),
.B(n_576),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_548),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_397),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_337),
.C(n_375),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_319),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_287),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_172),
.B(n_287),
.C(n_550),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_240),
.C(n_264),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_173),
.B(n_336),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_197),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_188),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_175),
.B(n_188),
.C(n_197),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_184),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_184),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_214),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_198),
.B(n_214),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_206),
.B(n_416),
.Y(n_415)
);

OAI21xp33_ASAP7_75t_SL g425 ( 
.A1(n_206),
.A2(n_415),
.B(n_426),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_206),
.A2(n_216),
.B1(n_467),
.B2(n_470),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_206),
.B(n_514),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_221),
.B1(n_228),
.B2(n_233),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_215),
.A2(n_233),
.B(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_215),
.A2(n_450),
.B1(n_460),
.B2(n_461),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_215),
.A2(n_266),
.B(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_216),
.B(n_270),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_216),
.A2(n_295),
.B(n_344),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_216),
.A2(n_435),
.B(n_439),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_216),
.A2(n_451),
.B1(n_470),
.B2(n_483),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_219),
.A2(n_221),
.B(n_299),
.Y(n_334)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_224),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_226),
.Y(n_298)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_230),
.Y(n_294)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_230),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_232),
.Y(n_469)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_240),
.B(n_264),
.Y(n_336)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_249),
.C(n_255),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_241),
.B(n_255),
.Y(n_322)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_249),
.B(n_322),
.Y(n_321)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OA21x2_ASAP7_75t_L g349 ( 
.A1(n_256),
.A2(n_257),
.B(n_302),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_259),
.Y(n_498)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_262),
.Y(n_497)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_276),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_265),
.B(n_276),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_286),
.Y(n_276)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_278),
.Y(n_301)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_282),
.Y(n_304)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_282),
.Y(n_432)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_282),
.Y(n_445)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_283),
.Y(n_428)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVxp33_ASAP7_75t_L g387 ( 
.A(n_286),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_288),
.B(n_309),
.C(n_318),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_309),
.B1(n_310),
.B2(n_318),
.Y(n_289)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_290),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_300),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_291),
.B(n_300),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_299),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_292),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_295),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_311),
.B(n_313),
.C(n_317),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_317),
.Y(n_312)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_335),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_320),
.B(n_335),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.C(n_325),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_321),
.B(n_545),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_323),
.A2(n_324),
.B1(n_325),
.B2(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_325),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_331),
.C(n_333),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_326),
.B(n_538),
.Y(n_537)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_331),
.A2(n_332),
.B1(n_334),
.B2(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_334),
.Y(n_539)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g548 ( 
.A1(n_338),
.A2(n_549),
.B(n_551),
.C(n_552),
.D(n_553),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_339),
.B(n_340),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_340)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_341),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_351),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_342),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_343),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_342)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_343),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_343),
.A2(n_350),
.B1(n_391),
.B2(n_393),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_343),
.B(n_349),
.Y(n_394)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_344),
.Y(n_461)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx12f_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

AOI21xp33_ASAP7_75t_L g567 ( 
.A1(n_350),
.A2(n_393),
.B(n_568),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_372),
.C(n_377),
.Y(n_376)
);

XNOR2x1_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_371),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_365),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_355),
.Y(n_384)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_360),
.Y(n_364)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_365),
.B(n_371),
.C(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_367),
.Y(n_392)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_375),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_378),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_376),
.B(n_378),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_381),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_379),
.B(n_395),
.C(n_571),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_389),
.B1(n_395),
.B2(n_396),
.Y(n_381)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_382),
.Y(n_395)
);

OAI21xp33_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_385),
.B(n_388),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_383),
.B(n_385),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_388),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_388),
.A2(n_562),
.B1(n_565),
.B2(n_575),
.Y(n_574)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_389),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_389),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_394),
.Y(n_389)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_391),
.Y(n_393)
);

INVxp33_ASAP7_75t_L g568 ( 
.A(n_394),
.Y(n_568)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_542),
.B(n_547),
.Y(n_397)
);

AOI21x1_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_527),
.B(n_541),
.Y(n_398)
);

OAI21x1_ASAP7_75t_SL g399 ( 
.A1(n_400),
.A2(n_489),
.B(n_526),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_447),
.B(n_488),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_433),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_402),
.B(n_433),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_423),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_403),
.A2(n_423),
.B1(n_424),
.B2(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_403),
.Y(n_463)
);

OAI32xp33_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_406),
.A3(n_411),
.B1(n_415),
.B2(n_417),
.Y(n_403)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_409),
.Y(n_459)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_410),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx5_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_440),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_434),
.B(n_441),
.C(n_446),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_435),
.Y(n_460)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_446),
.Y(n_440)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_442),
.Y(n_494)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_448),
.A2(n_464),
.B(n_487),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_462),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_SL g487 ( 
.A(n_449),
.B(n_462),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_465),
.A2(n_481),
.B(n_486),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_477),
.Y(n_465)
);

INVx6_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx6_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_482),
.B(n_485),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_482),
.B(n_485),
.Y(n_486)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_490),
.B(n_491),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_504),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_499),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_493),
.Y(n_529)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_495),
.Y(n_535)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_499),
.Y(n_530)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_504),
.B(n_529),
.C(n_530),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_524),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_505),
.B(n_524),
.Y(n_533)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_521),
.Y(n_518)
);

INVx6_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_531),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_528),
.B(n_531),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_532),
.A2(n_536),
.B1(n_537),
.B2(n_540),
.Y(n_531)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_532),
.Y(n_540)
);

XOR2x1_ASAP7_75t_SL g532 ( 
.A(n_533),
.B(n_534),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_533),
.B(n_534),
.C(n_536),
.Y(n_543)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_543),
.B(n_544),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_543),
.B(n_544),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_555),
.B(n_569),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_555),
.A2(n_577),
.B(n_578),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_560),
.Y(n_555)
);

NAND2xp33_ASAP7_75t_SL g578 ( 
.A(n_556),
.B(n_560),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_565),
.C(n_566),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_562),
.Y(n_575)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_563),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_566),
.A2(n_567),
.B1(n_573),
.B2(n_574),
.Y(n_572)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_570),
.B(n_572),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_570),
.B(n_572),
.Y(n_577)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);


endmodule