module fake_jpeg_25814_n_23 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_23);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_23;

wire n_13;
wire n_21;
wire n_10;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_9),
.A2(n_6),
.B1(n_2),
.B2(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_13),
.B(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_15),
.Y(n_17)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_11),
.B1(n_10),
.B2(n_3),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_19),
.B1(n_15),
.B2(n_12),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_16),
.A2(n_12),
.B1(n_10),
.B2(n_5),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_21),
.C(n_1),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_22),
.A2(n_1),
.B1(n_3),
.B2(n_7),
.Y(n_23)
);


endmodule