module fake_jpeg_26280_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_7),
.B(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_39),
.Y(n_51)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_21),
.B1(n_27),
.B2(n_18),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_47),
.A2(n_35),
.B1(n_23),
.B2(n_26),
.Y(n_98)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_21),
.B1(n_27),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_35),
.B1(n_18),
.B2(n_21),
.Y(n_69)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_52),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_24),
.Y(n_55)
);

OR2x2_ASAP7_75t_SL g81 ( 
.A(n_55),
.B(n_54),
.Y(n_81)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_60),
.Y(n_86)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_75),
.Y(n_114)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_67),
.B(n_71),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_69),
.A2(n_82),
.B1(n_24),
.B2(n_16),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_25),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_70),
.B(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_73),
.B(n_84),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_74),
.Y(n_112)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_80),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_25),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_81),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_51),
.B1(n_27),
.B2(n_37),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_79),
.A2(n_83),
.B1(n_98),
.B2(n_23),
.Y(n_107)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_30),
.B1(n_29),
.B2(n_17),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_17),
.B1(n_30),
.B2(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_40),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_40),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_41),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_88),
.Y(n_134)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_51),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_91),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_33),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_93),
.Y(n_132)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_25),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_100),
.C(n_22),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_56),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_96),
.Y(n_133)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_33),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_25),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_31),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_54),
.B(n_17),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_111),
.B1(n_78),
.B2(n_104),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_26),
.B1(n_23),
.B2(n_30),
.Y(n_111)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_125),
.B1(n_92),
.B2(n_86),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_83),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_78),
.A2(n_17),
.B1(n_30),
.B2(n_29),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_129),
.Y(n_141)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

AOI32xp33_ASAP7_75t_L g130 ( 
.A1(n_81),
.A2(n_22),
.A3(n_35),
.B1(n_29),
.B2(n_16),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_130),
.A2(n_110),
.B(n_127),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_135),
.B(n_136),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_122),
.B(n_19),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_129),
.B1(n_120),
.B2(n_131),
.Y(n_179)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_138),
.B(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_70),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_147),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_110),
.A2(n_70),
.B1(n_103),
.B2(n_88),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_142),
.A2(n_144),
.B1(n_154),
.B2(n_115),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_143),
.A2(n_148),
.B(n_152),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_128),
.A2(n_72),
.B1(n_75),
.B2(n_80),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_156),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_104),
.B(n_86),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_153),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_107),
.A2(n_100),
.B1(n_95),
.B2(n_94),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_151),
.A2(n_155),
.B1(n_106),
.B2(n_97),
.Y(n_169)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_111),
.A2(n_100),
.B1(n_95),
.B2(n_92),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_117),
.B(n_64),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_161),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_89),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_160),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_113),
.B(n_19),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_118),
.B(n_64),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_105),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_132),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_90),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_152),
.A2(n_109),
.B(n_124),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_106),
.B(n_109),
.Y(n_168)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_178),
.B1(n_179),
.B2(n_186),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_108),
.B(n_131),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_177),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_68),
.Y(n_172)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_116),
.B(n_118),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_139),
.Y(n_205)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_181),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_145),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_137),
.A2(n_151),
.B1(n_155),
.B2(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_182),
.Y(n_226)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_184),
.Y(n_216)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_135),
.A2(n_115),
.B1(n_108),
.B2(n_116),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_189),
.Y(n_221)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_147),
.A2(n_26),
.B1(n_34),
.B2(n_2),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_191),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_34),
.Y(n_193)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_138),
.B(n_7),
.C(n_14),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_9),
.C(n_14),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_160),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_201),
.B(n_205),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_209),
.Y(n_244)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_165),
.B(n_162),
.CI(n_9),
.CON(n_209),
.SN(n_209)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_212),
.Y(n_237)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_8),
.C(n_15),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_157),
.C(n_8),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_224),
.C(n_225),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_168),
.A2(n_157),
.B1(n_9),
.B2(n_2),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_169),
.B1(n_186),
.B2(n_172),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_197),
.B1(n_191),
.B2(n_188),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_217),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_194),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_219),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_166),
.B(n_10),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_196),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_180),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_223),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_187),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_178),
.B(n_10),
.C(n_3),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_165),
.B(n_11),
.C(n_4),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_167),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_173),
.Y(n_228)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_229),
.A2(n_238),
.B1(n_242),
.B2(n_221),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_218),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_243),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_168),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_200),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_233),
.B(n_250),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_176),
.Y(n_235)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_170),
.C(n_174),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_236),
.B(n_249),
.C(n_208),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_201),
.B(n_172),
.CI(n_175),
.CON(n_241),
.SN(n_241)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_251),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_202),
.A2(n_183),
.B1(n_171),
.B2(n_181),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

AND2x2_ASAP7_75t_SL g245 ( 
.A(n_200),
.B(n_189),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_204),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_202),
.B(n_185),
.C(n_4),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_220),
.B(n_5),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_207),
.A2(n_0),
.B(n_6),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_253),
.B(n_266),
.Y(n_281)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_257),
.B(n_259),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_213),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_258),
.B(n_265),
.Y(n_288)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_228),
.B(n_199),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_262),
.B(n_264),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_211),
.B1(n_207),
.B2(n_203),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_263),
.A2(n_270),
.B1(n_249),
.B2(n_254),
.Y(n_274)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_230),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_224),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_209),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_267),
.B(n_268),
.Y(n_286)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_211),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_269),
.B(n_271),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_277),
.B1(n_241),
.B2(n_210),
.Y(n_290)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_276),
.Y(n_296)
);

INVx13_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_261),
.A2(n_245),
.B1(n_247),
.B2(n_240),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_206),
.Y(n_278)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_282),
.Y(n_299)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

A2O1A1O1Ixp25_ASAP7_75t_L g283 ( 
.A1(n_252),
.A2(n_241),
.B(n_269),
.C(n_265),
.D(n_258),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_250),
.Y(n_292)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_284),
.B(n_231),
.Y(n_295)
);

OAI211xp5_ASAP7_75t_L g285 ( 
.A1(n_252),
.A2(n_244),
.B(n_237),
.C(n_209),
.Y(n_285)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_225),
.Y(n_291)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_291),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_292),
.B(n_283),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_231),
.C(n_226),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_293),
.B(n_300),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_272),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_14),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_295),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_286),
.A2(n_251),
.B(n_226),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_302),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_234),
.C(n_215),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_6),
.C(n_12),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_301),
.B(n_274),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_278),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_305),
.Y(n_314)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_291),
.A2(n_273),
.B1(n_276),
.B2(n_280),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_312),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_299),
.B(n_297),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_301),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_315),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_293),
.C(n_300),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_318),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_319),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_289),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_15),
.Y(n_319)
);

NOR3xp33_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_307),
.C(n_312),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_306),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_313),
.B(n_309),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_324),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_326),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_327),
.A2(n_323),
.B(n_321),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_325),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_281),
.Y(n_330)
);


endmodule