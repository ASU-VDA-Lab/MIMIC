module real_aes_9177_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_725;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_359;
wire n_156;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g178 ( .A1(n_0), .A2(n_179), .B(n_182), .C(n_186), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_1), .B(n_170), .Y(n_189) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_3), .B(n_180), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_4), .A2(n_139), .B(n_501), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_5), .A2(n_144), .B(n_147), .C(n_528), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_6), .A2(n_139), .B(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_7), .B(n_170), .Y(n_507) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_8), .A2(n_172), .B(n_247), .Y(n_246) );
AND2x6_ASAP7_75t_L g144 ( .A(n_9), .B(n_145), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_10), .A2(n_144), .B(n_147), .C(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g541 ( .A(n_11), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_12), .B(n_115), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_12), .B(n_42), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_13), .B(n_185), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_14), .A2(n_104), .B1(n_116), .B2(n_740), .Y(n_103) );
INVx1_ASAP7_75t_L g165 ( .A(n_15), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_16), .B(n_180), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_17), .A2(n_181), .B(n_561), .C(n_563), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_18), .B(n_170), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_19), .B(n_159), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g146 ( .A1(n_20), .A2(n_147), .B(n_150), .C(n_158), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_21), .A2(n_184), .B(n_240), .C(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_22), .B(n_185), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_23), .A2(n_41), .B1(n_730), .B2(n_731), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_23), .Y(n_731) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_24), .B(n_185), .Y(n_515) );
CKINVDCx16_ASAP7_75t_R g475 ( .A(n_25), .Y(n_475) );
INVx1_ASAP7_75t_L g514 ( .A(n_26), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_27), .A2(n_147), .B(n_158), .C(n_250), .Y(n_249) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_28), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_29), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_30), .A2(n_79), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_30), .Y(n_128) );
INVx1_ASAP7_75t_L g492 ( .A(n_31), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_32), .A2(n_139), .B(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g142 ( .A(n_33), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_34), .A2(n_198), .B(n_199), .C(n_203), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_35), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_36), .A2(n_184), .B(n_504), .C(n_506), .Y(n_503) );
INVxp67_ASAP7_75t_L g493 ( .A(n_37), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_38), .B(n_252), .Y(n_251) );
CKINVDCx14_ASAP7_75t_R g502 ( .A(n_39), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_40), .A2(n_147), .B(n_158), .C(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_41), .Y(n_730) );
INVx1_ASAP7_75t_L g115 ( .A(n_42), .Y(n_115) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_43), .A2(n_186), .B(n_539), .C(n_540), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_44), .B(n_138), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_45), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_46), .B(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_47), .B(n_180), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_48), .B(n_139), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_49), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_50), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_51), .A2(n_198), .B(n_203), .C(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g183 ( .A(n_52), .Y(n_183) );
INVx1_ASAP7_75t_L g226 ( .A(n_53), .Y(n_226) );
INVx1_ASAP7_75t_L g547 ( .A(n_54), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_55), .B(n_139), .Y(n_223) );
AOI222xp33_ASAP7_75t_L g457 ( .A1(n_56), .A2(n_458), .B1(n_725), .B2(n_726), .C1(n_732), .C2(n_737), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_57), .Y(n_167) );
CKINVDCx14_ASAP7_75t_R g537 ( .A(n_58), .Y(n_537) );
INVx1_ASAP7_75t_L g145 ( .A(n_59), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_60), .B(n_139), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_61), .B(n_170), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_62), .A2(n_157), .B(n_213), .C(n_215), .Y(n_212) );
INVx1_ASAP7_75t_L g164 ( .A(n_63), .Y(n_164) );
INVx1_ASAP7_75t_SL g505 ( .A(n_64), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_65), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_66), .B(n_180), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_67), .B(n_170), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_68), .B(n_181), .Y(n_237) );
INVx1_ASAP7_75t_L g478 ( .A(n_69), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g176 ( .A(n_70), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_71), .B(n_152), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_72), .A2(n_147), .B(n_203), .C(n_266), .Y(n_265) );
CKINVDCx16_ASAP7_75t_R g211 ( .A(n_73), .Y(n_211) );
INVx1_ASAP7_75t_L g112 ( .A(n_74), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_75), .A2(n_139), .B(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_76), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_77), .A2(n_139), .B(n_558), .Y(n_557) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_78), .A2(n_125), .B1(n_126), .B2(n_129), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_78), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_79), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_80), .A2(n_138), .B(n_488), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g511 ( .A(n_81), .Y(n_511) );
INVx1_ASAP7_75t_L g559 ( .A(n_82), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_83), .B(n_155), .Y(n_154) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_84), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_84), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_85), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_86), .A2(n_139), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g562 ( .A(n_87), .Y(n_562) );
INVx2_ASAP7_75t_L g162 ( .A(n_88), .Y(n_162) );
INVx1_ASAP7_75t_L g529 ( .A(n_89), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_90), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_91), .B(n_185), .Y(n_238) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_92), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g448 ( .A(n_92), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g461 ( .A(n_92), .B(n_450), .Y(n_461) );
INVx2_ASAP7_75t_L g463 ( .A(n_92), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_93), .A2(n_147), .B(n_203), .C(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_94), .B(n_139), .Y(n_196) );
INVx1_ASAP7_75t_L g200 ( .A(n_95), .Y(n_200) );
INVxp67_ASAP7_75t_L g216 ( .A(n_96), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_97), .B(n_172), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g233 ( .A(n_99), .Y(n_233) );
INVx1_ASAP7_75t_L g267 ( .A(n_100), .Y(n_267) );
INVx2_ASAP7_75t_L g550 ( .A(n_101), .Y(n_550) );
AND2x2_ASAP7_75t_L g228 ( .A(n_102), .B(n_161), .Y(n_228) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx5_ASAP7_75t_SL g740 ( .A(n_106), .Y(n_740) );
AND2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_113), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g450 ( .A(n_109), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVxp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_456), .Y(n_116) );
BUFx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_118), .B(n_452), .C(n_457), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_445), .B(n_452), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_130), .B1(n_443), .B2(n_444), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_124), .Y(n_443) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g444 ( .A(n_130), .Y(n_444) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_130), .A2(n_733), .B1(n_734), .B2(n_735), .Y(n_732) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_131), .B(n_379), .Y(n_130) );
NOR5xp2_ASAP7_75t_L g131 ( .A(n_132), .B(n_310), .C(n_339), .D(n_359), .E(n_366), .Y(n_131) );
OAI211xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_190), .B(n_254), .C(n_297), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_134), .A2(n_382), .B1(n_384), .B2(n_385), .Y(n_381) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_169), .Y(n_134) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_135), .Y(n_257) );
AND2x4_ASAP7_75t_L g290 ( .A(n_135), .B(n_291), .Y(n_290) );
INVx5_ASAP7_75t_L g308 ( .A(n_135), .Y(n_308) );
AND2x2_ASAP7_75t_L g317 ( .A(n_135), .B(n_309), .Y(n_317) );
AND2x2_ASAP7_75t_L g329 ( .A(n_135), .B(n_194), .Y(n_329) );
AND2x2_ASAP7_75t_L g425 ( .A(n_135), .B(n_293), .Y(n_425) );
OR2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_166), .Y(n_135) );
AOI21xp5_ASAP7_75t_SL g136 ( .A1(n_137), .A2(n_146), .B(n_159), .Y(n_136) );
BUFx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_144), .Y(n_139) );
NAND2x1p5_ASAP7_75t_L g234 ( .A(n_140), .B(n_144), .Y(n_234) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
INVx1_ASAP7_75t_L g157 ( .A(n_141), .Y(n_157) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
INVx1_ASAP7_75t_L g241 ( .A(n_142), .Y(n_241) );
INVx1_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_143), .Y(n_153) );
INVx3_ASAP7_75t_L g181 ( .A(n_143), .Y(n_181) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_143), .Y(n_185) );
INVx1_ASAP7_75t_L g252 ( .A(n_143), .Y(n_252) );
BUFx3_ASAP7_75t_L g158 ( .A(n_144), .Y(n_158) );
INVx4_ASAP7_75t_SL g188 ( .A(n_144), .Y(n_188) );
INVx5_ASAP7_75t_L g177 ( .A(n_147), .Y(n_177) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
BUFx3_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_148), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_154), .B(n_156), .Y(n_150) );
INVx2_ASAP7_75t_L g155 ( .A(n_152), .Y(n_155) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx4_ASAP7_75t_L g214 ( .A(n_153), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_155), .A2(n_200), .B(n_201), .C(n_202), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_155), .A2(n_202), .B(n_226), .C(n_227), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_155), .A2(n_478), .B(n_479), .C(n_480), .Y(n_477) );
O2A1O1Ixp5_ASAP7_75t_L g528 ( .A1(n_155), .A2(n_480), .B(n_529), .C(n_530), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_156), .A2(n_180), .B(n_514), .C(n_515), .Y(n_513) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_157), .B(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_160), .B(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g168 ( .A(n_161), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_161), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_161), .A2(n_223), .B(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_161), .A2(n_234), .B(n_511), .C(n_512), .Y(n_510) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_161), .A2(n_535), .B(n_542), .Y(n_534) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_162), .B(n_163), .Y(n_161) );
AND2x2_ASAP7_75t_L g173 ( .A(n_162), .B(n_163), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_168), .A2(n_525), .B(n_531), .Y(n_524) );
INVx2_ASAP7_75t_L g291 ( .A(n_169), .Y(n_291) );
AND2x2_ASAP7_75t_L g309 ( .A(n_169), .B(n_263), .Y(n_309) );
AND2x2_ASAP7_75t_L g328 ( .A(n_169), .B(n_262), .Y(n_328) );
AND2x2_ASAP7_75t_L g368 ( .A(n_169), .B(n_308), .Y(n_368) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_174), .B(n_189), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_171), .B(n_205), .Y(n_204) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_171), .A2(n_232), .B(n_242), .Y(n_231) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_171), .A2(n_264), .B(n_272), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_171), .B(n_273), .Y(n_272) );
AO21x2_ASAP7_75t_L g473 ( .A1(n_171), .A2(n_474), .B(n_481), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_171), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_171), .B(n_532), .Y(n_531) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_172), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_172), .A2(n_248), .B(n_249), .Y(n_247) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g244 ( .A(n_173), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_SL g175 ( .A1(n_176), .A2(n_177), .B(n_178), .C(n_188), .Y(n_175) );
INVx2_ASAP7_75t_L g198 ( .A(n_177), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_177), .A2(n_188), .B(n_211), .C(n_212), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_SL g488 ( .A1(n_177), .A2(n_188), .B(n_489), .C(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_177), .A2(n_188), .B(n_502), .C(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_SL g536 ( .A1(n_177), .A2(n_188), .B(n_537), .C(n_538), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_SL g546 ( .A1(n_177), .A2(n_188), .B(n_547), .C(n_548), .Y(n_546) );
O2A1O1Ixp33_ASAP7_75t_SL g558 ( .A1(n_177), .A2(n_188), .B(n_559), .C(n_560), .Y(n_558) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_180), .B(n_216), .Y(n_215) );
OAI22xp33_ASAP7_75t_L g491 ( .A1(n_180), .A2(n_214), .B1(n_492), .B2(n_493), .Y(n_491) );
INVx5_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_181), .B(n_541), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_183), .B(n_184), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_184), .B(n_505), .Y(n_504) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g539 ( .A(n_185), .Y(n_539) );
INVx2_ASAP7_75t_L g480 ( .A(n_186), .Y(n_480) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_187), .Y(n_202) );
INVx1_ASAP7_75t_L g563 ( .A(n_187), .Y(n_563) );
INVx1_ASAP7_75t_L g203 ( .A(n_188), .Y(n_203) );
INVxp67_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_192), .B(n_218), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AOI322xp5_ASAP7_75t_L g427 ( .A1(n_193), .A2(n_229), .A3(n_282), .B1(n_290), .B2(n_344), .C1(n_428), .C2(n_431), .Y(n_427) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_206), .Y(n_193) );
INVx5_ASAP7_75t_L g259 ( .A(n_194), .Y(n_259) );
AND2x2_ASAP7_75t_L g276 ( .A(n_194), .B(n_261), .Y(n_276) );
BUFx2_ASAP7_75t_L g354 ( .A(n_194), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_194), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g431 ( .A(n_194), .B(n_338), .Y(n_431) );
OR2x6_ASAP7_75t_L g194 ( .A(n_195), .B(n_204), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_206), .B(n_220), .Y(n_285) );
INVx1_ASAP7_75t_L g312 ( .A(n_206), .Y(n_312) );
AND2x2_ASAP7_75t_L g325 ( .A(n_206), .B(n_245), .Y(n_325) );
AND2x2_ASAP7_75t_L g426 ( .A(n_206), .B(n_344), .Y(n_426) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OR2x2_ASAP7_75t_L g280 ( .A(n_207), .B(n_220), .Y(n_280) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_207), .Y(n_288) );
OR2x2_ASAP7_75t_L g295 ( .A(n_207), .B(n_245), .Y(n_295) );
AND2x2_ASAP7_75t_L g305 ( .A(n_207), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_207), .B(n_231), .Y(n_334) );
INVxp67_ASAP7_75t_L g358 ( .A(n_207), .Y(n_358) );
AND2x2_ASAP7_75t_L g365 ( .A(n_207), .B(n_229), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_207), .B(n_245), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_207), .B(n_230), .Y(n_391) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_217), .Y(n_207) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_208), .A2(n_500), .B(n_507), .Y(n_499) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_208), .A2(n_545), .B(n_551), .Y(n_544) );
OA21x2_ASAP7_75t_L g556 ( .A1(n_208), .A2(n_557), .B(n_564), .Y(n_556) );
O2A1O1Ixp33_ASAP7_75t_L g266 ( .A1(n_213), .A2(n_267), .B(n_268), .C(n_269), .Y(n_266) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_214), .B(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_214), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_229), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_220), .B(n_246), .Y(n_335) );
OR2x2_ASAP7_75t_L g357 ( .A(n_220), .B(n_230), .Y(n_357) );
AND2x2_ASAP7_75t_L g370 ( .A(n_220), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_220), .B(n_325), .Y(n_376) );
OAI211xp5_ASAP7_75t_SL g380 ( .A1(n_220), .A2(n_381), .B(n_386), .C(n_395), .Y(n_380) );
AND2x2_ASAP7_75t_L g441 ( .A(n_220), .B(n_245), .Y(n_441) );
INVx5_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
OR2x2_ASAP7_75t_L g294 ( .A(n_221), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_221), .B(n_300), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_221), .B(n_289), .Y(n_301) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_221), .Y(n_303) );
OR2x2_ASAP7_75t_L g314 ( .A(n_221), .B(n_230), .Y(n_314) );
AND2x2_ASAP7_75t_SL g319 ( .A(n_221), .B(n_305), .Y(n_319) );
AND2x2_ASAP7_75t_L g344 ( .A(n_221), .B(n_230), .Y(n_344) );
AND2x2_ASAP7_75t_L g364 ( .A(n_221), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g402 ( .A(n_221), .B(n_229), .Y(n_402) );
OR2x2_ASAP7_75t_L g405 ( .A(n_221), .B(n_391), .Y(n_405) );
OR2x6_ASAP7_75t_L g221 ( .A(n_222), .B(n_228), .Y(n_221) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_245), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g348 ( .A1(n_230), .A2(n_349), .B(n_352), .C(n_358), .Y(n_348) );
INVx5_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_231), .B(n_245), .Y(n_279) );
AND2x2_ASAP7_75t_L g283 ( .A(n_231), .B(n_246), .Y(n_283) );
OR2x2_ASAP7_75t_L g289 ( .A(n_231), .B(n_245), .Y(n_289) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_235), .Y(n_232) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_234), .A2(n_475), .B(n_476), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_234), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_239), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_239), .A2(n_251), .B(n_253), .Y(n_250) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx2_ASAP7_75t_L g485 ( .A(n_244), .Y(n_485) );
INVx1_ASAP7_75t_SL g306 ( .A(n_245), .Y(n_306) );
OR2x2_ASAP7_75t_L g434 ( .A(n_245), .B(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_274), .B(n_277), .C(n_286), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AOI31xp33_ASAP7_75t_L g359 ( .A1(n_256), .A2(n_360), .A3(n_362), .B(n_363), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_257), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_258), .B(n_290), .Y(n_296) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_259), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g316 ( .A(n_259), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g321 ( .A(n_259), .B(n_291), .Y(n_321) );
AND2x2_ASAP7_75t_L g331 ( .A(n_259), .B(n_290), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_259), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g351 ( .A(n_259), .B(n_308), .Y(n_351) );
AND2x2_ASAP7_75t_L g356 ( .A(n_259), .B(n_328), .Y(n_356) );
OR2x2_ASAP7_75t_L g375 ( .A(n_259), .B(n_261), .Y(n_375) );
OR2x2_ASAP7_75t_L g377 ( .A(n_259), .B(n_378), .Y(n_377) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_259), .Y(n_424) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g324 ( .A(n_261), .B(n_291), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_261), .B(n_308), .Y(n_347) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx2_ASAP7_75t_L g293 ( .A(n_263), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_271), .Y(n_264) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx3_ASAP7_75t_L g506 ( .A(n_270), .Y(n_506) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g384 ( .A(n_276), .B(n_308), .Y(n_384) );
AOI322xp5_ASAP7_75t_L g386 ( .A1(n_276), .A2(n_290), .A3(n_328), .B1(n_387), .B2(n_388), .C1(n_389), .C2(n_392), .Y(n_386) );
INVx1_ASAP7_75t_L g394 ( .A(n_276), .Y(n_394) );
NAND2xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
INVx1_ASAP7_75t_SL g388 ( .A(n_278), .Y(n_388) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
OR2x2_ASAP7_75t_L g340 ( .A(n_279), .B(n_285), .Y(n_340) );
INVx1_ASAP7_75t_L g371 ( .A(n_279), .Y(n_371) );
INVx2_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OAI32xp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_290), .A3(n_292), .B1(n_294), .B2(n_296), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
AOI21xp33_ASAP7_75t_SL g326 ( .A1(n_289), .A2(n_304), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g341 ( .A(n_290), .Y(n_341) );
AND2x4_ASAP7_75t_L g338 ( .A(n_291), .B(n_308), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_291), .B(n_374), .Y(n_373) );
AOI322xp5_ASAP7_75t_L g403 ( .A1(n_292), .A2(n_319), .A3(n_338), .B1(n_371), .B2(n_404), .C1(n_406), .C2(n_407), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g432 ( .A1(n_292), .A2(n_369), .B1(n_433), .B2(n_434), .C(n_436), .Y(n_432) );
AND2x2_ASAP7_75t_L g320 ( .A(n_293), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g300 ( .A(n_295), .Y(n_300) );
OR2x2_ASAP7_75t_L g372 ( .A(n_295), .B(n_357), .Y(n_372) );
OAI31xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_301), .A3(n_302), .B(n_307), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_298), .A2(n_331), .B1(n_332), .B2(n_336), .Y(n_330) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g343 ( .A(n_300), .B(n_344), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_302), .A2(n_343), .B1(n_396), .B2(n_399), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g385 ( .A(n_305), .B(n_354), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_305), .B(n_344), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_306), .B(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g419 ( .A(n_306), .B(n_357), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_307), .A2(n_402), .B1(n_415), .B2(n_418), .Y(n_414) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx2_ASAP7_75t_L g323 ( .A(n_308), .Y(n_323) );
AND2x2_ASAP7_75t_L g406 ( .A(n_308), .B(n_328), .Y(n_406) );
OR2x2_ASAP7_75t_L g408 ( .A(n_308), .B(n_375), .Y(n_408) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_308), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_309), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_309), .B(n_354), .Y(n_362) );
OAI211xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_315), .B(n_318), .C(n_330), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_320), .B1(n_322), .B2(n_325), .C(n_326), .Y(n_318) );
INVxp67_ASAP7_75t_L g430 ( .A(n_321), .Y(n_430) );
INVx1_ASAP7_75t_L g397 ( .A(n_322), .Y(n_397) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AND2x2_ASAP7_75t_L g361 ( .A(n_323), .B(n_328), .Y(n_361) );
INVx1_ASAP7_75t_L g378 ( .A(n_324), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_324), .B(n_351), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g393 ( .A(n_328), .Y(n_393) );
AND2x2_ASAP7_75t_L g399 ( .A(n_328), .B(n_354), .Y(n_399) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx1_ASAP7_75t_SL g387 ( .A(n_335), .Y(n_387) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_338), .B(n_374), .Y(n_398) );
OAI221xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_342), .B2(n_345), .C(n_348), .Y(n_339) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g435 ( .A(n_344), .Y(n_435) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g353 ( .A(n_347), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_351), .B(n_410), .Y(n_409) );
AOI21xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_355), .B(n_357), .Y(n_352) );
OAI211xp5_ASAP7_75t_SL g400 ( .A1(n_355), .A2(n_401), .B(n_403), .C(n_409), .Y(n_400) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g412 ( .A(n_357), .Y(n_412) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI222xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B1(n_372), .B2(n_373), .C1(n_376), .C2(n_377), .Y(n_366) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g442 ( .A(n_373), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_374), .B(n_417), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_374), .A2(n_421), .B1(n_423), .B2(n_426), .Y(n_420) );
INVx2_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
NOR4xp25_ASAP7_75t_L g379 ( .A(n_380), .B(n_400), .C(n_413), .D(n_432), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_382), .B(n_412), .Y(n_422) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g389 ( .A(n_387), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_390), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_420), .C(n_427), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx2_ASAP7_75t_L g429 ( .A(n_425), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
OAI21xp5_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_439), .B(n_442), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_444), .A2(n_459), .B1(n_462), .B2(n_464), .Y(n_458) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g455 ( .A(n_448), .Y(n_455) );
NOR2x2_ASAP7_75t_L g739 ( .A(n_449), .B(n_463), .Y(n_739) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g462 ( .A(n_450), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g733 ( .A(n_460), .Y(n_733) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g736 ( .A(n_462), .Y(n_736) );
INVx2_ASAP7_75t_L g734 ( .A(n_464), .Y(n_734) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_659), .Y(n_464) );
NAND5xp2_ASAP7_75t_L g465 ( .A(n_466), .B(n_588), .C(n_618), .D(n_639), .E(n_645), .Y(n_465) );
AOI221xp5_ASAP7_75t_SL g466 ( .A1(n_467), .A2(n_521), .B1(n_552), .B2(n_554), .C(n_565), .Y(n_466) );
INVxp67_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_518), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_496), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_SL g639 ( .A1(n_471), .A2(n_508), .B(n_640), .C(n_643), .Y(n_639) );
AND2x2_ASAP7_75t_L g709 ( .A(n_471), .B(n_509), .Y(n_709) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_483), .Y(n_471) );
AND2x2_ASAP7_75t_L g567 ( .A(n_472), .B(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g571 ( .A(n_472), .B(n_568), .Y(n_571) );
OR2x2_ASAP7_75t_L g597 ( .A(n_472), .B(n_509), .Y(n_597) );
AND2x2_ASAP7_75t_L g599 ( .A(n_472), .B(n_499), .Y(n_599) );
AND2x2_ASAP7_75t_L g617 ( .A(n_472), .B(n_498), .Y(n_617) );
INVx1_ASAP7_75t_L g650 ( .A(n_472), .Y(n_650) );
INVx2_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
BUFx2_ASAP7_75t_L g520 ( .A(n_473), .Y(n_520) );
AND2x2_ASAP7_75t_L g553 ( .A(n_473), .B(n_499), .Y(n_553) );
AND2x2_ASAP7_75t_L g706 ( .A(n_473), .B(n_509), .Y(n_706) );
AND2x2_ASAP7_75t_L g587 ( .A(n_483), .B(n_497), .Y(n_587) );
OR2x2_ASAP7_75t_L g591 ( .A(n_483), .B(n_509), .Y(n_591) );
AND2x2_ASAP7_75t_L g616 ( .A(n_483), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_SL g663 ( .A(n_483), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_483), .B(n_625), .Y(n_711) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_486), .B(n_494), .Y(n_483) );
INVx1_ASAP7_75t_L g569 ( .A(n_484), .Y(n_569) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OA21x2_ASAP7_75t_L g568 ( .A1(n_487), .A2(n_495), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
OAI322xp33_ASAP7_75t_L g712 ( .A1(n_496), .A2(n_648), .A3(n_671), .B1(n_692), .B2(n_713), .C1(n_715), .C2(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_497), .B(n_568), .Y(n_715) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_508), .Y(n_497) );
AND2x2_ASAP7_75t_L g519 ( .A(n_498), .B(n_520), .Y(n_519) );
AND2x4_ASAP7_75t_L g584 ( .A(n_498), .B(n_509), .Y(n_584) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g625 ( .A(n_499), .B(n_509), .Y(n_625) );
AND2x2_ASAP7_75t_L g669 ( .A(n_499), .B(n_508), .Y(n_669) );
AND2x2_ASAP7_75t_L g552 ( .A(n_508), .B(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g570 ( .A(n_508), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_508), .B(n_599), .Y(n_723) );
INVx3_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g518 ( .A(n_509), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_509), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g637 ( .A(n_509), .B(n_568), .Y(n_637) );
AND2x2_ASAP7_75t_L g664 ( .A(n_509), .B(n_599), .Y(n_664) );
OR2x2_ASAP7_75t_L g720 ( .A(n_509), .B(n_571), .Y(n_720) );
OR2x6_ASAP7_75t_L g509 ( .A(n_510), .B(n_516), .Y(n_509) );
INVx1_ASAP7_75t_SL g606 ( .A(n_518), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_519), .B(n_637), .Y(n_638) );
AND2x2_ASAP7_75t_L g672 ( .A(n_519), .B(n_662), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_519), .B(n_595), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_519), .B(n_717), .Y(n_716) );
OAI31xp33_ASAP7_75t_L g690 ( .A1(n_521), .A2(n_552), .A3(n_691), .B(n_693), .Y(n_690) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_533), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_522), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g673 ( .A(n_522), .B(n_608), .Y(n_673) );
OR2x2_ASAP7_75t_L g680 ( .A(n_522), .B(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g692 ( .A(n_522), .B(n_581), .Y(n_692) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
OR2x2_ASAP7_75t_L g626 ( .A(n_523), .B(n_627), .Y(n_626) );
BUFx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g554 ( .A(n_524), .B(n_555), .Y(n_554) );
INVx4_ASAP7_75t_L g575 ( .A(n_524), .Y(n_575) );
AND2x2_ASAP7_75t_L g612 ( .A(n_524), .B(n_556), .Y(n_612) );
AND2x2_ASAP7_75t_L g611 ( .A(n_533), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_SL g681 ( .A(n_533), .Y(n_681) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_543), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_534), .B(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g581 ( .A(n_534), .B(n_544), .Y(n_581) );
INVx2_ASAP7_75t_L g601 ( .A(n_534), .Y(n_601) );
AND2x2_ASAP7_75t_L g615 ( .A(n_534), .B(n_544), .Y(n_615) );
AND2x2_ASAP7_75t_L g622 ( .A(n_534), .B(n_578), .Y(n_622) );
BUFx3_ASAP7_75t_L g632 ( .A(n_534), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_534), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g577 ( .A(n_543), .Y(n_577) );
AND2x2_ASAP7_75t_L g585 ( .A(n_543), .B(n_575), .Y(n_585) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g555 ( .A(n_544), .B(n_556), .Y(n_555) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_544), .Y(n_609) );
INVx2_ASAP7_75t_SL g592 ( .A(n_553), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_553), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_553), .B(n_662), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_554), .B(n_632), .Y(n_685) );
INVx1_ASAP7_75t_SL g719 ( .A(n_554), .Y(n_719) );
INVx1_ASAP7_75t_SL g627 ( .A(n_555), .Y(n_627) );
INVx1_ASAP7_75t_SL g578 ( .A(n_556), .Y(n_578) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_556), .Y(n_589) );
OR2x2_ASAP7_75t_L g600 ( .A(n_556), .B(n_575), .Y(n_600) );
AND2x2_ASAP7_75t_L g614 ( .A(n_556), .B(n_575), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_556), .B(n_604), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_570), .B(n_572), .C(n_583), .Y(n_565) );
AOI31xp33_ASAP7_75t_L g682 ( .A1(n_566), .A2(n_683), .A3(n_684), .B(n_685), .Y(n_682) );
AND2x2_ASAP7_75t_L g655 ( .A(n_567), .B(n_584), .Y(n_655) );
BUFx3_ASAP7_75t_L g595 ( .A(n_568), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_568), .B(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g631 ( .A(n_568), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_568), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g586 ( .A(n_571), .Y(n_586) );
OAI222xp33_ASAP7_75t_L g695 ( .A1(n_571), .A2(n_696), .B1(n_699), .B2(n_700), .C1(n_701), .C2(n_702), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_579), .Y(n_572) );
INVx1_ASAP7_75t_L g701 ( .A(n_573), .Y(n_701) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_575), .B(n_578), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_575), .B(n_601), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_575), .B(n_576), .Y(n_671) );
INVx1_ASAP7_75t_L g722 ( .A(n_575), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_576), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g724 ( .A(n_576), .Y(n_724) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx2_ASAP7_75t_L g604 ( .A(n_577), .Y(n_604) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_578), .Y(n_647) );
AOI32xp33_ASAP7_75t_L g583 ( .A1(n_579), .A2(n_584), .A3(n_585), .B1(n_586), .B2(n_587), .Y(n_583) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_581), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g658 ( .A(n_581), .Y(n_658) );
OR2x2_ASAP7_75t_L g699 ( .A(n_581), .B(n_600), .Y(n_699) );
INVx1_ASAP7_75t_L g635 ( .A(n_582), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_584), .B(n_595), .Y(n_620) );
INVx3_ASAP7_75t_L g629 ( .A(n_584), .Y(n_629) );
AOI322xp5_ASAP7_75t_L g645 ( .A1(n_584), .A2(n_629), .A3(n_646), .B1(n_648), .B2(n_651), .C1(n_655), .C2(n_656), .Y(n_645) );
AND2x2_ASAP7_75t_L g621 ( .A(n_585), .B(n_622), .Y(n_621) );
INVxp67_ASAP7_75t_L g698 ( .A(n_585), .Y(n_698) );
A2O1A1O1Ixp25_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B(n_593), .C(n_601), .D(n_602), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_589), .B(n_632), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
OAI221xp5_ASAP7_75t_L g602 ( .A1(n_591), .A2(n_603), .B1(n_606), .B2(n_607), .C(n_610), .Y(n_602) );
INVx1_ASAP7_75t_SL g717 ( .A(n_591), .Y(n_717) );
AOI21xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_598), .B(n_600), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_595), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI221xp5_ASAP7_75t_SL g687 ( .A1(n_597), .A2(n_681), .B1(n_688), .B2(n_689), .C(n_690), .Y(n_687) );
OAI222xp33_ASAP7_75t_L g718 ( .A1(n_598), .A2(n_719), .B1(n_720), .B2(n_721), .C1(n_723), .C2(n_724), .Y(n_718) );
AND2x2_ASAP7_75t_L g676 ( .A(n_599), .B(n_662), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_599), .A2(n_614), .B(n_661), .Y(n_688) );
INVx1_ASAP7_75t_L g702 ( .A(n_599), .Y(n_702) );
INVx2_ASAP7_75t_SL g605 ( .A(n_600), .Y(n_605) );
AND2x2_ASAP7_75t_L g608 ( .A(n_601), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_SL g642 ( .A(n_604), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_604), .B(n_614), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_605), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_605), .B(n_615), .Y(n_644) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OAI21xp5_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_613), .B(n_616), .Y(n_610) );
INVx1_ASAP7_75t_SL g628 ( .A(n_612), .Y(n_628) );
AND2x2_ASAP7_75t_L g675 ( .A(n_612), .B(n_658), .Y(n_675) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
AND2x2_ASAP7_75t_L g714 ( .A(n_614), .B(n_632), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_615), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g700 ( .A(n_616), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_621), .B1(n_623), .B2(n_630), .C(n_633), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_626), .B1(n_628), .B2(n_629), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI22xp33_ASAP7_75t_L g633 ( .A1(n_627), .A2(n_634), .B1(n_636), .B2(n_638), .Y(n_633) );
OR2x2_ASAP7_75t_L g704 ( .A(n_628), .B(n_632), .Y(n_704) );
OR2x2_ASAP7_75t_L g707 ( .A(n_628), .B(n_642), .Y(n_707) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OAI221xp5_ASAP7_75t_L g703 ( .A1(n_649), .A2(n_704), .B1(n_705), .B2(n_707), .C(n_708), .Y(n_703) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND3xp33_ASAP7_75t_SL g659 ( .A(n_660), .B(n_674), .C(n_686), .Y(n_659) );
AOI222xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_665), .B1(n_667), .B2(n_670), .C1(n_672), .C2(n_673), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_662), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g684 ( .A(n_664), .Y(n_684) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVxp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B1(n_677), .B2(n_679), .C(n_682), .Y(n_674) );
INVx1_ASAP7_75t_L g689 ( .A(n_675), .Y(n_689) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OAI21xp33_ASAP7_75t_L g708 ( .A1(n_679), .A2(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
NOR5xp2_ASAP7_75t_L g686 ( .A(n_687), .B(n_695), .C(n_703), .D(n_712), .E(n_718), .Y(n_686) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OR2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVxp67_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx3_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
endmodule