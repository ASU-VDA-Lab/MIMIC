module real_jpeg_18379_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_412;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_1),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_2),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_2),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_2),
.A2(n_99),
.B1(n_131),
.B2(n_278),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_2),
.A2(n_99),
.B1(n_342),
.B2(n_343),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_2),
.A2(n_99),
.B1(n_399),
.B2(n_402),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_3),
.A2(n_158),
.B1(n_162),
.B2(n_167),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_3),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_3),
.A2(n_167),
.B1(n_242),
.B2(n_263),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_4),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_4),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_4),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g378 ( 
.A(n_4),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_5),
.Y(n_144)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_5),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g423 ( 
.A(n_5),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_6),
.A2(n_146),
.B1(n_150),
.B2(n_153),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_6),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_6),
.A2(n_153),
.B1(n_238),
.B2(n_241),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_7),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_7),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_7),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_7),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_7),
.Y(n_340)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_7),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_8),
.A2(n_96),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_8),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_8),
.A2(n_111),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_8),
.A2(n_111),
.B1(n_159),
.B2(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_9),
.Y(n_134)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_10),
.A2(n_114),
.A3(n_117),
.B1(n_121),
.B2(n_129),
.Y(n_113)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_10),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_10),
.A2(n_128),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_10),
.B(n_35),
.Y(n_297)
);

OAI32xp33_ASAP7_75t_L g316 ( 
.A1(n_10),
.A2(n_317),
.A3(n_321),
.B1(n_322),
.B2(n_325),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_10),
.A2(n_128),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_10),
.B(n_65),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_10),
.B(n_423),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_10),
.B(n_200),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_11),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_23)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_11),
.A2(n_29),
.B1(n_300),
.B2(n_304),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_11),
.A2(n_29),
.B1(n_388),
.B2(n_394),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_11),
.A2(n_29),
.B1(n_425),
.B2(n_429),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_13),
.A2(n_202),
.B1(n_203),
.B2(n_205),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_13),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_13),
.A2(n_202),
.B1(n_227),
.B2(n_231),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_13),
.A2(n_202),
.B1(n_272),
.B2(n_274),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_14),
.Y(n_140)
);

BUFx4f_ASAP7_75t_L g149 ( 
.A(n_14),
.Y(n_149)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_14),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_14),
.Y(n_186)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_283),
.Y(n_16)
);

OAI21xp33_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_246),
.B(n_281),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_18),
.B(n_247),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_168),
.C(n_223),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_19),
.B(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_112),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_62),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_21),
.B(n_62),
.C(n_112),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_33),
.B1(n_35),
.B2(n_55),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_23),
.A2(n_34),
.B1(n_211),
.B2(n_215),
.Y(n_210)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_26),
.Y(n_214)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_27),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_28),
.Y(n_120)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_31),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_56)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_34),
.A2(n_56),
.B1(n_215),
.B2(n_277),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_45),
.Y(n_34)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_35),
.Y(n_215)
);

AO22x2_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_35)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_36),
.Y(n_352)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_37),
.Y(n_305)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_37),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_42),
.Y(n_273)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_57),
.A2(n_61),
.B1(n_218),
.B2(n_222),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_57),
.A2(n_61),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_57),
.A2(n_61),
.B1(n_162),
.B2(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_60),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_93),
.B(n_106),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_64),
.A2(n_94),
.B1(n_107),
.B2(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_64),
.A2(n_108),
.B(n_270),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_64),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_64),
.A2(n_107),
.B1(n_299),
.B2(n_346),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_78),
.Y(n_64)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_65),
.B(n_271),
.Y(n_270)
);

AO22x2_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B1(n_72),
.B2(n_75),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_71),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_71),
.Y(n_324)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_73),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_73),
.Y(n_264)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_73),
.Y(n_337)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_74),
.Y(n_193)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_74),
.Y(n_244)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_83),
.B1(n_86),
.B2(n_89),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_85),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_85),
.Y(n_275)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_97),
.Y(n_222)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_97),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_103),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_107),
.Y(n_307)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_109),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_135),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_113),
.B(n_135),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_128),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_128),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_128),
.B(n_182),
.Y(n_375)
);

OAI21xp33_ASAP7_75t_SL g384 ( 
.A1(n_128),
.A2(n_375),
.B(n_385),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_128),
.A2(n_137),
.B1(n_422),
.B2(n_424),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_145),
.B1(n_154),
.B2(n_157),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_136),
.A2(n_157),
.B(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_136),
.A2(n_225),
.B(n_332),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_136),
.A2(n_411),
.B1(n_415),
.B2(n_416),
.Y(n_410)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_137),
.B(n_226),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_137),
.A2(n_398),
.B(n_404),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_137),
.A2(n_412),
.B1(n_424),
.B2(n_437),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_140),
.Y(n_258)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_142),
.B(n_226),
.Y(n_225)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_143),
.Y(n_439)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_145),
.A2(n_259),
.B(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_148),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_149),
.Y(n_230)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_149),
.Y(n_401)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_149),
.Y(n_428)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_156),
.Y(n_256)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_160),
.Y(n_403)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_160),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_161),
.Y(n_166)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_164),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_168),
.B(n_223),
.Y(n_309)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_210),
.C(n_216),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_169),
.B(n_216),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_191),
.B(n_199),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_170),
.A2(n_183),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_170),
.A2(n_183),
.B1(n_334),
.B2(n_341),
.Y(n_333)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_171),
.B(n_201),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_171),
.A2(n_357),
.B(n_358),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_171),
.A2(n_200),
.B1(n_384),
.B2(n_387),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_171),
.A2(n_200),
.B1(n_335),
.B2(n_387),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_183),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_176),
.B1(n_178),
.B2(n_182),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_174),
.Y(n_370)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_175),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_175),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx8_ASAP7_75t_L g374 ( 
.A(n_177),
.Y(n_374)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_182),
.Y(n_344)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_183),
.B(n_191),
.Y(n_358)
);

OA22x2_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_186),
.Y(n_381)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_197),
.Y(n_321)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_200),
.B(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_210),
.B(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_217),
.A2(n_299),
.B1(n_306),
.B2(n_307),
.Y(n_298)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_235),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_224),
.B(n_235),
.Y(n_267)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_245),
.Y(n_235)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

BUFx2_ASAP7_75t_SL g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_265),
.B1(n_266),
.B2(n_280),
.Y(n_249)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_260),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_259),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_252),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx4_ASAP7_75t_SL g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_255),
.Y(n_295)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_255),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_257),
.Y(n_332)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_258),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_276),
.Y(n_268)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_310),
.B(n_456),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_308),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_286),
.B(n_308),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.C(n_291),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_287),
.B(n_452),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_291),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_296),
.C(n_298),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_292),
.A2(n_296),
.B1(n_297),
.B2(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_292),
.Y(n_362)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_298),
.B(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI21x1_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_450),
.B(n_455),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_364),
.B(n_449),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_353),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_314),
.B(n_353),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_333),
.C(n_345),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_315),
.B(n_447),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_331),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_316),
.B(n_331),
.Y(n_355)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_333),
.B(n_345),
.Y(n_447)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_341),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_342),
.Y(n_386)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_359),
.B1(n_360),
.B2(n_363),
.Y(n_353)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_354),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_355),
.B(n_356),
.C(n_359),
.Y(n_454)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_444),
.B(n_448),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_408),
.B(n_443),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_396),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_367),
.B(n_396),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_382),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_368),
.A2(n_382),
.B1(n_383),
.B2(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_368),
.Y(n_418)
);

OAI32xp33_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_371),
.A3(n_372),
.B1(n_375),
.B2(n_376),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_379),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_405),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_397),
.B(n_406),
.C(n_407),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_398),
.Y(n_415)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

OAI21x1_ASAP7_75t_SL g408 ( 
.A1(n_409),
.A2(n_419),
.B(n_442),
.Y(n_408)
);

NOR2x1_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_417),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_410),
.B(n_417),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_435),
.B(n_441),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_430),
.Y(n_420)
);

BUFx12f_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_434),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_436),
.B(n_440),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_436),
.B(n_440),
.Y(n_441)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx5_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_445),
.B(n_446),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_454),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_451),
.B(n_454),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);


endmodule