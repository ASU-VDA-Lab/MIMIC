module fake_jpeg_3415_n_291 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_291);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_45),
.B(n_49),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_47),
.B(n_57),
.Y(n_77)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_51),
.B(n_53),
.Y(n_98)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_0),
.C(n_2),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_32),
.Y(n_81)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_15),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_59),
.Y(n_100)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_30),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_32),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_3),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_4),
.Y(n_83)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_31),
.B1(n_20),
.B2(n_35),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_67),
.A2(n_78),
.B1(n_37),
.B2(n_33),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_20),
.B1(n_35),
.B2(n_27),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_69),
.A2(n_56),
.B(n_28),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_24),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_74),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_26),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_79),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_31),
.B1(n_27),
.B2(n_17),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_83),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_23),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_29),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_94),
.Y(n_110)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_39),
.B1(n_25),
.B2(n_23),
.Y(n_93)
);

AO22x2_ASAP7_75t_L g131 ( 
.A1(n_93),
.A2(n_100),
.B1(n_92),
.B2(n_101),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_29),
.Y(n_94)
);

BUFx16f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_17),
.C(n_36),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_54),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_102),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_46),
.B(n_36),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_41),
.B(n_22),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_62),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_107),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_46),
.B(n_22),
.Y(n_107)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_62),
.C(n_37),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_108),
.B(n_122),
.C(n_95),
.Y(n_171)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

NAND2xp33_ASAP7_75t_SL g157 ( 
.A(n_113),
.B(n_131),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_115),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_135),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_28),
.B(n_63),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_132),
.B(n_136),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_46),
.C(n_42),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_39),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_42),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_130),
.B(n_142),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_98),
.A2(n_65),
.B(n_48),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_4),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_8),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_37),
.B(n_34),
.C(n_9),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_137),
.B(n_139),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_70),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_93),
.A2(n_50),
.B(n_34),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_96),
.A2(n_50),
.B1(n_37),
.B2(n_33),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_71),
.B1(n_91),
.B2(n_90),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g139 ( 
.A1(n_96),
.A2(n_37),
.A3(n_33),
.B1(n_9),
.B2(n_10),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_70),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_87),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g141 ( 
.A1(n_69),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_141),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_73),
.B(n_5),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_173),
.B1(n_114),
.B2(n_115),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_80),
.B1(n_106),
.B2(n_75),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_146),
.A2(n_140),
.B1(n_135),
.B2(n_143),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_86),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_167),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_150),
.B(n_165),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_95),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_154),
.B(n_159),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_71),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_174),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_106),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_166),
.B(n_115),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_112),
.B(n_87),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_123),
.B(n_84),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_175),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_172),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_117),
.B(n_75),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_110),
.B(n_91),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_109),
.B(n_90),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_11),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_128),
.Y(n_191)
);

OR2x2_ASAP7_75t_SL g177 ( 
.A(n_171),
.B(n_122),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_177),
.A2(n_155),
.B(n_147),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_156),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_183),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_108),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_127),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_172),
.C(n_162),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_144),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_191),
.Y(n_224)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_190),
.A2(n_173),
.B1(n_148),
.B2(n_163),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_125),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_195),
.B(n_196),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_121),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_144),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_198),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_127),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_147),
.A2(n_134),
.B1(n_141),
.B2(n_131),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_199),
.A2(n_169),
.B1(n_185),
.B2(n_197),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_114),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_202),
.Y(n_210)
);

AND2x6_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_132),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_133),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_205),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

AO22x1_ASAP7_75t_L g205 ( 
.A1(n_157),
.A2(n_131),
.B1(n_139),
.B2(n_113),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_215),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_177),
.C(n_194),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_199),
.A2(n_169),
.B1(n_157),
.B2(n_146),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_214),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_193),
.A2(n_145),
.B1(n_172),
.B2(n_148),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_184),
.B(n_150),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_220),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_131),
.B1(n_158),
.B2(n_153),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_189),
.A2(n_182),
.B(n_192),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_225),
.B(n_227),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_205),
.A2(n_131),
.B1(n_153),
.B2(n_158),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_226),
.B1(n_179),
.B2(n_178),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_189),
.A2(n_160),
.B(n_166),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_160),
.B1(n_164),
.B2(n_165),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_192),
.A2(n_151),
.B(n_152),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_202),
.A2(n_118),
.B1(n_11),
.B2(n_13),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_228),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_180),
.A2(n_186),
.B(n_194),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_212),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_238),
.B1(n_222),
.B2(n_213),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_200),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_231),
.B(n_237),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_234),
.C(n_206),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_183),
.C(n_178),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_181),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_216),
.A2(n_209),
.B1(n_223),
.B2(n_217),
.Y(n_238)
);

OAI322xp33_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_181),
.A3(n_188),
.B1(n_204),
.B2(n_190),
.C1(n_187),
.C2(n_13),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_246),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_224),
.B(n_188),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_245),
.Y(n_260)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_118),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_243),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_254),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_252),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_215),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_255),
.B1(n_258),
.B2(n_240),
.Y(n_268)
);

BUFx12_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_228),
.B1(n_210),
.B2(n_209),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_242),
.A2(n_208),
.B1(n_210),
.B2(n_214),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_226),
.C(n_225),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_232),
.C(n_242),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_248),
.B(n_238),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_265),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_266),
.Y(n_273)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_259),
.A2(n_232),
.B(n_240),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_234),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_265),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_258),
.A2(n_227),
.B(n_241),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_270),
.A2(n_247),
.B1(n_260),
.B2(n_241),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_278),
.C(n_263),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_235),
.B(n_244),
.C(n_249),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_277),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_SL g275 ( 
.A1(n_262),
.A2(n_230),
.B(n_220),
.C(n_218),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_275),
.A2(n_254),
.B(n_276),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_251),
.C(n_252),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_236),
.C(n_219),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_281),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_236),
.C(n_219),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_283),
.A2(n_274),
.B(n_275),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_282),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_272),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_288),
.C(n_286),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_275),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_254),
.Y(n_291)
);


endmodule