module fake_jpeg_1118_n_552 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_552);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_552;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_53),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_55),
.B(n_77),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_24),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_68),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_24),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_64),
.Y(n_120)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_65),
.Y(n_122)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_66),
.Y(n_164)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_28),
.B(n_17),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_70),
.Y(n_162)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g143 ( 
.A(n_73),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_28),
.B(n_18),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_78),
.B(n_88),
.Y(n_134)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_80),
.Y(n_161)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_81),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_31),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_37),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_90),
.B(n_94),
.Y(n_141)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_16),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_43),
.B(n_16),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_97),
.B(n_102),
.Y(n_144)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_14),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_14),
.Y(n_128)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_103),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_19),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_104),
.B(n_105),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_50),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_45),
.B(n_43),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_107),
.B(n_128),
.Y(n_183)
);

OR2x4_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_41),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_117),
.Y(n_185)
);

HAxp5_ASAP7_75t_SL g125 ( 
.A(n_82),
.B(n_41),
.CON(n_125),
.SN(n_125)
);

BUFx8_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

AND2x4_ASAP7_75t_L g129 ( 
.A(n_71),
.B(n_44),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_129),
.B(n_145),
.C(n_46),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_65),
.B(n_43),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_41),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_66),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_135),
.Y(n_175)
);

INVx6_ASAP7_75t_SL g132 ( 
.A(n_95),
.Y(n_132)
);

CKINVDCx12_ASAP7_75t_R g180 ( 
.A(n_132),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_73),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_67),
.A2(n_45),
.B1(n_44),
.B2(n_69),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_151),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_98),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_140),
.B(n_159),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_56),
.A2(n_45),
.B(n_52),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_102),
.A2(n_50),
.B1(n_46),
.B2(n_36),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_148),
.A2(n_80),
.B1(n_92),
.B2(n_86),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_87),
.B(n_46),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_54),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_89),
.A2(n_41),
.B1(n_29),
.B2(n_50),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_163),
.A2(n_41),
.B1(n_29),
.B2(n_85),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_103),
.B(n_23),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_165),
.B(n_34),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_168),
.B(n_170),
.Y(n_247)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_134),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_171),
.Y(n_245)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_173),
.Y(n_275)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_116),
.B(n_115),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_176),
.B(n_186),
.Y(n_256)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_177),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_124),
.Y(n_178)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_178),
.Y(n_243)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_181),
.A2(n_210),
.B1(n_211),
.B2(n_215),
.Y(n_276)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_112),
.Y(n_182)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_182),
.Y(n_273)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_42),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_187),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_188),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_189),
.Y(n_242)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_190),
.Y(n_244)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_191),
.Y(n_259)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_138),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_193),
.Y(n_233)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_194),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_197),
.Y(n_267)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_198),
.Y(n_271)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_146),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_199),
.Y(n_250)
);

AO22x1_ASAP7_75t_SL g200 ( 
.A1(n_117),
.A2(n_72),
.B1(n_96),
.B2(n_62),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_207),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_120),
.B(n_35),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_202),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_120),
.B(n_119),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_122),
.B(n_35),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

CKINVDCx12_ASAP7_75t_R g205 ( 
.A(n_160),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_205),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_122),
.B(n_34),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_208),
.Y(n_240)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_110),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_209),
.B(n_212),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_147),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_114),
.B(n_52),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_214),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_138),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_129),
.A2(n_29),
.B1(n_36),
.B2(n_50),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_106),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_217),
.Y(n_251)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_149),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_108),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_221),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_149),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_219),
.A2(n_220),
.B1(n_224),
.B2(n_225),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_129),
.A2(n_29),
.B1(n_36),
.B2(n_42),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_111),
.B(n_33),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_222),
.B(n_223),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_151),
.B(n_33),
.Y(n_223)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_112),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_160),
.B(n_26),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_226),
.A2(n_227),
.B1(n_123),
.B2(n_118),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_185),
.B(n_144),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_228),
.B(n_254),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_148),
.B1(n_163),
.B2(n_161),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_230),
.A2(n_236),
.B1(n_266),
.B2(n_270),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_144),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_234),
.B(n_248),
.C(n_180),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_167),
.A2(n_152),
.B1(n_161),
.B2(n_155),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_172),
.A2(n_23),
.B1(n_26),
.B2(n_164),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_238),
.A2(n_252),
.B1(n_268),
.B2(n_200),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_183),
.B(n_125),
.C(n_157),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_167),
.A2(n_60),
.B1(n_75),
.B2(n_84),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_185),
.B(n_155),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_175),
.B(n_152),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_262),
.B(n_264),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_167),
.A2(n_139),
.B1(n_123),
.B2(n_118),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_263),
.A2(n_182),
.B1(n_224),
.B2(n_218),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_196),
.B(n_139),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_181),
.A2(n_58),
.B1(n_166),
.B2(n_126),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_215),
.A2(n_166),
.B1(n_126),
.B2(n_108),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_220),
.A2(n_101),
.B(n_83),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_272),
.A2(n_74),
.B(n_188),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_200),
.B(n_160),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_274),
.B(n_217),
.Y(n_311)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_243),
.Y(n_279)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_279),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_280),
.B(n_295),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_282),
.A2(n_292),
.B1(n_323),
.B2(n_5),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_261),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_283),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_284),
.B(n_299),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_232),
.B(n_178),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_285),
.B(n_294),
.Y(n_354)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_237),
.Y(n_286)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_286),
.Y(n_334)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_237),
.Y(n_287)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_287),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_245),
.B(n_193),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_289),
.Y(n_326)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_243),
.Y(n_290)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_290),
.Y(n_344)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_291),
.Y(n_329)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_293),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_245),
.B(n_216),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_260),
.B(n_278),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_275),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_296),
.B(n_297),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_240),
.B(n_260),
.Y(n_297)
);

NOR2x1_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_212),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_298),
.A2(n_244),
.B(n_47),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_258),
.B(n_234),
.C(n_247),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_228),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_300),
.B(n_303),
.Y(n_348)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_246),
.Y(n_302)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_302),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_241),
.B(n_187),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_254),
.B(n_169),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_304),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_197),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_305),
.B(n_313),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_184),
.C(n_179),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_306),
.B(n_317),
.Y(n_366)
);

AND2x6_ASAP7_75t_L g307 ( 
.A(n_258),
.B(n_13),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_307),
.B(n_311),
.Y(n_331)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_308),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_236),
.A2(n_227),
.B1(n_211),
.B2(n_219),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_309),
.A2(n_319),
.B(n_242),
.Y(n_342)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_231),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_256),
.B(n_210),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_312),
.B(n_316),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_235),
.B(n_199),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_229),
.B(n_174),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_314),
.B(n_322),
.Y(n_363)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_246),
.Y(n_315)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_315),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_262),
.B(n_274),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_230),
.B(n_195),
.C(n_189),
.Y(n_317)
);

INVx13_ASAP7_75t_L g318 ( 
.A(n_233),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_318),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_239),
.A2(n_95),
.B1(n_47),
.B2(n_59),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_320),
.A2(n_265),
.B1(n_267),
.B2(n_273),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_239),
.B(n_0),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_321),
.B(n_325),
.Y(n_364)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_229),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_231),
.Y(n_323)
);

A2O1A1O1Ixp25_ASAP7_75t_L g324 ( 
.A1(n_239),
.A2(n_61),
.B(n_47),
.C(n_2),
.D(n_4),
.Y(n_324)
);

A2O1A1Ixp33_ASAP7_75t_L g339 ( 
.A1(n_324),
.A2(n_251),
.B(n_250),
.C(n_267),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_259),
.B(n_0),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_298),
.A2(n_272),
.B(n_276),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_327),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_319),
.A2(n_277),
.B(n_270),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_328),
.B(n_330),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_298),
.A2(n_316),
.B(n_288),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_281),
.A2(n_268),
.B1(n_266),
.B2(n_250),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_338),
.A2(n_340),
.B1(n_345),
.B2(n_361),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_339),
.B(n_352),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_311),
.A2(n_259),
.B1(n_265),
.B2(n_242),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_341),
.A2(n_343),
.B1(n_359),
.B2(n_302),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_347),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_317),
.A2(n_273),
.B1(n_249),
.B2(n_257),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_288),
.A2(n_261),
.B1(n_249),
.B2(n_253),
.Y(n_345)
);

OAI32xp33_ASAP7_75t_L g347 ( 
.A1(n_299),
.A2(n_257),
.A3(n_244),
.B1(n_253),
.B2(n_47),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_349),
.B(n_320),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_301),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_352)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_357),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_301),
.A2(n_5),
.B(n_6),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_358),
.B(n_352),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_321),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_304),
.A2(n_280),
.B1(n_307),
.B2(n_303),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_326),
.B(n_285),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_368),
.B(n_376),
.Y(n_434)
);

OAI32xp33_ASAP7_75t_L g369 ( 
.A1(n_348),
.A2(n_304),
.A3(n_290),
.B1(n_279),
.B2(n_312),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_392),
.Y(n_407)
);

INVx13_ASAP7_75t_L g371 ( 
.A(n_329),
.Y(n_371)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_371),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_284),
.C(n_306),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_372),
.B(n_374),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_353),
.Y(n_373)
);

NOR3xp33_ASAP7_75t_L g425 ( 
.A(n_373),
.B(n_382),
.C(n_388),
.Y(n_425)
);

MAJx2_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_297),
.C(n_322),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_354),
.B(n_296),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_354),
.B(n_293),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_377),
.B(n_385),
.Y(n_415)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_333),
.Y(n_378)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_378),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_380),
.A2(n_349),
.B(n_339),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_363),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_333),
.Y(n_383)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_383),
.Y(n_416)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_344),
.Y(n_384)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_384),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_332),
.B(n_308),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_330),
.B(n_291),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_386),
.B(n_387),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_335),
.B(n_348),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_363),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_335),
.B(n_291),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_400),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_332),
.B(n_310),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_390),
.B(n_397),
.Y(n_422)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_344),
.Y(n_391)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_391),
.Y(n_429)
);

AO22x1_ASAP7_75t_L g392 ( 
.A1(n_361),
.A2(n_324),
.B1(n_286),
.B2(n_287),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_346),
.Y(n_393)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_393),
.Y(n_430)
);

NOR3xp33_ASAP7_75t_L g431 ( 
.A(n_396),
.B(n_398),
.C(n_364),
.Y(n_431)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_346),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_337),
.Y(n_398)
);

AND2x6_ASAP7_75t_L g399 ( 
.A(n_331),
.B(n_318),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_399),
.B(n_401),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_323),
.C(n_315),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_337),
.B(n_283),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_402),
.B(n_355),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_338),
.A2(n_283),
.B1(n_318),
.B2(n_9),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_403),
.A2(n_355),
.B1(n_359),
.B2(n_329),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_406),
.B(n_418),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_381),
.A2(n_327),
.B1(n_328),
.B2(n_331),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_408),
.A2(n_417),
.B1(n_421),
.B2(n_340),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_387),
.B(n_362),
.Y(n_409)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_409),
.B(n_414),
.C(n_431),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_412),
.B(n_370),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_400),
.B(n_362),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_381),
.A2(n_349),
.B1(n_343),
.B2(n_367),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_371),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_419),
.A2(n_403),
.B1(n_375),
.B2(n_391),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_370),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_420),
.B(n_435),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_379),
.A2(n_366),
.B1(n_367),
.B2(n_345),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_369),
.B(n_356),
.Y(n_424)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_424),
.Y(n_446)
);

OAI32xp33_ASAP7_75t_L g426 ( 
.A1(n_379),
.A2(n_356),
.A3(n_347),
.B1(n_350),
.B2(n_365),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_426),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_394),
.A2(n_342),
.B(n_358),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_427),
.A2(n_412),
.B(n_424),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_389),
.B(n_364),
.Y(n_428)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_428),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_341),
.Y(n_432)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_432),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_378),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_405),
.B(n_372),
.C(n_374),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_436),
.B(n_438),
.C(n_439),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_405),
.B(n_386),
.C(n_380),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_410),
.B(n_370),
.C(n_394),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_440),
.A2(n_443),
.B(n_456),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_441),
.A2(n_442),
.B1(n_451),
.B2(n_452),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_417),
.A2(n_392),
.B1(n_395),
.B2(n_375),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_410),
.B(n_392),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_407),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_420),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_447),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_408),
.A2(n_421),
.B1(n_411),
.B2(n_407),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_404),
.B(n_383),
.C(n_397),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_453),
.B(n_413),
.C(n_430),
.Y(n_466)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_422),
.Y(n_454)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_454),
.Y(n_467)
);

BUFx12f_ASAP7_75t_L g455 ( 
.A(n_418),
.Y(n_455)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_455),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_434),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_457),
.B(n_458),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_434),
.B(n_393),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_428),
.B(n_399),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_459),
.B(n_460),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_411),
.A2(n_384),
.B1(n_351),
.B2(n_334),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_433),
.Y(n_461)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_461),
.Y(n_472)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_422),
.Y(n_462)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_462),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_466),
.B(n_469),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_459),
.B(n_415),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_468),
.B(n_416),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_432),
.C(n_427),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_477),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_438),
.B(n_415),
.C(n_433),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_473),
.B(n_476),
.C(n_485),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_453),
.B(n_439),
.C(n_440),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_445),
.B(n_413),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_440),
.B(n_430),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_479),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_452),
.B(n_429),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_480),
.B(n_419),
.C(n_334),
.Y(n_503)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_444),
.Y(n_481)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_481),
.Y(n_488)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_446),
.Y(n_482)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_482),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_447),
.A2(n_425),
.B(n_435),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_484),
.A2(n_441),
.B(n_423),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_448),
.B(n_429),
.C(n_423),
.Y(n_485)
);

A2O1A1O1Ixp25_ASAP7_75t_L g487 ( 
.A1(n_479),
.A2(n_447),
.B(n_437),
.C(n_460),
.D(n_449),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_487),
.A2(n_491),
.B(n_498),
.Y(n_505)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_465),
.Y(n_490)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_490),
.Y(n_511)
);

FAx1_ASAP7_75t_L g491 ( 
.A(n_470),
.B(n_464),
.CI(n_437),
.CON(n_491),
.SN(n_491)
);

FAx1_ASAP7_75t_SL g508 ( 
.A(n_491),
.B(n_469),
.CI(n_464),
.CON(n_508),
.SN(n_508)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_442),
.Y(n_492)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_492),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_484),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_495),
.B(n_496),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_450),
.C(n_416),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_471),
.B(n_455),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_497),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_498),
.A2(n_478),
.B(n_480),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_499),
.A2(n_501),
.B1(n_472),
.B2(n_336),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_455),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_500),
.B(n_466),
.Y(n_510)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_467),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_503),
.B(n_477),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_504),
.B(n_517),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_505),
.A2(n_513),
.B(n_493),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_493),
.B(n_474),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_507),
.B(n_486),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_508),
.B(n_509),
.Y(n_519)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_510),
.Y(n_528)
);

A2O1A1Ixp33_ASAP7_75t_L g513 ( 
.A1(n_487),
.A2(n_475),
.B(n_483),
.C(n_474),
.Y(n_513)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_515),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_494),
.B(n_463),
.C(n_365),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_516),
.B(n_518),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_494),
.B(n_463),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_491),
.A2(n_351),
.B1(n_350),
.B2(n_336),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_516),
.B(n_502),
.C(n_496),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_520),
.B(n_507),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_522),
.A2(n_508),
.B(n_8),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_523),
.B(n_524),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_504),
.B(n_486),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_512),
.A2(n_488),
.B1(n_489),
.B2(n_500),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_525),
.A2(n_527),
.B1(n_529),
.B2(n_513),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_514),
.A2(n_497),
.B1(n_503),
.B2(n_351),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g529 ( 
.A(n_510),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_528),
.A2(n_506),
.B(n_517),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_532),
.A2(n_535),
.B(n_537),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_533),
.B(n_534),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_521),
.B(n_509),
.C(n_511),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_520),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_536),
.A2(n_538),
.B(n_526),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_529),
.B(n_518),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_539),
.B(n_542),
.Y(n_545)
);

BUFx24_ASAP7_75t_SL g542 ( 
.A(n_531),
.Y(n_542)
);

AO21x1_ASAP7_75t_L g543 ( 
.A1(n_540),
.A2(n_519),
.B(n_521),
.Y(n_543)
);

AOI322xp5_ASAP7_75t_L g546 ( 
.A1(n_543),
.A2(n_530),
.A3(n_519),
.B1(n_508),
.B2(n_523),
.C1(n_524),
.C2(n_7),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_541),
.B(n_531),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_544),
.B(n_8),
.C(n_9),
.Y(n_547)
);

AO21x1_ASAP7_75t_SL g548 ( 
.A1(n_546),
.A2(n_547),
.B(n_9),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_548),
.A2(n_545),
.B1(n_10),
.B2(n_11),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_11),
.C(n_12),
.Y(n_551)
);

AO21x1_ASAP7_75t_L g552 ( 
.A1(n_551),
.A2(n_12),
.B(n_497),
.Y(n_552)
);


endmodule