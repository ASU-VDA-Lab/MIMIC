module fake_ariane_1827_n_37 (n_8, n_3, n_2, n_7, n_5, n_1, n_0, n_6, n_9, n_4, n_37);

input n_8;
input n_3;
input n_2;
input n_7;
input n_5;
input n_1;
input n_0;
input n_6;
input n_9;
input n_4;

output n_37;

wire n_24;
wire n_22;
wire n_13;
wire n_27;
wire n_20;
wire n_29;
wire n_17;
wire n_18;
wire n_32;
wire n_28;
wire n_11;
wire n_34;
wire n_26;
wire n_14;
wire n_36;
wire n_33;
wire n_19;
wire n_30;
wire n_31;
wire n_16;
wire n_12;
wire n_15;
wire n_21;
wire n_23;
wire n_35;
wire n_10;
wire n_25;

CKINVDCx5p33_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

CKINVDCx5p33_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx5p33_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_3),
.B(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_2),
.Y(n_21)
);

AND2x2_ASAP7_75t_SL g22 ( 
.A(n_18),
.B(n_2),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

OAI211xp5_ASAP7_75t_SL g24 ( 
.A1(n_21),
.A2(n_13),
.B(n_16),
.C(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

AOI21xp33_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_12),
.B(n_17),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_26),
.B1(n_17),
.B2(n_19),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_20),
.B1(n_23),
.B2(n_16),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g29 ( 
.A(n_27),
.B(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

AOI221xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_30),
.B1(n_24),
.B2(n_11),
.C(n_7),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_30),
.B1(n_11),
.B2(n_6),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_3),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_4),
.Y(n_34)
);

OAI221xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_11),
.B1(n_8),
.B2(n_9),
.C(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_34),
.B1(n_11),
.B2(n_8),
.Y(n_37)
);


endmodule