module fake_jpeg_25954_n_106 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_10),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_27),
.Y(n_42)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_21),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_32),
.B(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_30),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_23),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_31),
.A2(n_14),
.B1(n_15),
.B2(n_23),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_15),
.B1(n_14),
.B2(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_27),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_53),
.C(n_26),
.Y(n_65)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_39),
.B1(n_42),
.B2(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_12),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_17),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_28),
.B1(n_40),
.B2(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_22),
.B(n_16),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_61),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_69),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_64),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_56),
.B1(n_54),
.B2(n_48),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_76),
.C(n_58),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_71),
.B(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_58),
.B1(n_53),
.B2(n_65),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_45),
.B(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_77),
.B(n_79),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_46),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_50),
.C(n_51),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_87),
.B(n_67),
.Y(n_90)
);

AO221x1_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_59),
.B1(n_68),
.B2(n_64),
.C(n_3),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_67),
.B1(n_73),
.B2(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

A2O1A1O1Ixp25_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_76),
.B(n_70),
.C(n_71),
.D(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_93),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_81),
.B(n_86),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_92),
.C(n_81),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_80),
.C(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_7),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_SL g101 ( 
.A1(n_98),
.A2(n_94),
.B(n_97),
.C(n_8),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_100),
.B(n_6),
.Y(n_102)
);

OAI221xp5_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_16),
.B1(n_24),
.B2(n_18),
.C(n_13),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_102),
.C(n_0),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_6),
.A3(n_13),
.B1(n_2),
.B2(n_4),
.C1(n_0),
.C2(n_1),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_103),
.A2(n_104),
.B(n_1),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_16),
.Y(n_106)
);


endmodule