module fake_jpeg_6358_n_124 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_124);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_27),
.B(n_28),
.Y(n_53)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_29),
.A2(n_33),
.B1(n_20),
.B2(n_12),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_30),
.B(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_26),
.B(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_31),
.B(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_2),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

AOI21xp33_ASAP7_75t_L g35 ( 
.A1(n_23),
.A2(n_2),
.B(n_7),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_21),
.B(n_18),
.C(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_11),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_40),
.B(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_25),
.Y(n_39)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_15),
.A2(n_7),
.B(n_8),
.C(n_11),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_39),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

CKINVDCx12_ASAP7_75t_R g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_49),
.Y(n_69)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_50),
.B(n_55),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_27),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_56),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_27),
.A2(n_14),
.B1(n_13),
.B2(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_59),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_14),
.B1(n_13),
.B2(n_19),
.Y(n_55)
);

OR2x2_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_8),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_29),
.A2(n_19),
.B1(n_24),
.B2(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_28),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_24),
.C(n_36),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_28),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_76),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_46),
.Y(n_88)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_49),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_89),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_45),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_75),
.C(n_64),
.Y(n_92)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_41),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_66),
.B(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_95),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_68),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_78),
.B(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_99),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_78),
.B(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_83),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_100),
.B(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

A2O1A1O1Ixp25_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_89),
.B(n_99),
.C(n_92),
.D(n_67),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_67),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_76),
.B1(n_67),
.B2(n_86),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_108),
.B1(n_44),
.B2(n_60),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_91),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_102),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_70),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_109),
.B(n_101),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_117),
.A3(n_109),
.B1(n_105),
.B2(n_93),
.C1(n_58),
.C2(n_82),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_119),
.A2(n_114),
.B1(n_85),
.B2(n_101),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_121),
.C(n_120),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_41),
.Y(n_124)
);


endmodule