module fake_jpeg_7236_n_136 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_136);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_12),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_8),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_27),
.B(n_32),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_72),
.Y(n_90)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_78),
.Y(n_100)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_0),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_46),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_87),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_64),
.B1(n_54),
.B2(n_59),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_84),
.A2(n_94),
.B1(n_99),
.B2(n_11),
.Y(n_114)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

AO22x2_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_49),
.B1(n_41),
.B2(n_43),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_100),
.B1(n_90),
.B2(n_15),
.Y(n_111)
);

AO22x1_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_108)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_95),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_59),
.B1(n_65),
.B2(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_52),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_66),
.C(n_47),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_97),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_61),
.B1(n_60),
.B2(n_58),
.Y(n_99)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_48),
.B1(n_53),
.B2(n_50),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_104),
.B(n_107),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_118)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_45),
.B1(n_30),
.B2(n_31),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_5),
.B1(n_6),
.B2(n_10),
.Y(n_109)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_121),
.B1(n_116),
.B2(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_119),
.B1(n_115),
.B2(n_112),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_114),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_111),
.C(n_107),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_125),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_118),
.B1(n_101),
.B2(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_13),
.C(n_24),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_26),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_28),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_33),
.C(n_36),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_37),
.Y(n_136)
);


endmodule