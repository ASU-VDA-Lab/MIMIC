module fake_netlist_1_11553_n_666 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_666);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_666;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_649;
wire n_276;
wire n_526;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g75 ( .A(n_60), .Y(n_75) );
BUFx3_ASAP7_75t_L g76 ( .A(n_65), .Y(n_76) );
XOR2xp5_ASAP7_75t_L g77 ( .A(n_62), .B(n_5), .Y(n_77) );
HB1xp67_ASAP7_75t_L g78 ( .A(n_3), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_8), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_16), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_7), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_10), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_38), .Y(n_83) );
NOR2xp33_ASAP7_75t_L g84 ( .A(n_37), .B(n_46), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_64), .Y(n_85) );
NOR2xp67_ASAP7_75t_L g86 ( .A(n_58), .B(n_29), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_1), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_47), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_13), .Y(n_89) );
INVxp33_ASAP7_75t_L g90 ( .A(n_19), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_66), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_31), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_11), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_44), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_34), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_73), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_42), .Y(n_97) );
HB1xp67_ASAP7_75t_L g98 ( .A(n_14), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_1), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_41), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_33), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_54), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_22), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_18), .B(n_49), .Y(n_104) );
INVx2_ASAP7_75t_SL g105 ( .A(n_40), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_25), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_28), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_71), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_30), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_5), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_69), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_43), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_6), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_24), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_21), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_50), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_20), .Y(n_117) );
CKINVDCx14_ASAP7_75t_R g118 ( .A(n_70), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_48), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_57), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_75), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_119), .B(n_0), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_119), .B(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_120), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g125 ( .A(n_105), .B(n_2), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_113), .B(n_2), .Y(n_126) );
AND2x6_ASAP7_75t_L g127 ( .A(n_76), .B(n_35), .Y(n_127) );
INVx3_ASAP7_75t_L g128 ( .A(n_120), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_75), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_103), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_78), .Y(n_131) );
AND2x2_ASAP7_75t_SL g132 ( .A(n_98), .B(n_36), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_80), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_85), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_105), .B(n_3), .Y(n_135) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_83), .A2(n_39), .B(n_72), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_76), .Y(n_138) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_83), .A2(n_32), .B(n_68), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_90), .B(n_4), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_102), .B(n_4), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_88), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_87), .B(n_6), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_97), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_102), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_108), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_97), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_89), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_93), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_92), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g151 ( .A1(n_93), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_94), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_108), .Y(n_153) );
AOI22x1_ASAP7_75t_SL g154 ( .A1(n_82), .A2(n_12), .B1(n_15), .B2(n_17), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_111), .Y(n_155) );
INVx2_ASAP7_75t_SL g156 ( .A(n_111), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_118), .B(n_12), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_95), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_100), .Y(n_159) );
BUFx12f_ASAP7_75t_L g160 ( .A(n_96), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_101), .Y(n_161) );
NAND2xp33_ASAP7_75t_L g162 ( .A(n_127), .B(n_112), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_160), .Y(n_163) );
INVx2_ASAP7_75t_SL g164 ( .A(n_141), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_133), .B(n_91), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_133), .B(n_117), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_138), .Y(n_167) );
INVx2_ASAP7_75t_SL g168 ( .A(n_137), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_128), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_128), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_124), .A2(n_79), .B1(n_81), .B2(n_116), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_138), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_131), .B(n_99), .Y(n_174) );
NOR2x1p5_ASAP7_75t_L g175 ( .A(n_160), .B(n_99), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_138), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_134), .B(n_161), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_138), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_141), .B(n_86), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_134), .B(n_107), .Y(n_180) );
AND2x6_ASAP7_75t_L g181 ( .A(n_141), .B(n_84), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_138), .Y(n_182) );
BUFx4f_ASAP7_75t_L g183 ( .A(n_132), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_128), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_138), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_145), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
INVx1_ASAP7_75t_SL g188 ( .A(n_126), .Y(n_188) );
OR2x6_ASAP7_75t_L g189 ( .A(n_126), .B(n_77), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_145), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_142), .B(n_115), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_145), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_145), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_128), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_124), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_145), .Y(n_196) );
BUFx3_ASAP7_75t_L g197 ( .A(n_146), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_142), .B(n_161), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_148), .B(n_115), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_156), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_156), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_146), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_146), .Y(n_203) );
BUFx4f_ASAP7_75t_L g204 ( .A(n_132), .Y(n_204) );
INVx1_ASAP7_75t_SL g205 ( .A(n_157), .Y(n_205) );
INVx5_ASAP7_75t_L g206 ( .A(n_127), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_135), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_148), .B(n_114), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_150), .A2(n_110), .B1(n_112), .B2(n_114), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_146), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_121), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_146), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_121), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_150), .B(n_109), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_146), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_152), .B(n_109), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_152), .B(n_107), .Y(n_217) );
INVx4_ASAP7_75t_SL g218 ( .A(n_127), .Y(n_218) );
OR2x2_ASAP7_75t_L g219 ( .A(n_122), .B(n_77), .Y(n_219) );
INVx1_ASAP7_75t_SL g220 ( .A(n_157), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_207), .B(n_140), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_200), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_168), .B(n_123), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_191), .B(n_140), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_206), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_174), .B(n_159), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_191), .B(n_132), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_206), .B(n_218), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_206), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_169), .Y(n_230) );
INVx2_ASAP7_75t_SL g231 ( .A(n_206), .Y(n_231) );
INVxp67_ASAP7_75t_SL g232 ( .A(n_171), .Y(n_232) );
NOR2xp67_ASAP7_75t_L g233 ( .A(n_163), .B(n_143), .Y(n_233) );
OAI21xp5_ASAP7_75t_L g234 ( .A1(n_170), .A2(n_139), .B(n_136), .Y(n_234) );
NOR2xp33_ASAP7_75t_SL g235 ( .A(n_183), .B(n_130), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_208), .B(n_159), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_184), .Y(n_237) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_194), .A2(n_139), .B(n_136), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_208), .B(n_158), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_201), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_217), .B(n_158), .Y(n_241) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_205), .Y(n_242) );
BUFx3_ASAP7_75t_L g243 ( .A(n_181), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_217), .B(n_96), .Y(n_244) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_195), .A2(n_136), .B(n_139), .Y(n_245) );
INVxp67_ASAP7_75t_SL g246 ( .A(n_171), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_180), .B(n_106), .Y(n_247) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_220), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_199), .B(n_106), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_218), .B(n_153), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_214), .B(n_127), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_177), .B(n_147), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_183), .A2(n_127), .B1(n_125), .B2(n_144), .Y(n_253) );
NOR2x2_ASAP7_75t_L g254 ( .A(n_189), .B(n_154), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_173), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_171), .Y(n_256) );
AND2x4_ASAP7_75t_L g257 ( .A(n_179), .B(n_149), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_188), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_216), .B(n_127), .Y(n_259) );
AND2x6_ASAP7_75t_SL g260 ( .A(n_189), .B(n_154), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_211), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_173), .Y(n_262) );
NOR2xp67_ASAP7_75t_L g263 ( .A(n_163), .B(n_149), .Y(n_263) );
INVx2_ASAP7_75t_SL g264 ( .A(n_218), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_198), .B(n_147), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_204), .A2(n_127), .B1(n_147), .B2(n_144), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_165), .B(n_179), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_178), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_165), .B(n_144), .Y(n_269) );
NAND2x1_ASAP7_75t_L g270 ( .A(n_164), .B(n_136), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_213), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_164), .B(n_153), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_179), .B(n_166), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_219), .B(n_151), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_176), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_204), .B(n_153), .Y(n_276) );
INVx2_ASAP7_75t_SL g277 ( .A(n_181), .Y(n_277) );
BUFx4_ASAP7_75t_L g278 ( .A(n_189), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_178), .Y(n_279) );
AND2x6_ASAP7_75t_SL g280 ( .A(n_166), .B(n_104), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_209), .B(n_147), .Y(n_281) );
INVxp67_ASAP7_75t_L g282 ( .A(n_209), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_223), .B(n_162), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_258), .B(n_162), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_233), .B(n_175), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_270), .A2(n_139), .B(n_186), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_225), .Y(n_287) );
NOR2xp33_ASAP7_75t_R g288 ( .A(n_235), .B(n_181), .Y(n_288) );
INVx2_ASAP7_75t_SL g289 ( .A(n_242), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_257), .B(n_172), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_248), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_256), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_221), .B(n_172), .Y(n_293) );
CKINVDCx8_ASAP7_75t_R g294 ( .A(n_260), .Y(n_294) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_245), .A2(n_196), .B(n_187), .Y(n_295) );
AOI21x1_ASAP7_75t_L g296 ( .A1(n_251), .A2(n_196), .B(n_186), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_259), .A2(n_185), .B(n_187), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_L g298 ( .A1(n_281), .A2(n_144), .B(n_129), .C(n_155), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_252), .B(n_265), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_252), .B(n_181), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_256), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_256), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_265), .B(n_181), .Y(n_303) );
AOI22xp33_ASAP7_75t_SL g304 ( .A1(n_257), .A2(n_129), .B1(n_155), .B2(n_153), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_234), .A2(n_185), .B(n_192), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_257), .A2(n_153), .B1(n_212), .B2(n_176), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_274), .B(n_153), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g308 ( .A1(n_226), .A2(n_197), .B(n_212), .C(n_193), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_238), .A2(n_276), .B(n_272), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_243), .B(n_193), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_243), .B(n_197), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_225), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_274), .B(n_190), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_SL g314 ( .A1(n_276), .A2(n_210), .B(n_203), .C(n_192), .Y(n_314) );
INVx4_ASAP7_75t_L g315 ( .A(n_225), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_272), .A2(n_210), .B(n_203), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_227), .A2(n_190), .B1(n_182), .B2(n_215), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_230), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g319 ( .A1(n_282), .A2(n_182), .B1(n_202), .B2(n_215), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_267), .B(n_224), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_273), .B(n_215), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_225), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_244), .B(n_215), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_277), .B(n_202), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_254), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_222), .B(n_23), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_230), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_247), .B(n_202), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_254), .Y(n_329) );
AO31x2_ASAP7_75t_L g330 ( .A1(n_298), .A2(n_239), .A3(n_241), .B(n_236), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_299), .B(n_263), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_290), .A2(n_266), .B1(n_277), .B2(n_271), .Y(n_332) );
CKINVDCx14_ASAP7_75t_R g333 ( .A(n_325), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_286), .A2(n_228), .B(n_232), .Y(n_334) );
O2A1O1Ixp33_ASAP7_75t_SL g335 ( .A1(n_308), .A2(n_250), .B(n_269), .C(n_261), .Y(n_335) );
OAI21x1_ASAP7_75t_L g336 ( .A1(n_295), .A2(n_250), .B(n_275), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_309), .A2(n_228), .B(n_246), .Y(n_337) );
A2O1A1Ixp33_ASAP7_75t_L g338 ( .A1(n_283), .A2(n_240), .B(n_237), .C(n_253), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_289), .Y(n_339) );
AO31x2_ASAP7_75t_L g340 ( .A1(n_305), .A2(n_237), .A3(n_279), .B(n_268), .Y(n_340) );
OR2x6_ASAP7_75t_L g341 ( .A(n_329), .B(n_278), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_307), .Y(n_342) );
AO32x2_ASAP7_75t_L g343 ( .A1(n_317), .A2(n_280), .A3(n_264), .B1(n_231), .B2(n_167), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_293), .A2(n_249), .B(n_231), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_318), .Y(n_345) );
AOI21xp5_ASAP7_75t_SL g346 ( .A1(n_326), .A2(n_264), .B(n_229), .Y(n_346) );
AND2x6_ASAP7_75t_L g347 ( .A(n_326), .B(n_229), .Y(n_347) );
OAI21x1_ASAP7_75t_L g348 ( .A1(n_296), .A2(n_275), .B(n_279), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_291), .Y(n_349) );
AO31x2_ASAP7_75t_L g350 ( .A1(n_321), .A2(n_268), .A3(n_262), .B(n_255), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_320), .B(n_275), .Y(n_351) );
INVx2_ASAP7_75t_SL g352 ( .A(n_285), .Y(n_352) );
O2A1O1Ixp33_ASAP7_75t_L g353 ( .A1(n_300), .A2(n_303), .B(n_313), .C(n_284), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_290), .B(n_229), .Y(n_354) );
A2O1A1Ixp33_ASAP7_75t_L g355 ( .A1(n_328), .A2(n_262), .B(n_255), .C(n_202), .Y(n_355) );
OA21x2_ASAP7_75t_L g356 ( .A1(n_297), .A2(n_167), .B(n_229), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_306), .Y(n_357) );
NOR2x1_ASAP7_75t_R g358 ( .A(n_294), .B(n_167), .Y(n_358) );
OAI221xp5_ASAP7_75t_L g359 ( .A1(n_304), .A2(n_167), .B1(n_27), .B2(n_45), .C(n_51), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_331), .B(n_285), .Y(n_360) );
OA21x2_ASAP7_75t_L g361 ( .A1(n_348), .A2(n_323), .B(n_319), .Y(n_361) );
CKINVDCx8_ASAP7_75t_R g362 ( .A(n_341), .Y(n_362) );
AO31x2_ASAP7_75t_L g363 ( .A1(n_355), .A2(n_327), .A3(n_316), .B(n_302), .Y(n_363) );
AO21x2_ASAP7_75t_L g364 ( .A1(n_335), .A2(n_314), .B(n_324), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_341), .A2(n_288), .B1(n_301), .B2(n_292), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_347), .Y(n_366) );
A2O1A1Ixp33_ASAP7_75t_L g367 ( .A1(n_353), .A2(n_311), .B(n_310), .C(n_312), .Y(n_367) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_347), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_340), .Y(n_369) );
OAI21x1_ASAP7_75t_L g370 ( .A1(n_336), .A2(n_322), .B(n_312), .Y(n_370) );
INVx5_ASAP7_75t_L g371 ( .A(n_347), .Y(n_371) );
AOI21xp5_ASAP7_75t_L g372 ( .A1(n_334), .A2(n_322), .B(n_312), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_339), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_340), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_349), .Y(n_375) );
AOI222xp33_ASAP7_75t_L g376 ( .A1(n_342), .A2(n_315), .B1(n_322), .B2(n_287), .C1(n_55), .C2(n_56), .Y(n_376) );
BUFx8_ASAP7_75t_L g377 ( .A(n_352), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_337), .A2(n_287), .B(n_315), .Y(n_378) );
BUFx8_ASAP7_75t_L g379 ( .A(n_343), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_354), .B(n_287), .Y(n_380) );
CKINVDCx6p67_ASAP7_75t_R g381 ( .A(n_358), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_344), .A2(n_26), .B(n_52), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g383 ( .A1(n_332), .A2(n_53), .B1(n_59), .B2(n_61), .C(n_63), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_333), .A2(n_67), .B1(n_74), .B2(n_351), .Y(n_384) );
OA21x2_ASAP7_75t_L g385 ( .A1(n_338), .A2(n_357), .B(n_359), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_369), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_369), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_374), .B(n_330), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_374), .Y(n_389) );
AO21x2_ASAP7_75t_L g390 ( .A1(n_367), .A2(n_346), .B(n_330), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_370), .Y(n_391) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_370), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_385), .B(n_330), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_385), .B(n_343), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_361), .Y(n_395) );
AO21x2_ASAP7_75t_L g396 ( .A1(n_367), .A2(n_340), .B(n_345), .Y(n_396) );
OA21x2_ASAP7_75t_L g397 ( .A1(n_372), .A2(n_356), .B(n_343), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_375), .B(n_350), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_360), .A2(n_373), .B1(n_365), .B2(n_383), .C(n_384), .Y(n_399) );
INVx2_ASAP7_75t_SL g400 ( .A(n_371), .Y(n_400) );
OR2x2_ASAP7_75t_SL g401 ( .A(n_368), .B(n_356), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_363), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_371), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_361), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_378), .A2(n_350), .B(n_385), .Y(n_405) );
AO21x2_ASAP7_75t_L g406 ( .A1(n_364), .A2(n_350), .B(n_382), .Y(n_406) );
OA21x2_ASAP7_75t_L g407 ( .A1(n_380), .A2(n_361), .B(n_379), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_363), .Y(n_408) );
INVx3_ASAP7_75t_L g409 ( .A(n_371), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_363), .B(n_371), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_363), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_379), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_381), .A2(n_379), .B1(n_376), .B2(n_377), .Y(n_413) );
INVx2_ASAP7_75t_SL g414 ( .A(n_371), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_366), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_366), .B(n_368), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_364), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_368), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_366), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_418), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_388), .B(n_368), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_388), .B(n_364), .Y(n_422) );
AO21x2_ASAP7_75t_L g423 ( .A1(n_405), .A2(n_362), .B(n_381), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_413), .A2(n_362), .B1(n_377), .B2(n_399), .C(n_398), .Y(n_424) );
NOR2x1p5_ASAP7_75t_L g425 ( .A(n_403), .B(n_377), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_388), .B(n_393), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_393), .B(n_386), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_398), .B(n_393), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_386), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_387), .B(n_394), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_412), .B(n_419), .Y(n_431) );
INVxp67_ASAP7_75t_SL g432 ( .A(n_389), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_389), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_387), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_389), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_395), .Y(n_436) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_403), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_394), .B(n_412), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_410), .B(n_416), .Y(n_439) );
INVx3_ASAP7_75t_L g440 ( .A(n_392), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_394), .B(n_410), .Y(n_441) );
INVxp67_ASAP7_75t_SL g442 ( .A(n_395), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_395), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_403), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_400), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_404), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_410), .B(n_402), .Y(n_447) );
OAI211xp5_ASAP7_75t_L g448 ( .A1(n_413), .A2(n_399), .B(n_415), .C(n_419), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_402), .B(n_396), .Y(n_449) );
INVx3_ASAP7_75t_L g450 ( .A(n_392), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_400), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_404), .Y(n_452) );
INVx5_ASAP7_75t_L g453 ( .A(n_403), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_396), .B(n_411), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_396), .B(n_411), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_396), .B(n_411), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_404), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_391), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_401), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_401), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_407), .B(n_408), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_408), .B(n_390), .Y(n_462) );
INVx4_ASAP7_75t_L g463 ( .A(n_409), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_415), .B(n_416), .Y(n_464) );
BUFx2_ASAP7_75t_L g465 ( .A(n_407), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_400), .Y(n_466) );
INVx3_ASAP7_75t_L g467 ( .A(n_392), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_416), .B(n_408), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_429), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_424), .B(n_416), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_428), .B(n_407), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_429), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_426), .B(n_416), .Y(n_473) );
INVx3_ASAP7_75t_L g474 ( .A(n_463), .Y(n_474) );
INVx3_ASAP7_75t_L g475 ( .A(n_463), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_453), .B(n_414), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_426), .B(n_418), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_424), .A2(n_405), .B(n_414), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_434), .Y(n_479) );
AND4x1_ASAP7_75t_L g480 ( .A(n_425), .B(n_414), .C(n_409), .D(n_407), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_427), .B(n_409), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_438), .B(n_407), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_434), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_428), .B(n_409), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_438), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_446), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_447), .B(n_390), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_441), .B(n_390), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_427), .B(n_390), .Y(n_489) );
NOR2xp33_ASAP7_75t_R g490 ( .A(n_420), .B(n_392), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_421), .B(n_397), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_421), .B(n_397), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_441), .B(n_397), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_448), .B(n_397), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_447), .B(n_397), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_430), .B(n_406), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_431), .Y(n_497) );
INVxp67_ASAP7_75t_L g498 ( .A(n_445), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_430), .B(n_417), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_451), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_439), .B(n_417), .Y(n_501) );
AND2x2_ASAP7_75t_SL g502 ( .A(n_465), .B(n_392), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_448), .B(n_406), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_466), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_425), .A2(n_406), .B1(n_417), .B2(n_391), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_459), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_446), .Y(n_507) );
BUFx3_ASAP7_75t_L g508 ( .A(n_453), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_422), .B(n_406), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_422), .B(n_391), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_459), .B(n_392), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_439), .B(n_392), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_460), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_460), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_439), .B(n_449), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_449), .B(n_435), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_433), .B(n_435), .Y(n_517) );
NOR2xp33_ASAP7_75t_SL g518 ( .A(n_463), .B(n_453), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_432), .B(n_439), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_432), .B(n_433), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_468), .B(n_462), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_444), .B(n_437), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_436), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_468), .B(n_462), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_468), .B(n_455), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_486), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_525), .B(n_456), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_518), .B(n_453), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_485), .B(n_461), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_506), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_516), .B(n_461), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_471), .B(n_433), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_525), .B(n_455), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_524), .B(n_454), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_524), .B(n_454), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_486), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_510), .B(n_435), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_498), .Y(n_538) );
O2A1O1Ixp33_ASAP7_75t_SL g539 ( .A1(n_476), .A2(n_444), .B(n_464), .C(n_436), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_521), .B(n_456), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_469), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_507), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_476), .A2(n_423), .B(n_442), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_507), .Y(n_544) );
AND2x4_ASAP7_75t_L g545 ( .A(n_474), .B(n_465), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_474), .B(n_468), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_497), .B(n_464), .Y(n_547) );
AOI211xp5_ASAP7_75t_L g548 ( .A1(n_470), .A2(n_452), .B(n_443), .C(n_442), .Y(n_548) );
OAI222xp33_ASAP7_75t_L g549 ( .A1(n_482), .A2(n_463), .B1(n_453), .B2(n_443), .C1(n_452), .C2(n_457), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_521), .B(n_446), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_484), .B(n_453), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_472), .B(n_423), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_495), .B(n_457), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_495), .B(n_457), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_515), .B(n_458), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_479), .B(n_423), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_483), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_520), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_513), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_514), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_515), .B(n_458), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_493), .B(n_458), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_487), .B(n_423), .Y(n_563) );
OAI21xp33_ASAP7_75t_L g564 ( .A1(n_494), .A2(n_503), .B(n_509), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_500), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_487), .B(n_440), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_482), .B(n_440), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_504), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_523), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_499), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_496), .B(n_440), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_477), .B(n_453), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_491), .B(n_440), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_481), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_492), .B(n_450), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_530), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_538), .B(n_480), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_527), .B(n_512), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_527), .B(n_512), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_564), .B(n_494), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_559), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_533), .B(n_473), .Y(n_582) );
NAND2x1p5_ASAP7_75t_L g583 ( .A(n_528), .B(n_475), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_560), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_541), .Y(n_585) );
AND2x2_ASAP7_75t_SL g586 ( .A(n_545), .B(n_502), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_548), .B(n_490), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_531), .B(n_519), .Y(n_588) );
INVx2_ASAP7_75t_SL g589 ( .A(n_558), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_562), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_563), .A2(n_470), .B1(n_501), .B2(n_489), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_562), .Y(n_592) );
OAI332xp33_ASAP7_75t_L g593 ( .A1(n_547), .A2(n_488), .A3(n_511), .B1(n_517), .B2(n_478), .B3(n_490), .C1(n_502), .C2(n_505), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_574), .B(n_499), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_563), .A2(n_501), .B1(n_522), .B2(n_474), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_532), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_531), .B(n_475), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_565), .B(n_508), .Y(n_598) );
INVxp67_ASAP7_75t_L g599 ( .A(n_568), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_532), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_570), .B(n_475), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_529), .B(n_505), .Y(n_602) );
INVx3_ASAP7_75t_L g603 ( .A(n_545), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_558), .B(n_501), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_570), .B(n_508), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_533), .B(n_450), .Y(n_606) );
AND2x4_ASAP7_75t_L g607 ( .A(n_545), .B(n_450), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_529), .B(n_450), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_541), .Y(n_609) );
NAND4xp75_ASAP7_75t_L g610 ( .A(n_543), .B(n_467), .C(n_551), .D(n_572), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_588), .Y(n_611) );
OAI322xp33_ASAP7_75t_L g612 ( .A1(n_580), .A2(n_571), .A3(n_552), .B1(n_556), .B2(n_537), .C1(n_569), .C2(n_557), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_577), .A2(n_566), .B1(n_567), .B2(n_575), .Y(n_613) );
A2O1A1Ixp33_ASAP7_75t_L g614 ( .A1(n_586), .A2(n_546), .B(n_540), .C(n_534), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_585), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_592), .B(n_553), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_592), .B(n_553), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_602), .B(n_540), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_600), .B(n_554), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_602), .B(n_534), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_580), .B(n_535), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_609), .B(n_554), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_576), .Y(n_623) );
INVxp67_ASAP7_75t_L g624 ( .A(n_598), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_581), .Y(n_625) );
INVxp67_ASAP7_75t_L g626 ( .A(n_589), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_600), .B(n_535), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_591), .B(n_550), .Y(n_628) );
A2O1A1Ixp33_ASAP7_75t_L g629 ( .A1(n_603), .A2(n_546), .B(n_567), .C(n_550), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_578), .B(n_561), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_584), .Y(n_631) );
AOI21xp33_ASAP7_75t_L g632 ( .A1(n_599), .A2(n_557), .B(n_571), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_616), .Y(n_633) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_623), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_614), .A2(n_587), .B(n_539), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g636 ( .A1(n_626), .A2(n_583), .B(n_610), .Y(n_636) );
A2O1A1Ixp33_ASAP7_75t_SL g637 ( .A1(n_632), .A2(n_603), .B(n_605), .C(n_595), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_629), .B(n_583), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_622), .Y(n_639) );
OAI221xp5_ASAP7_75t_SL g640 ( .A1(n_613), .A2(n_597), .B1(n_601), .B2(n_608), .C(n_594), .Y(n_640) );
OAI21xp5_ASAP7_75t_L g641 ( .A1(n_632), .A2(n_549), .B(n_608), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_624), .A2(n_604), .B1(n_590), .B2(n_596), .C(n_537), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_628), .A2(n_606), .B1(n_575), .B2(n_573), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_612), .A2(n_593), .B(n_607), .Y(n_644) );
INVx1_ASAP7_75t_SL g645 ( .A(n_617), .Y(n_645) );
OAI211xp5_ASAP7_75t_L g646 ( .A1(n_637), .A2(n_621), .B(n_620), .C(n_618), .Y(n_646) );
NAND4xp25_ASAP7_75t_L g647 ( .A(n_644), .B(n_611), .C(n_627), .D(n_631), .Y(n_647) );
A2O1A1Ixp33_ASAP7_75t_L g648 ( .A1(n_635), .A2(n_619), .B(n_622), .C(n_625), .Y(n_648) );
O2A1O1Ixp5_ASAP7_75t_L g649 ( .A1(n_638), .A2(n_615), .B(n_607), .C(n_546), .Y(n_649) );
A2O1A1Ixp33_ASAP7_75t_L g650 ( .A1(n_636), .A2(n_630), .B(n_582), .C(n_579), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_633), .Y(n_651) );
AOI211xp5_ASAP7_75t_SL g652 ( .A1(n_640), .A2(n_593), .B(n_566), .C(n_573), .Y(n_652) );
OR3x2_ASAP7_75t_L g653 ( .A(n_647), .B(n_639), .C(n_641), .Y(n_653) );
NOR2xp67_ASAP7_75t_L g654 ( .A(n_646), .B(n_634), .Y(n_654) );
NOR3xp33_ASAP7_75t_L g655 ( .A(n_649), .B(n_642), .C(n_634), .Y(n_655) );
OAI211xp5_ASAP7_75t_L g656 ( .A1(n_648), .A2(n_643), .B(n_645), .C(n_561), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_654), .Y(n_657) );
NAND3xp33_ASAP7_75t_SL g658 ( .A(n_655), .B(n_652), .C(n_650), .Y(n_658) );
AND2x4_ASAP7_75t_L g659 ( .A(n_657), .B(n_651), .Y(n_659) );
AND3x4_ASAP7_75t_L g660 ( .A(n_658), .B(n_653), .C(n_656), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_659), .Y(n_661) );
OAI22x1_ASAP7_75t_L g662 ( .A1(n_661), .A2(n_660), .B1(n_526), .B2(n_536), .Y(n_662) );
AO221x1_ASAP7_75t_L g663 ( .A1(n_662), .A2(n_467), .B1(n_526), .B2(n_536), .C(n_542), .Y(n_663) );
XNOR2xp5_ASAP7_75t_L g664 ( .A(n_663), .B(n_555), .Y(n_664) );
OA22x2_ASAP7_75t_L g665 ( .A1(n_664), .A2(n_555), .B1(n_542), .B2(n_544), .Y(n_665) );
AOI211xp5_ASAP7_75t_L g666 ( .A1(n_665), .A2(n_467), .B(n_544), .C(n_661), .Y(n_666) );
endmodule