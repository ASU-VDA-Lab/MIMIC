module fake_jpeg_30981_n_47 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_4),
.B(n_1),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_21),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_15),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_22),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_0),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_19),
.A2(n_18),
.B1(n_15),
.B2(n_16),
.Y(n_23)
);

NOR2x1_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_17),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_28),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_24),
.B1(n_16),
.B2(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_21),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_12),
.B1(n_18),
.B2(n_11),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_24),
.C(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_29),
.C(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_14),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_27),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_27),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_12),
.C(n_13),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_39),
.Y(n_41)
);

BUFx24_ASAP7_75t_SL g42 ( 
.A(n_40),
.Y(n_42)
);

OAI321xp33_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_34),
.A3(n_37),
.B1(n_6),
.B2(n_8),
.C(n_9),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_3),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_5),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_41),
.Y(n_47)
);


endmodule