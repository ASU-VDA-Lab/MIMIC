module fake_netlist_6_3066_n_1803 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1803);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1803;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_1214;
wire n_835;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_SL g169 ( 
.A(n_148),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_128),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_3),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_26),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_167),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_75),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_50),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_9),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_31),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_124),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_7),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_76),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_21),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_110),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_31),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_59),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_64),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_26),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_57),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_55),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_27),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_139),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_83),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_93),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_134),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_155),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_15),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_45),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_89),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_140),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_73),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_107),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_37),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_60),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_37),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_143),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_118),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_56),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_40),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_56),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_126),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_52),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_17),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_101),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_27),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_111),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_109),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_51),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_106),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_52),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_55),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_35),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_17),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_72),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_34),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_135),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_0),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_141),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_87),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_123),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_133),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_138),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_51),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_144),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_164),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_129),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_130),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_145),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_9),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_131),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_20),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_156),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_115),
.Y(n_244)
);

BUFx2_ASAP7_75t_SL g245 ( 
.A(n_29),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_43),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_99),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_40),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_25),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_6),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_44),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_8),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_127),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_20),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_13),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_154),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_50),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_94),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_42),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_90),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_39),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_150),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_54),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_16),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_168),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_5),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_46),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_105),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_48),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_54),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_104),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_152),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_39),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_63),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_98),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_62),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_53),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_15),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_0),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_146),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_29),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_5),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_149),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_84),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_35),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_81),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_2),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_14),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_28),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_21),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_157),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_11),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_57),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_43),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_61),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_153),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_30),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_77),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_36),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_28),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_11),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_108),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_24),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_44),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_142),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_147),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_88),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_166),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_112),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_67),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_114),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_18),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_91),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_78),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_3),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_19),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_116),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_102),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_96),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_137),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_36),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_22),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_4),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_34),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_1),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_68),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_47),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_71),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_33),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_25),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_42),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_69),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_45),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_38),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_163),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_92),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_228),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_294),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_246),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_287),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_228),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_228),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_287),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_173),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_198),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_228),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_228),
.Y(n_347)
);

BUFx6f_ASAP7_75t_SL g348 ( 
.A(n_247),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_296),
.B(n_1),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_199),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_206),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_313),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_228),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_313),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_271),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_228),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_173),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_231),
.B(n_2),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_209),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_173),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_173),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_213),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_219),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_335),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_176),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_323),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_323),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_323),
.Y(n_368)
);

INVxp33_ASAP7_75t_SL g369 ( 
.A(n_176),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_335),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_229),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_R g372 ( 
.A(n_276),
.B(n_66),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_222),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_170),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_178),
.B(n_4),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_268),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_222),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_229),
.B(n_6),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_189),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_261),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_261),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_223),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_177),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_177),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_229),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_174),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_226),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_175),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_177),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_240),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_179),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_285),
.B(n_7),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_177),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_181),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_180),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_247),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_180),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_189),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_197),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_180),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_231),
.B(n_8),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_180),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_210),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_210),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_247),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_249),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_256),
.B(n_275),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_256),
.B(n_10),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_252),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_259),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_287),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_275),
.B(n_10),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_267),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_210),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_201),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_270),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_202),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_277),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_210),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_234),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_302),
.B(n_12),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_279),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_288),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_234),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_234),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_203),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_290),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_302),
.B(n_12),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_374),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_357),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_386),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_388),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_391),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_371),
.B(n_172),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_341),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_394),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_342),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_399),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_415),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_338),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_352),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_357),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_417),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_426),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_349),
.B(n_178),
.Y(n_445)
);

NAND3xp33_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_248),
.C(n_221),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_346),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_385),
.B(n_187),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_360),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_345),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_373),
.B(n_221),
.Y(n_451)
);

INVx6_ASAP7_75t_L g452 ( 
.A(n_344),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_345),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_378),
.B(n_192),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_350),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_350),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_351),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_351),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_337),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_359),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_359),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_347),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_362),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_360),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_361),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_353),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_361),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_354),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_337),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_369),
.B(n_211),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_R g471 ( 
.A(n_362),
.B(n_205),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_393),
.Y(n_472)
);

NAND3xp33_ASAP7_75t_L g473 ( 
.A(n_428),
.B(n_248),
.C(n_234),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_356),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_344),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_L g476 ( 
.A(n_363),
.B(n_266),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_363),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_382),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_348),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_393),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_365),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_395),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_356),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_382),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_387),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_366),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_366),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_395),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_376),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_376),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_383),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_407),
.B(n_169),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_387),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_384),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_389),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_355),
.B(n_262),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_367),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_369),
.B(n_211),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_397),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_400),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_402),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_364),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_377),
.B(n_171),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_390),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_367),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_403),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_390),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_440),
.Y(n_508)
);

INVx4_ASAP7_75t_SL g509 ( 
.A(n_452),
.Y(n_509)
);

OR2x6_ASAP7_75t_L g510 ( 
.A(n_481),
.B(n_340),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_471),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_489),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_489),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_452),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_446),
.A2(n_401),
.B1(n_412),
.B2(n_408),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_492),
.B(n_404),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_454),
.B(n_368),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_446),
.A2(n_358),
.B1(n_255),
.B2(n_334),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_489),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_434),
.B(n_414),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_448),
.B(n_406),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_473),
.A2(n_454),
.B1(n_255),
.B2(n_334),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_445),
.B(n_406),
.Y(n_523)
);

BUFx4f_ASAP7_75t_L g524 ( 
.A(n_452),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_445),
.B(n_409),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_459),
.Y(n_526)
);

OAI221xp5_ASAP7_75t_L g527 ( 
.A1(n_473),
.A2(n_392),
.B1(n_329),
.B2(n_339),
.C(n_171),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_437),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_437),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_454),
.B(n_419),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_475),
.B(n_380),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_454),
.B(n_310),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_486),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_479),
.B(n_310),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_490),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_452),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_452),
.B(n_420),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_429),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_435),
.Y(n_539)
);

NOR2x1p5_ASAP7_75t_L g540 ( 
.A(n_475),
.B(n_396),
.Y(n_540)
);

OR2x6_ASAP7_75t_L g541 ( 
.A(n_450),
.B(n_477),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_475),
.B(n_409),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_479),
.B(n_310),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_496),
.A2(n_413),
.B1(n_423),
.B2(n_422),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_451),
.B(n_381),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_437),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_476),
.B(n_410),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_490),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_504),
.B(n_410),
.Y(n_549)
);

BUFx4f_ASAP7_75t_L g550 ( 
.A(n_435),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_447),
.Y(n_551)
);

INVx4_ASAP7_75t_SL g552 ( 
.A(n_435),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_447),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_441),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_490),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_447),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_486),
.B(n_310),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_468),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_435),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_462),
.B(n_424),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_462),
.B(n_466),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_469),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_435),
.Y(n_563)
);

OR2x6_ASAP7_75t_L g564 ( 
.A(n_507),
.B(n_343),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_469),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_469),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_462),
.B(n_425),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_435),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_451),
.B(n_413),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_502),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_430),
.B(n_416),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_503),
.A2(n_182),
.B1(n_250),
.B2(n_300),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_486),
.Y(n_573)
);

CKINVDCx16_ASAP7_75t_R g574 ( 
.A(n_470),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_453),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_474),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_430),
.B(n_416),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_466),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_503),
.B(n_411),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_474),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_466),
.B(n_418),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_442),
.B(n_418),
.Y(n_582)
);

BUFx6f_ASAP7_75t_SL g583 ( 
.A(n_491),
.Y(n_583)
);

AND2x2_ASAP7_75t_SL g584 ( 
.A(n_470),
.B(n_266),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_483),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_483),
.A2(n_184),
.B1(n_214),
.B2(n_188),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_442),
.B(n_422),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_455),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_449),
.B(n_423),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_491),
.B(n_245),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_486),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_486),
.B(n_427),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_464),
.B(n_427),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_486),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_465),
.B(n_396),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_SL g596 ( 
.A(n_456),
.B(n_242),
.Y(n_596)
);

INVx6_ASAP7_75t_L g597 ( 
.A(n_487),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_431),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_498),
.A2(n_254),
.B1(n_264),
.B2(n_293),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_467),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_495),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_487),
.Y(n_602)
);

INVxp33_ASAP7_75t_L g603 ( 
.A(n_498),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_457),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_467),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_458),
.B(n_379),
.Y(n_606)
);

INVxp33_ASAP7_75t_L g607 ( 
.A(n_506),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_460),
.B(n_405),
.Y(n_608)
);

INVx5_ASAP7_75t_L g609 ( 
.A(n_487),
.Y(n_609)
);

OAI22xp33_ASAP7_75t_L g610 ( 
.A1(n_461),
.A2(n_251),
.B1(n_257),
.B2(n_263),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_487),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_472),
.B(n_405),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_463),
.B(n_398),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_478),
.B(n_344),
.Y(n_614)
);

NAND2x1p5_ASAP7_75t_L g615 ( 
.A(n_497),
.B(n_194),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_484),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_480),
.B(n_319),
.Y(n_617)
);

BUFx10_ASAP7_75t_L g618 ( 
.A(n_485),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_493),
.B(n_289),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_432),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_482),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_500),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_488),
.B(n_348),
.Y(n_623)
);

INVx6_ASAP7_75t_L g624 ( 
.A(n_487),
.Y(n_624)
);

INVx5_ASAP7_75t_L g625 ( 
.A(n_487),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_494),
.B(n_348),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_494),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_505),
.B(n_372),
.Y(n_628)
);

CKINVDCx8_ASAP7_75t_R g629 ( 
.A(n_433),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_499),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_499),
.B(n_320),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_505),
.B(n_195),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_501),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_501),
.B(n_208),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_505),
.A2(n_282),
.B1(n_273),
.B2(n_269),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_506),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_500),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_436),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_500),
.B(n_212),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_505),
.B(n_196),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_505),
.A2(n_224),
.B1(n_333),
.B2(n_216),
.Y(n_641)
);

BUFx10_ASAP7_75t_L g642 ( 
.A(n_438),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_505),
.B(n_497),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_497),
.A2(n_266),
.B1(n_235),
.B2(n_284),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_497),
.B(n_200),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_444),
.Y(n_646)
);

NAND3xp33_ASAP7_75t_L g647 ( 
.A(n_515),
.B(n_297),
.C(n_292),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_627),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_517),
.B(n_207),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_521),
.B(n_215),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_521),
.B(n_204),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_516),
.B(n_217),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_581),
.B(n_278),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_512),
.Y(n_654)
);

INVx8_ASAP7_75t_L g655 ( 
.A(n_541),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_508),
.B(n_439),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_510),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_630),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_512),
.Y(n_659)
);

NOR2xp67_ASAP7_75t_L g660 ( 
.A(n_511),
.B(n_443),
.Y(n_660)
);

AO22x1_ASAP7_75t_L g661 ( 
.A1(n_523),
.A2(n_312),
.B1(n_191),
.B2(n_190),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_523),
.B(n_281),
.C(n_299),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_601),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_629),
.Y(n_664)
);

NAND3xp33_ASAP7_75t_L g665 ( 
.A(n_515),
.B(n_321),
.C(n_331),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_584),
.B(n_268),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_569),
.B(n_370),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_579),
.B(n_375),
.Y(n_668)
);

NAND2x1p5_ASAP7_75t_L g669 ( 
.A(n_514),
.B(n_272),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_600),
.B(n_274),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_584),
.B(n_268),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_525),
.B(n_268),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_525),
.B(n_268),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_605),
.B(n_283),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_539),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_633),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_513),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_531),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_538),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_636),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_608),
.B(n_375),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_613),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_589),
.B(n_183),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_524),
.B(n_268),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_531),
.B(n_291),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_621),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_519),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_614),
.B(n_289),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_599),
.A2(n_266),
.B1(n_263),
.B2(n_325),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_519),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_530),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_547),
.A2(n_225),
.B1(n_332),
.B2(n_328),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_593),
.B(n_571),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_638),
.B(n_305),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_599),
.B(n_308),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_571),
.B(n_183),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_526),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_547),
.A2(n_218),
.B1(n_326),
.B2(n_318),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_545),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_577),
.B(n_185),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_545),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_535),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_548),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_615),
.B(n_336),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_548),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_549),
.B(n_330),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_582),
.B(n_185),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_619),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_582),
.B(n_220),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_587),
.B(n_514),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_587),
.B(n_227),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_560),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_592),
.A2(n_265),
.B1(n_230),
.B2(n_232),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_518),
.A2(n_522),
.B1(n_572),
.B2(n_527),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_579),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_615),
.B(n_233),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_567),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_540),
.B(n_186),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_536),
.B(n_520),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_542),
.B(n_236),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_595),
.B(n_237),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_595),
.B(n_238),
.Y(n_722)
);

INVxp67_ASAP7_75t_SL g723 ( 
.A(n_539),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_607),
.B(n_289),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_555),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_607),
.B(n_239),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_SL g727 ( 
.A(n_618),
.B(n_242),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_555),
.Y(n_728)
);

BUFx8_ASAP7_75t_L g729 ( 
.A(n_583),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_603),
.B(n_186),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_L g731 ( 
.A(n_537),
.B(n_634),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_590),
.B(n_193),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_631),
.B(n_241),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_631),
.B(n_639),
.Y(n_734)
);

OR2x6_ASAP7_75t_L g735 ( 
.A(n_575),
.B(n_251),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_562),
.Y(n_736)
);

INVx5_ASAP7_75t_L g737 ( 
.A(n_539),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_562),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_603),
.B(n_193),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_544),
.B(n_243),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_518),
.A2(n_325),
.B1(n_257),
.B2(n_190),
.Y(n_741)
);

AO221x1_ASAP7_75t_L g742 ( 
.A1(n_610),
.A2(n_262),
.B1(n_330),
.B2(n_304),
.C(n_312),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_SL g743 ( 
.A(n_618),
.B(n_262),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_539),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_565),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_565),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_617),
.B(n_244),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_579),
.B(n_307),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_522),
.A2(n_191),
.B1(n_330),
.B2(n_304),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_592),
.B(n_253),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_572),
.A2(n_304),
.B1(n_324),
.B2(n_322),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_566),
.B(n_306),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_606),
.B(n_327),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_628),
.A2(n_258),
.B1(n_317),
.B2(n_260),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_612),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_534),
.A2(n_280),
.B1(n_286),
.B2(n_295),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_563),
.B(n_298),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_566),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_590),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_568),
.B(n_314),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_534),
.B(n_309),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_576),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_543),
.B(n_311),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_576),
.B(n_311),
.Y(n_764)
);

AND2x2_ASAP7_75t_SL g765 ( 
.A(n_574),
.B(n_85),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_580),
.B(n_307),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_644),
.A2(n_315),
.B1(n_303),
.B2(n_301),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_L g768 ( 
.A(n_543),
.B(n_316),
.C(n_16),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_642),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_580),
.B(n_80),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_585),
.B(n_79),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_585),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_620),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_561),
.B(n_82),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_590),
.Y(n_775)
);

NOR2xp67_ASAP7_75t_L g776 ( 
.A(n_588),
.B(n_165),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_533),
.B(n_74),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_586),
.A2(n_13),
.B1(n_18),
.B2(n_19),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_532),
.A2(n_86),
.B1(n_161),
.B2(n_158),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_532),
.A2(n_70),
.B1(n_151),
.B2(n_136),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_528),
.B(n_65),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_622),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_642),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_611),
.B(n_594),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_510),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_637),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_611),
.B(n_58),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_550),
.A2(n_553),
.B(n_529),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_510),
.B(n_22),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_693),
.B(n_556),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_693),
.B(n_551),
.Y(n_791)
);

AO32x1_ASAP7_75t_L g792 ( 
.A1(n_697),
.A2(n_637),
.A3(n_578),
.B1(n_546),
.B2(n_591),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_664),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_651),
.B(n_753),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_651),
.B(n_570),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_719),
.A2(n_550),
.B(n_573),
.Y(n_796)
);

NOR3xp33_ASAP7_75t_L g797 ( 
.A(n_682),
.B(n_610),
.C(n_604),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_696),
.B(n_598),
.Y(n_798)
);

O2A1O1Ixp5_ASAP7_75t_L g799 ( 
.A1(n_672),
.A2(n_632),
.B(n_640),
.C(n_557),
.Y(n_799)
);

O2A1O1Ixp5_ASAP7_75t_L g800 ( 
.A1(n_672),
.A2(n_632),
.B(n_640),
.C(n_557),
.Y(n_800)
);

OR2x6_ASAP7_75t_SL g801 ( 
.A(n_679),
.B(n_596),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_724),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_788),
.A2(n_573),
.B(n_591),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_686),
.Y(n_804)
);

AOI21x1_ASAP7_75t_L g805 ( 
.A1(n_673),
.A2(n_643),
.B(n_645),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_R g806 ( 
.A(n_773),
.B(n_783),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_696),
.B(n_554),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_656),
.Y(n_808)
);

A2O1A1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_700),
.A2(n_623),
.B(n_626),
.C(n_586),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_675),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_SL g811 ( 
.A(n_741),
.B(n_558),
.C(n_616),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_785),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_734),
.B(n_559),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_700),
.B(n_564),
.C(n_646),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_677),
.Y(n_815)
);

O2A1O1Ixp33_ASAP7_75t_SL g816 ( 
.A1(n_673),
.A2(n_645),
.B(n_623),
.C(n_626),
.Y(n_816)
);

NAND2x1p5_ASAP7_75t_L g817 ( 
.A(n_675),
.B(n_559),
.Y(n_817)
);

AO21x1_ASAP7_75t_L g818 ( 
.A1(n_666),
.A2(n_644),
.B(n_641),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_707),
.A2(n_541),
.B1(n_635),
.B2(n_641),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_731),
.A2(n_559),
.B(n_602),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_706),
.B(n_541),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_666),
.A2(n_635),
.B(n_625),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_675),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_707),
.B(n_564),
.Y(n_824)
);

O2A1O1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_650),
.A2(n_564),
.B(n_583),
.C(n_30),
.Y(n_825)
);

AOI21x1_ASAP7_75t_L g826 ( 
.A1(n_684),
.A2(n_552),
.B(n_624),
.Y(n_826)
);

O2A1O1Ixp33_ASAP7_75t_SL g827 ( 
.A1(n_774),
.A2(n_552),
.B(n_509),
.C(n_597),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_710),
.A2(n_559),
.B(n_602),
.Y(n_828)
);

INVx3_ASAP7_75t_SL g829 ( 
.A(n_655),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_675),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_784),
.A2(n_602),
.B(n_609),
.Y(n_831)
);

NOR2xp67_ASAP7_75t_L g832 ( 
.A(n_708),
.B(n_730),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_744),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_737),
.A2(n_602),
.B(n_609),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_737),
.A2(n_609),
.B(n_625),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_691),
.B(n_509),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_664),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_737),
.A2(n_625),
.B(n_552),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_653),
.A2(n_23),
.B(n_24),
.C(n_32),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_688),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_648),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_712),
.B(n_624),
.Y(n_842)
);

BUFx12f_ASAP7_75t_L g843 ( 
.A(n_729),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_717),
.B(n_624),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_737),
.A2(n_597),
.B(n_100),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_714),
.B(n_597),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_669),
.A2(n_97),
.B(n_132),
.Y(n_847)
);

OAI21xp5_ASAP7_75t_L g848 ( 
.A1(n_671),
.A2(n_162),
.B(n_125),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_714),
.B(n_121),
.Y(n_849)
);

BUFx12f_ASAP7_75t_L g850 ( 
.A(n_729),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_653),
.A2(n_122),
.B1(n_120),
.B2(n_119),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_SL g852 ( 
.A(n_769),
.B(n_117),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_669),
.A2(n_113),
.B(n_103),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_667),
.Y(n_854)
);

AO21x1_ASAP7_75t_L g855 ( 
.A1(n_774),
.A2(n_23),
.B(n_32),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_755),
.B(n_33),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_744),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_709),
.B(n_38),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_681),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_652),
.B(n_41),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_711),
.A2(n_41),
.B1(n_46),
.B2(n_47),
.Y(n_861)
);

O2A1O1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_695),
.A2(n_750),
.B(n_766),
.C(n_764),
.Y(n_862)
);

NOR3xp33_ASAP7_75t_L g863 ( 
.A(n_740),
.B(n_48),
.C(n_49),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_683),
.B(n_49),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_683),
.B(n_53),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_723),
.A2(n_757),
.B(n_760),
.Y(n_866)
);

AND2x6_ASAP7_75t_L g867 ( 
.A(n_779),
.B(n_780),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_658),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_676),
.B(n_680),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_744),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_733),
.B(n_747),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_762),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_702),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_762),
.A2(n_772),
.B(n_728),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_744),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_715),
.Y(n_876)
);

AO22x1_ASAP7_75t_L g877 ( 
.A1(n_662),
.A2(n_789),
.B1(n_761),
.B2(n_763),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_765),
.B(n_730),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_739),
.B(n_689),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_739),
.A2(n_778),
.B1(n_722),
.B2(n_721),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_772),
.B(n_703),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_769),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_703),
.B(n_728),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_726),
.A2(n_777),
.B(n_787),
.Y(n_884)
);

INVx4_ASAP7_75t_L g885 ( 
.A(n_655),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_699),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_663),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_663),
.Y(n_888)
);

AND2x2_ASAP7_75t_SL g889 ( 
.A(n_765),
.B(n_689),
.Y(n_889)
);

OR2x6_ASAP7_75t_L g890 ( 
.A(n_655),
.B(n_657),
.Y(n_890)
);

BUFx4f_ASAP7_75t_L g891 ( 
.A(n_694),
.Y(n_891)
);

NOR3xp33_ASAP7_75t_L g892 ( 
.A(n_740),
.B(n_661),
.C(n_748),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_752),
.A2(n_782),
.B(n_786),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_668),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_761),
.B(n_763),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_735),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_736),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_752),
.A2(n_750),
.B(n_758),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_647),
.A2(n_665),
.B(n_748),
.C(n_649),
.Y(n_899)
);

O2A1O1Ixp5_ASAP7_75t_L g900 ( 
.A1(n_704),
.A2(n_716),
.B(n_766),
.C(n_764),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_701),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_695),
.A2(n_704),
.B(n_716),
.C(n_670),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_738),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_745),
.A2(n_746),
.B(n_654),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_674),
.B(n_649),
.Y(n_905)
);

NOR2x1_ASAP7_75t_R g906 ( 
.A(n_732),
.B(n_718),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_741),
.B(n_678),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_659),
.B(n_725),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_720),
.B(n_727),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_687),
.A2(n_705),
.B(n_690),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_781),
.A2(n_770),
.B(n_771),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_778),
.A2(n_685),
.B1(n_768),
.B2(n_742),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_685),
.B(n_759),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_781),
.A2(n_770),
.B(n_771),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_692),
.B(n_698),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_720),
.B(n_713),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_775),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_776),
.B(n_754),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_743),
.B(n_732),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_756),
.A2(n_718),
.B(n_749),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_749),
.B(n_767),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_789),
.A2(n_751),
.B(n_660),
.C(n_694),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_694),
.A2(n_751),
.B(n_735),
.Y(n_923)
);

OAI321xp33_ASAP7_75t_L g924 ( 
.A1(n_735),
.A2(n_651),
.A3(n_599),
.B1(n_700),
.B2(n_707),
.C(n_696),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_719),
.A2(n_524),
.B(n_550),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_651),
.B(n_693),
.Y(n_926)
);

INVx3_ASAP7_75t_SL g927 ( 
.A(n_679),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_693),
.B(n_734),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_719),
.A2(n_524),
.B(n_550),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_686),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_693),
.B(n_734),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_693),
.A2(n_651),
.B1(n_734),
.B2(n_700),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_693),
.B(n_734),
.Y(n_933)
);

OAI21xp33_ASAP7_75t_L g934 ( 
.A1(n_651),
.A2(n_445),
.B(n_696),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_651),
.B(n_693),
.Y(n_935)
);

BUFx4f_ASAP7_75t_L g936 ( 
.A(n_655),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_656),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_651),
.A2(n_693),
.B(n_650),
.C(n_671),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_SL g939 ( 
.A1(n_672),
.A2(n_673),
.B(n_774),
.C(n_666),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_656),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_719),
.A2(n_524),
.B(n_550),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_693),
.B(n_734),
.Y(n_942)
);

NAND2xp33_ASAP7_75t_L g943 ( 
.A(n_710),
.B(n_650),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_693),
.B(n_734),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_672),
.A2(n_673),
.B(n_693),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_651),
.B(n_693),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_651),
.A2(n_693),
.B(n_700),
.C(n_696),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_656),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_651),
.B(n_508),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_693),
.B(n_734),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_693),
.B(n_734),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_693),
.B(n_734),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_651),
.B(n_693),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_693),
.A2(n_651),
.B1(n_700),
.B2(n_696),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_693),
.B(n_734),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_651),
.B(n_693),
.Y(n_956)
);

AO32x1_ASAP7_75t_L g957 ( 
.A1(n_697),
.A2(n_231),
.A3(n_275),
.B1(n_256),
.B2(n_686),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_651),
.B(n_508),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_719),
.A2(n_524),
.B(n_550),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_693),
.B(n_734),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_651),
.B(n_693),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_949),
.B(n_958),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_926),
.B(n_935),
.Y(n_963)
);

BUFx12f_ASAP7_75t_L g964 ( 
.A(n_843),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_946),
.B(n_953),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_954),
.B(n_932),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_854),
.Y(n_967)
);

AOI221x1_ASAP7_75t_L g968 ( 
.A1(n_947),
.A2(n_934),
.B1(n_956),
.B2(n_961),
.C(n_892),
.Y(n_968)
);

AO21x2_ASAP7_75t_L g969 ( 
.A1(n_945),
.A2(n_895),
.B(n_803),
.Y(n_969)
);

NAND2x1p5_ASAP7_75t_L g970 ( 
.A(n_823),
.B(n_833),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_928),
.B(n_931),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_939),
.A2(n_943),
.B(n_813),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_798),
.B(n_808),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_938),
.A2(n_924),
.B(n_879),
.C(n_952),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_813),
.A2(n_914),
.B(n_911),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_928),
.B(n_931),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_933),
.B(n_942),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_805),
.A2(n_828),
.B(n_826),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_804),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_948),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_940),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_933),
.B(n_942),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_950),
.A2(n_952),
.B(n_951),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_823),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_866),
.A2(n_831),
.B(n_898),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_955),
.B(n_944),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_881),
.A2(n_883),
.B(n_796),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_841),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_881),
.A2(n_883),
.B(n_884),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_955),
.B(n_960),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_904),
.A2(n_910),
.B(n_817),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_832),
.B(n_889),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_823),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_849),
.A2(n_880),
.B(n_846),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_794),
.B(n_859),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_937),
.Y(n_996)
);

OR2x2_ASAP7_75t_L g997 ( 
.A(n_795),
.B(n_894),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_846),
.A2(n_799),
.B(n_800),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_871),
.A2(n_900),
.B(n_862),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_807),
.B(n_878),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_905),
.A2(n_959),
.B(n_941),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_833),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_925),
.A2(n_929),
.B(n_791),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_SL g1004 ( 
.A1(n_855),
.A2(n_848),
.B(n_902),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_790),
.A2(n_791),
.B(n_916),
.Y(n_1005)
);

AO21x2_ASAP7_75t_L g1006 ( 
.A1(n_790),
.A2(n_816),
.B(n_809),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_869),
.B(n_864),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_921),
.A2(n_915),
.B(n_822),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_869),
.B(n_864),
.Y(n_1009)
);

NAND2x1p5_ASAP7_75t_L g1010 ( 
.A(n_833),
.B(n_857),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_865),
.A2(n_842),
.B(n_844),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_865),
.B(n_877),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_920),
.A2(n_923),
.B(n_909),
.C(n_824),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_873),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_837),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_802),
.B(n_868),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_834),
.A2(n_872),
.B(n_838),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_930),
.B(n_907),
.Y(n_1018)
);

AOI21xp33_ASAP7_75t_L g1019 ( 
.A1(n_819),
.A2(n_840),
.B(n_918),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_842),
.A2(n_899),
.B(n_836),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_818),
.A2(n_792),
.B(n_908),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_860),
.A2(n_867),
.B(n_856),
.Y(n_1022)
);

AOI21x1_ASAP7_75t_L g1023 ( 
.A1(n_903),
.A2(n_860),
.B(n_888),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_792),
.A2(n_827),
.B(n_922),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_867),
.A2(n_856),
.B(n_912),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_897),
.Y(n_1026)
);

AOI221x1_ASAP7_75t_L g1027 ( 
.A1(n_863),
.A2(n_797),
.B1(n_861),
.B2(n_839),
.C(n_811),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_792),
.A2(n_887),
.B(n_858),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_814),
.B(n_919),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_857),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_887),
.B(n_897),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_821),
.B(n_867),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_847),
.A2(n_853),
.B(n_845),
.Y(n_1033)
);

AOI21x1_ASAP7_75t_L g1034 ( 
.A1(n_835),
.A2(n_917),
.B(n_876),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_793),
.B(n_901),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_927),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_867),
.B(n_886),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_810),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_867),
.B(n_913),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_851),
.A2(n_875),
.B(n_870),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_896),
.B(n_812),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_913),
.B(n_801),
.Y(n_1042)
);

NOR2x1_ASAP7_75t_SL g1043 ( 
.A(n_857),
.B(n_882),
.Y(n_1043)
);

O2A1O1Ixp5_ASAP7_75t_L g1044 ( 
.A1(n_830),
.A2(n_875),
.B(n_891),
.C(n_957),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_SL g1045 ( 
.A1(n_825),
.A2(n_885),
.B(n_882),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_891),
.A2(n_852),
.B(n_936),
.C(n_906),
.Y(n_1046)
);

AO31x2_ASAP7_75t_L g1047 ( 
.A1(n_957),
.A2(n_885),
.A3(n_890),
.B(n_936),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_957),
.A2(n_890),
.B(n_829),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_890),
.A2(n_806),
.B(n_850),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_926),
.B(n_935),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_SL g1051 ( 
.A(n_926),
.B(n_946),
.C(n_935),
.Y(n_1051)
);

NAND2x1_ASAP7_75t_L g1052 ( 
.A(n_823),
.B(n_833),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_820),
.A2(n_893),
.B(n_874),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_937),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_927),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_854),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_926),
.B(n_935),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_926),
.B(n_935),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_926),
.B(n_935),
.Y(n_1059)
);

AO31x2_ASAP7_75t_L g1060 ( 
.A1(n_947),
.A2(n_954),
.A3(n_880),
.B(n_818),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_926),
.B(n_935),
.Y(n_1061)
);

AO31x2_ASAP7_75t_L g1062 ( 
.A1(n_947),
.A2(n_954),
.A3(n_880),
.B(n_818),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_926),
.B(n_935),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_854),
.Y(n_1064)
);

O2A1O1Ixp5_ASAP7_75t_L g1065 ( 
.A1(n_954),
.A2(n_947),
.B(n_895),
.C(n_961),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_926),
.B(n_935),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_947),
.A2(n_954),
.B(n_932),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_939),
.A2(n_945),
.B(n_524),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_926),
.B(n_935),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_823),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_926),
.A2(n_946),
.B1(n_953),
.B2(n_935),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_815),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_940),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_947),
.A2(n_954),
.B(n_926),
.C(n_946),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_926),
.B(n_935),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_939),
.A2(n_945),
.B(n_524),
.Y(n_1076)
);

NAND2xp33_ASAP7_75t_SL g1077 ( 
.A(n_806),
.B(n_879),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_885),
.B(n_913),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_949),
.B(n_958),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_939),
.A2(n_945),
.B(n_524),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_947),
.A2(n_954),
.B(n_932),
.Y(n_1081)
);

AOI221xp5_ASAP7_75t_SL g1082 ( 
.A1(n_954),
.A2(n_926),
.B1(n_953),
.B2(n_946),
.C(n_935),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_947),
.A2(n_954),
.B(n_932),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_947),
.A2(n_954),
.B(n_932),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_939),
.A2(n_945),
.B(n_524),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_949),
.B(n_958),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_926),
.B(n_935),
.Y(n_1087)
);

OA21x2_ASAP7_75t_L g1088 ( 
.A1(n_945),
.A2(n_849),
.B(n_846),
.Y(n_1088)
);

OR2x6_ASAP7_75t_SL g1089 ( 
.A(n_954),
.B(n_679),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_926),
.B(n_935),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_926),
.A2(n_946),
.B(n_953),
.C(n_935),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_947),
.A2(n_954),
.B(n_932),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_947),
.A2(n_954),
.B(n_932),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_926),
.B(n_935),
.Y(n_1094)
);

AOI21xp33_ASAP7_75t_L g1095 ( 
.A1(n_926),
.A2(n_961),
.B(n_946),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_947),
.A2(n_935),
.B1(n_946),
.B2(n_926),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_947),
.A2(n_954),
.B(n_932),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_939),
.A2(n_945),
.B(n_524),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_926),
.B(n_935),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_939),
.A2(n_945),
.B(n_524),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_947),
.A2(n_935),
.B1(n_946),
.B2(n_926),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_926),
.B(n_935),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_926),
.B(n_935),
.Y(n_1103)
);

INVxp67_ASAP7_75t_L g1104 ( 
.A(n_948),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_926),
.B(n_935),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_954),
.B(n_932),
.Y(n_1106)
);

INVx5_ASAP7_75t_L g1107 ( 
.A(n_823),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_823),
.Y(n_1108)
);

AND2x6_ASAP7_75t_L g1109 ( 
.A(n_1002),
.B(n_1108),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1063),
.A2(n_1066),
.B1(n_1051),
.B2(n_1095),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_971),
.B(n_976),
.Y(n_1111)
);

OAI21xp33_ASAP7_75t_L g1112 ( 
.A1(n_1071),
.A2(n_965),
.B(n_963),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_979),
.Y(n_1113)
);

OAI21xp33_ASAP7_75t_L g1114 ( 
.A1(n_1050),
.A2(n_1058),
.B(n_1057),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_1055),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_988),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_962),
.B(n_1079),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_997),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_1077),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_964),
.Y(n_1120)
);

NAND2x1p5_ASAP7_75t_L g1121 ( 
.A(n_1107),
.B(n_1002),
.Y(n_1121)
);

NOR2x1_ASAP7_75t_L g1122 ( 
.A(n_995),
.B(n_1035),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_978),
.A2(n_987),
.B(n_991),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1086),
.B(n_973),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_977),
.B(n_982),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_967),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_1056),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_1036),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1059),
.B(n_1061),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1069),
.B(n_1075),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1087),
.B(n_1090),
.Y(n_1131)
);

CKINVDCx8_ASAP7_75t_R g1132 ( 
.A(n_1064),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_981),
.Y(n_1133)
);

INVx3_ASAP7_75t_SL g1134 ( 
.A(n_1015),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1094),
.B(n_1099),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_1041),
.Y(n_1136)
);

BUFx2_ASAP7_75t_SL g1137 ( 
.A(n_1078),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_981),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1000),
.B(n_1102),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_980),
.Y(n_1140)
);

NOR3xp33_ASAP7_75t_L g1141 ( 
.A(n_1051),
.B(n_1091),
.C(n_1105),
.Y(n_1141)
);

CKINVDCx11_ASAP7_75t_R g1142 ( 
.A(n_1089),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_980),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_1107),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_1103),
.B(n_1073),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1082),
.B(n_983),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_999),
.A2(n_1005),
.B(n_975),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1042),
.B(n_1104),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1005),
.A2(n_975),
.B(n_1076),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_1104),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_1096),
.B(n_1101),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1002),
.Y(n_1152)
);

INVx3_ASAP7_75t_SL g1153 ( 
.A(n_1078),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1029),
.B(n_1018),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_996),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1014),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1067),
.A2(n_1084),
.B1(n_1097),
.B2(n_1083),
.Y(n_1157)
);

NAND2x1_ASAP7_75t_L g1158 ( 
.A(n_1108),
.B(n_1038),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1046),
.B(n_1054),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_992),
.B(n_986),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1032),
.B(n_990),
.Y(n_1161)
);

AND2x2_ASAP7_75t_SL g1162 ( 
.A(n_1012),
.B(n_1039),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_966),
.B(n_1106),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1043),
.B(n_1037),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1072),
.Y(n_1165)
);

INVx4_ASAP7_75t_L g1166 ( 
.A(n_1107),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1081),
.A2(n_1092),
.B1(n_1093),
.B2(n_1074),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_1049),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1016),
.B(n_1007),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_1107),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1068),
.A2(n_1100),
.B(n_1098),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_983),
.B(n_1009),
.Y(n_1172)
);

CKINVDCx16_ASAP7_75t_R g1173 ( 
.A(n_1025),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_1052),
.Y(n_1174)
);

NAND3xp33_ASAP7_75t_L g1175 ( 
.A(n_1013),
.B(n_1074),
.C(n_968),
.Y(n_1175)
);

BUFx12f_ASAP7_75t_L g1176 ( 
.A(n_970),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1026),
.Y(n_1177)
);

BUFx12f_ASAP7_75t_L g1178 ( 
.A(n_970),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1068),
.A2(n_1100),
.B(n_1076),
.Y(n_1179)
);

NAND2x1p5_ASAP7_75t_L g1180 ( 
.A(n_984),
.B(n_993),
.Y(n_1180)
);

AO21x2_ASAP7_75t_L g1181 ( 
.A1(n_1004),
.A2(n_998),
.B(n_994),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_974),
.B(n_1008),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1031),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1022),
.B(n_1019),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_1060),
.B(n_1062),
.Y(n_1185)
);

INVx1_ASAP7_75t_SL g1186 ( 
.A(n_993),
.Y(n_1186)
);

INVxp67_ASAP7_75t_L g1187 ( 
.A(n_1049),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1065),
.B(n_1060),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1065),
.B(n_1060),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1088),
.A2(n_1085),
.B1(n_1080),
.B2(n_1098),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1048),
.Y(n_1191)
);

INVx4_ASAP7_75t_L g1192 ( 
.A(n_1030),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_1048),
.Y(n_1193)
);

INVx3_ASAP7_75t_SL g1194 ( 
.A(n_1030),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1070),
.B(n_1027),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1011),
.B(n_1023),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1070),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1060),
.B(n_1062),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1020),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1047),
.Y(n_1200)
);

OR2x6_ASAP7_75t_L g1201 ( 
.A(n_1045),
.B(n_1010),
.Y(n_1201)
);

NOR2xp67_ASAP7_75t_L g1202 ( 
.A(n_1034),
.B(n_1020),
.Y(n_1202)
);

AOI221x1_ASAP7_75t_L g1203 ( 
.A1(n_1024),
.A2(n_1003),
.B1(n_1001),
.B2(n_1021),
.C(n_1085),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_969),
.B(n_1088),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1080),
.A2(n_1003),
.B(n_972),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1062),
.B(n_1006),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1062),
.B(n_1006),
.Y(n_1207)
);

CKINVDCx16_ASAP7_75t_R g1208 ( 
.A(n_1040),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1028),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_972),
.A2(n_1001),
.B(n_969),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_989),
.Y(n_1211)
);

BUFx12f_ASAP7_75t_L g1212 ( 
.A(n_1047),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1047),
.Y(n_1213)
);

OR2x6_ASAP7_75t_L g1214 ( 
.A(n_1033),
.B(n_1024),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1047),
.Y(n_1215)
);

OR2x2_ASAP7_75t_L g1216 ( 
.A(n_1028),
.B(n_1021),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1033),
.B(n_1044),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1017),
.Y(n_1218)
);

NOR2x1_ASAP7_75t_SL g1219 ( 
.A(n_1044),
.B(n_1053),
.Y(n_1219)
);

AO21x1_ASAP7_75t_L g1220 ( 
.A1(n_1096),
.A2(n_954),
.B(n_1101),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1078),
.B(n_885),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_979),
.Y(n_1222)
);

INVx1_ASAP7_75t_SL g1223 ( 
.A(n_997),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1063),
.B(n_1066),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1091),
.A2(n_954),
.B(n_947),
.C(n_935),
.Y(n_1225)
);

OA21x2_ASAP7_75t_L g1226 ( 
.A1(n_998),
.A2(n_1024),
.B(n_1021),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1063),
.B(n_1066),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_967),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_967),
.Y(n_1229)
);

BUFx10_ASAP7_75t_L g1230 ( 
.A(n_1029),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_SL g1231 ( 
.A1(n_1067),
.A2(n_926),
.B(n_946),
.C(n_935),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1078),
.B(n_885),
.Y(n_1232)
);

INVx5_ASAP7_75t_L g1233 ( 
.A(n_1002),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_981),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1055),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1078),
.B(n_885),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_SL g1237 ( 
.A1(n_966),
.A2(n_947),
.B(n_954),
.C(n_1106),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1035),
.Y(n_1238)
);

INVx5_ASAP7_75t_L g1239 ( 
.A(n_1002),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1055),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1063),
.B(n_1066),
.Y(n_1241)
);

AOI21xp33_ASAP7_75t_L g1242 ( 
.A1(n_1096),
.A2(n_954),
.B(n_935),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_979),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_995),
.B(n_997),
.Y(n_1244)
);

NAND2x1p5_ASAP7_75t_L g1245 ( 
.A(n_1107),
.B(n_1002),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1078),
.B(n_885),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1002),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1055),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1063),
.B(n_1066),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1063),
.B(n_1066),
.Y(n_1250)
);

CKINVDCx8_ASAP7_75t_R g1251 ( 
.A(n_967),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_SL g1252 ( 
.A1(n_1067),
.A2(n_926),
.B(n_946),
.C(n_935),
.Y(n_1252)
);

AO21x1_ASAP7_75t_SL g1253 ( 
.A1(n_1182),
.A2(n_1242),
.B(n_1146),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1144),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1144),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1157),
.A2(n_1242),
.B1(n_1141),
.B2(n_1167),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1159),
.B(n_1221),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1113),
.Y(n_1258)
);

OR2x6_ASAP7_75t_L g1259 ( 
.A(n_1187),
.B(n_1201),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1157),
.A2(n_1167),
.B1(n_1220),
.B2(n_1112),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1225),
.A2(n_1151),
.B(n_1163),
.Y(n_1261)
);

OAI222xp33_ASAP7_75t_L g1262 ( 
.A1(n_1110),
.A2(n_1173),
.B1(n_1225),
.B2(n_1241),
.C1(n_1224),
.C2(n_1249),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1184),
.A2(n_1175),
.B1(n_1227),
.B2(n_1250),
.Y(n_1263)
);

CKINVDCx6p67_ASAP7_75t_R g1264 ( 
.A(n_1134),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_SL g1265 ( 
.A1(n_1224),
.A2(n_1241),
.B(n_1227),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1222),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1199),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_SL g1268 ( 
.A1(n_1208),
.A2(n_1230),
.B1(n_1250),
.B2(n_1249),
.Y(n_1268)
);

AOI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1202),
.A2(n_1217),
.B(n_1179),
.Y(n_1269)
);

OAI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1129),
.A2(n_1135),
.B1(n_1130),
.B2(n_1131),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1132),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1128),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_SL g1273 ( 
.A1(n_1172),
.A2(n_1146),
.B(n_1125),
.Y(n_1273)
);

BUFx8_ASAP7_75t_SL g1274 ( 
.A(n_1120),
.Y(n_1274)
);

BUFx10_ASAP7_75t_L g1275 ( 
.A(n_1221),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1143),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1126),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1117),
.B(n_1124),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1129),
.A2(n_1135),
.B1(n_1130),
.B2(n_1131),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1243),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1111),
.A2(n_1125),
.B1(n_1119),
.B2(n_1114),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1230),
.A2(n_1139),
.B1(n_1154),
.B2(n_1168),
.Y(n_1282)
);

NAND2x1p5_ASAP7_75t_L g1283 ( 
.A(n_1233),
.B(n_1239),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1182),
.A2(n_1160),
.B1(n_1169),
.B2(n_1161),
.Y(n_1284)
);

OAI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1111),
.A2(n_1145),
.B1(n_1118),
.B2(n_1223),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1166),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1156),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1165),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1177),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1244),
.B(n_1231),
.Y(n_1290)
);

AO21x1_ASAP7_75t_SL g1291 ( 
.A1(n_1198),
.A2(n_1172),
.B(n_1206),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1127),
.Y(n_1292)
);

NAND2x1p5_ASAP7_75t_L g1293 ( 
.A(n_1233),
.B(n_1239),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1142),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1234),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1228),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1162),
.A2(n_1181),
.B1(n_1223),
.B2(n_1118),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_SL g1298 ( 
.A(n_1115),
.Y(n_1298)
);

INVx1_ASAP7_75t_SL g1299 ( 
.A(n_1229),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1251),
.A2(n_1122),
.B1(n_1238),
.B2(n_1159),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1235),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1181),
.A2(n_1193),
.B1(n_1191),
.B2(n_1195),
.Y(n_1302)
);

INVx11_ASAP7_75t_L g1303 ( 
.A(n_1176),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1133),
.Y(n_1304)
);

OA21x2_ASAP7_75t_L g1305 ( 
.A1(n_1203),
.A2(n_1179),
.B(n_1171),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1240),
.Y(n_1306)
);

NAND2x1p5_ASAP7_75t_L g1307 ( 
.A(n_1233),
.B(n_1239),
.Y(n_1307)
);

AO21x1_ASAP7_75t_L g1308 ( 
.A1(n_1195),
.A2(n_1196),
.B(n_1147),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1150),
.A2(n_1140),
.B1(n_1138),
.B2(n_1136),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1183),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1148),
.B(n_1153),
.Y(n_1311)
);

INVx6_ASAP7_75t_L g1312 ( 
.A(n_1247),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1214),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_SL g1314 ( 
.A1(n_1171),
.A2(n_1206),
.B(n_1219),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1248),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1186),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1186),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1180),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1252),
.A2(n_1189),
.B1(n_1188),
.B2(n_1214),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1214),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1211),
.Y(n_1321)
);

AOI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1210),
.A2(n_1205),
.B(n_1147),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_1178),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1155),
.B(n_1137),
.Y(n_1324)
);

OAI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1209),
.A2(n_1185),
.B1(n_1237),
.B2(n_1198),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1194),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1232),
.Y(n_1327)
);

INVx4_ASAP7_75t_L g1328 ( 
.A(n_1247),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1236),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1164),
.A2(n_1246),
.B1(n_1201),
.B2(n_1209),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1164),
.A2(n_1212),
.B1(n_1190),
.B2(n_1226),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1205),
.A2(n_1149),
.B(n_1210),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1201),
.A2(n_1197),
.B1(n_1192),
.B2(n_1170),
.Y(n_1333)
);

BUFx4f_ASAP7_75t_SL g1334 ( 
.A(n_1152),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1207),
.B(n_1192),
.Y(n_1335)
);

INVx4_ASAP7_75t_L g1336 ( 
.A(n_1109),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1158),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1149),
.A2(n_1215),
.B(n_1190),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1109),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1121),
.A2(n_1245),
.B1(n_1174),
.B2(n_1216),
.Y(n_1340)
);

BUFx2_ASAP7_75t_SL g1341 ( 
.A(n_1109),
.Y(n_1341)
);

INVxp33_ASAP7_75t_L g1342 ( 
.A(n_1121),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1174),
.B(n_1204),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1226),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1109),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1245),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1200),
.Y(n_1347)
);

BUFx8_ASAP7_75t_L g1348 ( 
.A(n_1213),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1218),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1208),
.A2(n_727),
.B1(n_889),
.B2(n_470),
.Y(n_1350)
);

BUFx10_ASAP7_75t_L g1351 ( 
.A(n_1128),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1244),
.B(n_1118),
.Y(n_1352)
);

BUFx2_ASAP7_75t_R g1353 ( 
.A(n_1120),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1117),
.B(n_1124),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1126),
.Y(n_1355)
);

AOI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1151),
.A2(n_1076),
.B(n_1068),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1132),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1123),
.A2(n_985),
.B(n_987),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1157),
.A2(n_935),
.B1(n_946),
.B2(n_926),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1115),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1116),
.Y(n_1361)
);

CKINVDCx11_ASAP7_75t_R g1362 ( 
.A(n_1132),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1118),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1159),
.B(n_1221),
.Y(n_1364)
);

BUFx2_ASAP7_75t_R g1365 ( 
.A(n_1120),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1116),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1157),
.A2(n_935),
.B1(n_946),
.B2(n_926),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1348),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1291),
.B(n_1319),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1313),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1352),
.Y(n_1371)
);

AO31x2_ASAP7_75t_L g1372 ( 
.A1(n_1308),
.A2(n_1344),
.A3(n_1321),
.B(n_1320),
.Y(n_1372)
);

AO21x2_ASAP7_75t_L g1373 ( 
.A1(n_1322),
.A2(n_1314),
.B(n_1332),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1313),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1295),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1320),
.B(n_1259),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1347),
.B(n_1319),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1358),
.A2(n_1269),
.B(n_1356),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1256),
.B(n_1261),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1290),
.B(n_1302),
.Y(n_1380)
);

INVx3_ASAP7_75t_L g1381 ( 
.A(n_1338),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1295),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1302),
.B(n_1256),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1273),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1343),
.B(n_1260),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1338),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1348),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1266),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1343),
.B(n_1260),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1259),
.B(n_1257),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1348),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1257),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1276),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1325),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1325),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1305),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1258),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1257),
.Y(n_1398)
);

BUFx12f_ASAP7_75t_L g1399 ( 
.A(n_1362),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1276),
.Y(n_1400)
);

AO21x2_ASAP7_75t_L g1401 ( 
.A1(n_1270),
.A2(n_1335),
.B(n_1330),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1253),
.B(n_1263),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1267),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1280),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1289),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1267),
.B(n_1265),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1364),
.B(n_1349),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1305),
.A2(n_1340),
.B(n_1333),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1285),
.B(n_1297),
.Y(n_1409)
);

NAND2x1p5_ASAP7_75t_L g1410 ( 
.A(n_1336),
.B(n_1328),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1336),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1278),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1316),
.Y(n_1413)
);

OR2x6_ASAP7_75t_L g1414 ( 
.A(n_1341),
.B(n_1364),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1304),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1279),
.B(n_1263),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1310),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1364),
.B(n_1327),
.Y(n_1418)
);

OR2x6_ASAP7_75t_L g1419 ( 
.A(n_1300),
.B(n_1283),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1270),
.B(n_1281),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1287),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1339),
.Y(n_1422)
);

INVx1_ASAP7_75t_SL g1423 ( 
.A(n_1354),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1288),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1317),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1361),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1366),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1331),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1284),
.B(n_1297),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1359),
.B(n_1367),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1284),
.B(n_1282),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1339),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1268),
.B(n_1311),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1363),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1337),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_1312),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1283),
.A2(n_1307),
.B(n_1293),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1318),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1309),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1345),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1292),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1309),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1345),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1359),
.B(n_1367),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1307),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1296),
.B(n_1299),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1350),
.B(n_1277),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1324),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1396),
.B(n_1355),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1379),
.A2(n_1262),
.B1(n_1264),
.B2(n_1271),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1372),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1379),
.B(n_1346),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1406),
.B(n_1342),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1372),
.B(n_1254),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1372),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1372),
.B(n_1396),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1372),
.B(n_1255),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1403),
.Y(n_1458)
);

AOI222xp33_ASAP7_75t_L g1459 ( 
.A1(n_1444),
.A2(n_1362),
.B1(n_1294),
.B2(n_1271),
.C1(n_1357),
.C2(n_1298),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1386),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1369),
.B(n_1286),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1397),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1416),
.B(n_1329),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1381),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1369),
.B(n_1381),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1376),
.B(n_1323),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1394),
.B(n_1329),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1395),
.B(n_1323),
.Y(n_1468)
);

AND2x2_ASAP7_75t_SL g1469 ( 
.A(n_1383),
.B(n_1275),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1402),
.B(n_1370),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1377),
.B(n_1357),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1370),
.B(n_1374),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1374),
.B(n_1351),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1384),
.Y(n_1474)
);

AOI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1430),
.A2(n_1420),
.B1(n_1444),
.B2(n_1383),
.C(n_1395),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1377),
.B(n_1360),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1439),
.B(n_1442),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1375),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1374),
.B(n_1351),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1408),
.B(n_1306),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1408),
.B(n_1326),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1376),
.B(n_1326),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1376),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1382),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1401),
.B(n_1315),
.Y(n_1485)
);

OAI21xp33_ASAP7_75t_L g1486 ( 
.A1(n_1450),
.A2(n_1431),
.B(n_1380),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1451),
.A2(n_1378),
.B(n_1428),
.Y(n_1487)
);

OAI21xp5_ASAP7_75t_SL g1488 ( 
.A1(n_1450),
.A2(n_1431),
.B(n_1385),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1478),
.B(n_1393),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1475),
.A2(n_1419),
.B1(n_1380),
.B2(n_1403),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1465),
.B(n_1401),
.Y(n_1491)
);

NAND4xp25_ASAP7_75t_L g1492 ( 
.A(n_1475),
.B(n_1447),
.C(n_1439),
.D(n_1442),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1465),
.B(n_1401),
.Y(n_1493)
);

NAND3xp33_ASAP7_75t_L g1494 ( 
.A(n_1485),
.B(n_1428),
.C(n_1409),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1485),
.A2(n_1385),
.B(n_1389),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1465),
.B(n_1470),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1478),
.B(n_1371),
.Y(n_1497)
);

OAI21xp33_ASAP7_75t_L g1498 ( 
.A1(n_1485),
.A2(n_1389),
.B(n_1409),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1469),
.A2(n_1390),
.B1(n_1429),
.B2(n_1433),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1484),
.B(n_1400),
.Y(n_1500)
);

AOI21xp33_ASAP7_75t_L g1501 ( 
.A1(n_1453),
.A2(n_1433),
.B(n_1429),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1469),
.B(n_1407),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1458),
.B(n_1413),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1458),
.B(n_1476),
.Y(n_1504)
);

OAI221xp5_ASAP7_75t_SL g1505 ( 
.A1(n_1459),
.A2(n_1419),
.B1(n_1423),
.B2(n_1412),
.C(n_1446),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_R g1506 ( 
.A(n_1463),
.B(n_1272),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1462),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1483),
.B(n_1390),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1476),
.B(n_1425),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1483),
.B(n_1404),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1463),
.A2(n_1419),
.B1(n_1391),
.B2(n_1368),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1469),
.A2(n_1407),
.B1(n_1392),
.B2(n_1398),
.Y(n_1512)
);

NAND3xp33_ASAP7_75t_L g1513 ( 
.A(n_1459),
.B(n_1434),
.C(n_1446),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1469),
.A2(n_1407),
.B1(n_1398),
.B2(n_1392),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1453),
.A2(n_1419),
.B1(n_1368),
.B2(n_1391),
.Y(n_1515)
);

AOI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1467),
.A2(n_1419),
.B1(n_1407),
.B2(n_1448),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_R g1517 ( 
.A(n_1471),
.B(n_1272),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1482),
.B(n_1418),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1476),
.B(n_1415),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1472),
.B(n_1405),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1472),
.B(n_1405),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1471),
.B(n_1441),
.Y(n_1522)
);

AOI221xp5_ASAP7_75t_L g1523 ( 
.A1(n_1468),
.A2(n_1415),
.B1(n_1417),
.B2(n_1427),
.C(n_1421),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1472),
.B(n_1417),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1467),
.A2(n_1387),
.B1(n_1414),
.B2(n_1422),
.Y(n_1525)
);

NAND3xp33_ASAP7_75t_L g1526 ( 
.A(n_1468),
.B(n_1427),
.C(n_1421),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1460),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1481),
.A2(n_1392),
.B1(n_1398),
.B2(n_1418),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1471),
.B(n_1424),
.C(n_1426),
.Y(n_1529)
);

OAI221xp5_ASAP7_75t_L g1530 ( 
.A1(n_1477),
.A2(n_1294),
.B1(n_1387),
.B2(n_1443),
.C(n_1422),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1452),
.B(n_1424),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1481),
.A2(n_1437),
.B(n_1445),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1454),
.B(n_1373),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1473),
.B(n_1388),
.Y(n_1534)
);

OAI221xp5_ASAP7_75t_L g1535 ( 
.A1(n_1477),
.A2(n_1387),
.B1(n_1443),
.B2(n_1422),
.C(n_1414),
.Y(n_1535)
);

AOI211xp5_ASAP7_75t_SL g1536 ( 
.A1(n_1481),
.A2(n_1411),
.B(n_1432),
.C(n_1418),
.Y(n_1536)
);

NAND3xp33_ASAP7_75t_L g1537 ( 
.A(n_1480),
.B(n_1435),
.C(n_1438),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1454),
.B(n_1373),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1527),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1507),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1507),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1491),
.B(n_1454),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1527),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1520),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1496),
.B(n_1456),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1491),
.B(n_1457),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1520),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1521),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1510),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1496),
.B(n_1456),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1524),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1493),
.B(n_1457),
.Y(n_1552)
);

NAND2x1p5_ASAP7_75t_L g1553 ( 
.A(n_1502),
.B(n_1457),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1504),
.B(n_1449),
.Y(n_1554)
);

NOR2x1_ASAP7_75t_L g1555 ( 
.A(n_1526),
.B(n_1474),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1533),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1493),
.B(n_1456),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1533),
.B(n_1451),
.Y(n_1558)
);

INVxp67_ASAP7_75t_SL g1559 ( 
.A(n_1526),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1538),
.B(n_1451),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1537),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1529),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1529),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_1508),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1517),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1489),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1487),
.Y(n_1567)
);

NAND2x1_ASAP7_75t_L g1568 ( 
.A(n_1532),
.B(n_1474),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1531),
.B(n_1480),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1534),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1487),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1518),
.B(n_1464),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1503),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1498),
.B(n_1474),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1487),
.B(n_1455),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1500),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1573),
.B(n_1566),
.Y(n_1577)
);

AOI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1565),
.A2(n_1486),
.B1(n_1498),
.B2(n_1488),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1540),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1573),
.B(n_1522),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1557),
.B(n_1508),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1557),
.B(n_1536),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1557),
.B(n_1487),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1540),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1566),
.B(n_1519),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1545),
.B(n_1495),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1541),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1541),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1562),
.Y(n_1589)
);

INVxp67_ASAP7_75t_SL g1590 ( 
.A(n_1555),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1543),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1576),
.B(n_1497),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1545),
.B(n_1461),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1576),
.B(n_1494),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1543),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1545),
.B(n_1461),
.Y(n_1596)
);

OAI211xp5_ASAP7_75t_L g1597 ( 
.A1(n_1559),
.A2(n_1486),
.B(n_1513),
.C(n_1501),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1550),
.B(n_1461),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1549),
.Y(n_1599)
);

AND2x6_ASAP7_75t_SL g1600 ( 
.A(n_1565),
.B(n_1274),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1549),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1544),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1554),
.B(n_1399),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1550),
.B(n_1482),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1570),
.B(n_1509),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1564),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1544),
.Y(n_1607)
);

NOR2x1p5_ASAP7_75t_L g1608 ( 
.A(n_1568),
.B(n_1399),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1547),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1547),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1551),
.Y(n_1611)
);

INVxp67_ASAP7_75t_SL g1612 ( 
.A(n_1555),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_SL g1613 ( 
.A(n_1559),
.B(n_1505),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1551),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1562),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1548),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1579),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1578),
.B(n_1561),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1594),
.B(n_1561),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1613),
.B(n_1563),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1582),
.B(n_1558),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1589),
.Y(n_1622)
);

AND2x4_ASAP7_75t_SL g1623 ( 
.A(n_1582),
.B(n_1482),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1579),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1586),
.B(n_1558),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1586),
.B(n_1574),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1604),
.B(n_1558),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1584),
.Y(n_1628)
);

NAND3xp33_ASAP7_75t_L g1629 ( 
.A(n_1597),
.B(n_1513),
.C(n_1563),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1580),
.B(n_1574),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1600),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1584),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1604),
.B(n_1560),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1606),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1577),
.B(n_1554),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1592),
.B(n_1570),
.Y(n_1636)
);

NAND2x1p5_ASAP7_75t_L g1637 ( 
.A(n_1608),
.B(n_1568),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1587),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1581),
.B(n_1560),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1605),
.B(n_1569),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1585),
.B(n_1542),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1587),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1581),
.Y(n_1643)
);

NOR2x1_ASAP7_75t_L g1644 ( 
.A(n_1615),
.B(n_1530),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1588),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1606),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1588),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1590),
.A2(n_1612),
.B(n_1615),
.Y(n_1648)
);

OAI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1603),
.A2(n_1490),
.B1(n_1492),
.B2(n_1516),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1593),
.B(n_1560),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1602),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1602),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1599),
.Y(n_1653)
);

AOI32xp33_ASAP7_75t_L g1654 ( 
.A1(n_1583),
.A2(n_1575),
.A3(n_1511),
.B1(n_1572),
.B2(n_1515),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1607),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1593),
.B(n_1556),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1601),
.B(n_1542),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1607),
.B(n_1546),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1609),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1631),
.B(n_1274),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1621),
.B(n_1596),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1634),
.B(n_1596),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1647),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1634),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1644),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1646),
.Y(n_1666)
);

BUFx3_ASAP7_75t_L g1667 ( 
.A(n_1646),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1647),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1618),
.B(n_1598),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1622),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1619),
.B(n_1609),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1626),
.B(n_1610),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1621),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1637),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1623),
.Y(n_1675)
);

AND2x4_ASAP7_75t_SL g1676 ( 
.A(n_1643),
.B(n_1482),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1623),
.B(n_1598),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1617),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1620),
.B(n_1546),
.Y(n_1679)
);

BUFx2_ASAP7_75t_SL g1680 ( 
.A(n_1643),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1629),
.B(n_1552),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1624),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1630),
.B(n_1353),
.Y(n_1683)
);

CKINVDCx16_ASAP7_75t_R g1684 ( 
.A(n_1648),
.Y(n_1684)
);

AO21x2_ASAP7_75t_L g1685 ( 
.A1(n_1649),
.A2(n_1571),
.B(n_1567),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1653),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1628),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1639),
.B(n_1583),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1636),
.B(n_1552),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1651),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1641),
.B(n_1610),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1637),
.Y(n_1692)
);

INVxp67_ASAP7_75t_SL g1693 ( 
.A(n_1652),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1657),
.B(n_1611),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1632),
.Y(n_1695)
);

AOI32xp33_ASAP7_75t_L g1696 ( 
.A1(n_1665),
.A2(n_1649),
.A3(n_1625),
.B1(n_1654),
.B2(n_1575),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1668),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1668),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_R g1699 ( 
.A(n_1660),
.B(n_1301),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1670),
.B(n_1640),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1684),
.A2(n_1499),
.B1(n_1506),
.B2(n_1625),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1681),
.A2(n_1525),
.B1(n_1516),
.B2(n_1638),
.Y(n_1702)
);

OR4x1_ASAP7_75t_L g1703 ( 
.A(n_1663),
.B(n_1642),
.C(n_1645),
.D(n_1655),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1690),
.Y(n_1704)
);

OA21x2_ASAP7_75t_L g1705 ( 
.A1(n_1664),
.A2(n_1659),
.B(n_1571),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1674),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1678),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1674),
.B(n_1635),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1685),
.A2(n_1575),
.B1(n_1553),
.B2(n_1455),
.Y(n_1709)
);

NOR3xp33_ASAP7_75t_L g1710 ( 
.A(n_1686),
.B(n_1315),
.C(n_1523),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1685),
.A2(n_1658),
.B(n_1571),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1678),
.Y(n_1712)
);

XNOR2xp5_ASAP7_75t_L g1713 ( 
.A(n_1673),
.B(n_1466),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1667),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1682),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1692),
.B(n_1553),
.Y(n_1716)
);

OAI322xp33_ASAP7_75t_L g1717 ( 
.A1(n_1693),
.A2(n_1658),
.A3(n_1567),
.B1(n_1553),
.B2(n_1611),
.C1(n_1614),
.C2(n_1595),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1675),
.B(n_1639),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1675),
.B(n_1627),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1682),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1669),
.B(n_1627),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1687),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1714),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1714),
.B(n_1683),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1706),
.B(n_1664),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1699),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1718),
.B(n_1667),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1704),
.B(n_1666),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1707),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1721),
.B(n_1679),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1712),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1703),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1700),
.B(n_1689),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1708),
.B(n_1671),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1697),
.B(n_1675),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1715),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1710),
.B(n_1666),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1710),
.B(n_1661),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1701),
.B(n_1671),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1719),
.B(n_1661),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1701),
.B(n_1662),
.Y(n_1741)
);

INVx3_ASAP7_75t_L g1742 ( 
.A(n_1705),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1698),
.B(n_1680),
.Y(n_1743)
);

NOR3x1_ASAP7_75t_L g1744 ( 
.A(n_1737),
.B(n_1716),
.C(n_1720),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1732),
.A2(n_1696),
.B(n_1685),
.Y(n_1745)
);

OAI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1726),
.A2(n_1739),
.B1(n_1732),
.B2(n_1724),
.C(n_1738),
.Y(n_1746)
);

OAI21xp33_ASAP7_75t_L g1747 ( 
.A1(n_1741),
.A2(n_1709),
.B(n_1716),
.Y(n_1747)
);

AOI211x1_ASAP7_75t_SL g1748 ( 
.A1(n_1723),
.A2(n_1711),
.B(n_1680),
.C(n_1717),
.Y(n_1748)
);

NAND2x1_ASAP7_75t_L g1749 ( 
.A(n_1727),
.B(n_1677),
.Y(n_1749)
);

O2A1O1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1725),
.A2(n_1722),
.B(n_1709),
.C(n_1687),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_SL g1751 ( 
.A(n_1734),
.B(n_1699),
.Y(n_1751)
);

AND4x1_ASAP7_75t_L g1752 ( 
.A(n_1724),
.B(n_1702),
.C(n_1365),
.D(n_1695),
.Y(n_1752)
);

OAI21xp33_ASAP7_75t_L g1753 ( 
.A1(n_1741),
.A2(n_1713),
.B(n_1695),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_R g1754 ( 
.A(n_1723),
.B(n_1301),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1730),
.A2(n_1677),
.B1(n_1662),
.B2(n_1676),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1727),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1756),
.B(n_1728),
.Y(n_1757)
);

AND4x1_ASAP7_75t_L g1758 ( 
.A(n_1748),
.B(n_1743),
.C(n_1735),
.D(n_1736),
.Y(n_1758)
);

AOI211xp5_ASAP7_75t_L g1759 ( 
.A1(n_1745),
.A2(n_1743),
.B(n_1735),
.C(n_1731),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1751),
.B(n_1740),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1747),
.A2(n_1733),
.B1(n_1729),
.B2(n_1677),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1749),
.Y(n_1762)
);

NAND3xp33_ASAP7_75t_SL g1763 ( 
.A(n_1754),
.B(n_1750),
.C(n_1746),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1752),
.B(n_1672),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1753),
.Y(n_1765)
);

NOR3xp33_ASAP7_75t_L g1766 ( 
.A(n_1755),
.B(n_1742),
.C(n_1672),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1744),
.B(n_1662),
.Y(n_1767)
);

NAND5xp2_ASAP7_75t_L g1768 ( 
.A(n_1746),
.B(n_1512),
.C(n_1514),
.D(n_1553),
.E(n_1528),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1762),
.B(n_1676),
.Y(n_1769)
);

NOR3xp33_ASAP7_75t_L g1770 ( 
.A(n_1763),
.B(n_1742),
.C(n_1691),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1767),
.A2(n_1760),
.B(n_1759),
.Y(n_1771)
);

OAI211xp5_ASAP7_75t_SL g1772 ( 
.A1(n_1765),
.A2(n_1742),
.B(n_1691),
.C(n_1694),
.Y(n_1772)
);

NAND4xp75_ASAP7_75t_L g1773 ( 
.A(n_1761),
.B(n_1705),
.C(n_1298),
.D(n_1633),
.Y(n_1773)
);

OAI211xp5_ASAP7_75t_SL g1774 ( 
.A1(n_1757),
.A2(n_1694),
.B(n_1535),
.C(n_1705),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1766),
.B(n_1688),
.Y(n_1775)
);

AOI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1770),
.A2(n_1764),
.B1(n_1769),
.B2(n_1775),
.Y(n_1776)
);

NOR2x1_ASAP7_75t_L g1777 ( 
.A(n_1771),
.B(n_1772),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1773),
.B(n_1758),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1774),
.B(n_1688),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1775),
.Y(n_1780)
);

INVxp67_ASAP7_75t_SL g1781 ( 
.A(n_1775),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1775),
.Y(n_1782)
);

CKINVDCx20_ASAP7_75t_R g1783 ( 
.A(n_1776),
.Y(n_1783)
);

OAI221xp5_ASAP7_75t_SL g1784 ( 
.A1(n_1779),
.A2(n_1768),
.B1(n_1633),
.B2(n_1650),
.C(n_1656),
.Y(n_1784)
);

NAND3xp33_ASAP7_75t_L g1785 ( 
.A(n_1777),
.B(n_1688),
.C(n_1567),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_SL g1786 ( 
.A(n_1780),
.B(n_1410),
.C(n_1303),
.Y(n_1786)
);

NOR3xp33_ASAP7_75t_L g1787 ( 
.A(n_1781),
.B(n_1479),
.C(n_1473),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1782),
.Y(n_1788)
);

XNOR2xp5_ASAP7_75t_L g1789 ( 
.A(n_1783),
.B(n_1778),
.Y(n_1789)
);

XOR2xp5_ASAP7_75t_L g1790 ( 
.A(n_1786),
.B(n_1466),
.Y(n_1790)
);

AND2x4_ASAP7_75t_SL g1791 ( 
.A(n_1788),
.B(n_1656),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1791),
.Y(n_1792)
);

NOR3xp33_ASAP7_75t_L g1793 ( 
.A(n_1792),
.B(n_1789),
.C(n_1784),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1793),
.Y(n_1794)
);

BUFx2_ASAP7_75t_L g1795 ( 
.A(n_1793),
.Y(n_1795)
);

AOI21x1_ASAP7_75t_L g1796 ( 
.A1(n_1795),
.A2(n_1785),
.B(n_1790),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1794),
.B(n_1787),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1796),
.B(n_1650),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1797),
.A2(n_1614),
.B(n_1616),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1798),
.A2(n_1334),
.B1(n_1616),
.B2(n_1595),
.Y(n_1800)
);

AOI222xp33_ASAP7_75t_L g1801 ( 
.A1(n_1800),
.A2(n_1799),
.B1(n_1591),
.B2(n_1334),
.C1(n_1479),
.C2(n_1436),
.Y(n_1801)
);

OAI221xp5_ASAP7_75t_R g1802 ( 
.A1(n_1801),
.A2(n_1591),
.B1(n_1564),
.B2(n_1539),
.C(n_1410),
.Y(n_1802)
);

AOI211xp5_ASAP7_75t_L g1803 ( 
.A1(n_1802),
.A2(n_1436),
.B(n_1440),
.C(n_1479),
.Y(n_1803)
);


endmodule