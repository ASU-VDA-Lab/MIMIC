module fake_jpeg_3076_n_169 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_58),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_69),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_56),
.B1(n_58),
.B2(n_55),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_74),
.B1(n_54),
.B2(n_62),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_58),
.B1(n_49),
.B2(n_50),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_75),
.A2(n_63),
.B1(n_64),
.B2(n_62),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_48),
.B1(n_18),
.B2(n_21),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

OR2x2_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_86),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_91),
.Y(n_97)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_72),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_54),
.B1(n_47),
.B2(n_52),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_93),
.Y(n_99)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_57),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_110),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_46),
.B1(n_45),
.B2(n_52),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_105),
.B1(n_24),
.B2(n_41),
.Y(n_112)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_0),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_4),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_48),
.B1(n_2),
.B2(n_3),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_108),
.A2(n_111),
.B1(n_4),
.B2(n_5),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_1),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_101),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_79),
.B(n_3),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_48),
.B1(n_5),
.B2(n_6),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_114),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_118),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_117),
.Y(n_139)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_22),
.C(n_39),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_125),
.Y(n_137)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_122),
.A2(n_106),
.B1(n_108),
.B2(n_12),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_129),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_6),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_26),
.C(n_38),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_118),
.C(n_130),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_127),
.A2(n_13),
.B1(n_16),
.B2(n_28),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_128),
.A2(n_130),
.B(n_12),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_10),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_30),
.B(n_37),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_144),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_140),
.B(n_142),
.Y(n_148)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_115),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_29),
.B(n_15),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_31),
.B(n_34),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_150),
.B(n_133),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_13),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_152),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_153),
.A2(n_143),
.B(n_138),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_158),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_153),
.C(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_147),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_160),
.C(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_162),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_151),
.B1(n_135),
.B2(n_134),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_163),
.B(n_151),
.Y(n_165)
);

OAI221xp5_ASAP7_75t_SL g166 ( 
.A1(n_165),
.A2(n_157),
.B1(n_136),
.B2(n_137),
.C(n_145),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_139),
.C(n_35),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_167),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_42),
.Y(n_169)
);


endmodule