module fake_jpeg_3674_n_124 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_124);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_4),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_31),
.B(n_34),
.Y(n_58)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_9),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_41),
.Y(n_43)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_19),
.B(n_25),
.C(n_22),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_46),
.B(n_47),
.C(n_51),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_18),
.B1(n_23),
.B2(n_26),
.Y(n_46)
);

NOR2x1_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_28),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_27),
.B1(n_19),
.B2(n_25),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_42),
.B1(n_24),
.B2(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_20),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_61),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_29),
.A2(n_22),
.B1(n_21),
.B2(n_20),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_46),
.B1(n_30),
.B2(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_21),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_69),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_70),
.B1(n_75),
.B2(n_78),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_71),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_10),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_74),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_53),
.B(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_44),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_42),
.B1(n_41),
.B2(n_0),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_10),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_50),
.A2(n_41),
.B1(n_1),
.B2(n_0),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_53),
.B1(n_60),
.B2(n_49),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_89),
.B1(n_72),
.B2(n_69),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_49),
.B1(n_41),
.B2(n_11),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_66),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_94),
.Y(n_100)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_63),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_83),
.C(n_86),
.Y(n_101)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_99),
.A2(n_88),
.B(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_101),
.B(n_92),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_99),
.B(n_86),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_104),
.C(n_75),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_89),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_95),
.B(n_73),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_108),
.B(n_110),
.Y(n_113)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_111),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_100),
.B(n_2),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_104),
.C(n_102),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_112),
.C(n_105),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_117),
.C(n_114),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_105),
.C(n_62),
.Y(n_117)
);

AO21x1_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_119),
.B(n_80),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_80),
.B1(n_70),
.B2(n_65),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_79),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_3),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_12),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);


endmodule