module fake_jpeg_31690_n_502 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_502);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_502;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_29),
.B(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_56),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_61),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_60),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_29),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_62),
.B(n_83),
.Y(n_127)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_67),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_66),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_68),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_73),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_19),
.B(n_0),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_74),
.Y(n_159)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_76),
.B(n_87),
.Y(n_129)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx24_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_39),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_80),
.B(n_89),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_22),
.B(n_0),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_25),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_24),
.B(n_0),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_99),
.Y(n_138)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_24),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_18),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_18),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_49),
.Y(n_150)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_102),
.B(n_18),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_18),
.Y(n_103)
);

INVx6_ASAP7_75t_SL g124 ( 
.A(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_100),
.B(n_31),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_104),
.B(n_113),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_108),
.B(n_142),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_100),
.B(n_31),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_49),
.B1(n_28),
.B2(n_42),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_118),
.A2(n_157),
.B1(n_80),
.B2(n_63),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_60),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_119),
.B(n_132),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_77),
.B(n_1),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_122),
.B(n_26),
.C(n_54),
.Y(n_198)
);

INVx6_ASAP7_75t_SL g126 ( 
.A(n_60),
.Y(n_126)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_126),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_86),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_79),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_140),
.B(n_150),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_92),
.B(n_30),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_93),
.B(n_30),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_146),
.B(n_154),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_89),
.B(n_22),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_103),
.A2(n_49),
.B(n_28),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_163),
.B(n_139),
.C(n_118),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_103),
.A2(n_49),
.B1(n_42),
.B2(n_40),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_96),
.B(n_44),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_162),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_69),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_164),
.Y(n_261)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_165),
.Y(n_248)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_112),
.B1(n_85),
.B2(n_88),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_168),
.A2(n_209),
.B1(n_158),
.B2(n_155),
.Y(n_255)
);

NAND2xp33_ASAP7_75t_SL g169 ( 
.A(n_156),
.B(n_98),
.Y(n_169)
);

NAND2xp33_ASAP7_75t_SL g224 ( 
.A(n_169),
.B(n_174),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_127),
.B(n_44),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_170),
.B(n_201),
.Y(n_250)
);

AOI32xp33_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_109),
.A3(n_121),
.B1(n_106),
.B2(n_129),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_171),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_260)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_125),
.Y(n_172)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_172),
.Y(n_221)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_173),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_157),
.A2(n_82),
.B1(n_84),
.B2(n_90),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_175),
.A2(n_205),
.B1(n_144),
.B2(n_143),
.Y(n_239)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_178),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_179),
.Y(n_249)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_180),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_128),
.Y(n_181)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_181),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_122),
.B(n_27),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_186),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_105),
.B(n_27),
.Y(n_186)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_110),
.Y(n_188)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_188),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_95),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_192),
.C(n_198),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_139),
.B(n_75),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_195),
.Y(n_229)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_133),
.Y(n_191)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_191),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_115),
.B(n_91),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_141),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_194),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_111),
.B(n_78),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_196),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_197),
.A2(n_136),
.B1(n_152),
.B2(n_144),
.Y(n_233)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_200),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_151),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_116),
.B(n_26),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_207),
.Y(n_236)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_116),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_204),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_120),
.A2(n_59),
.B1(n_68),
.B2(n_66),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_151),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_120),
.A2(n_53),
.B1(n_52),
.B2(n_64),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_149),
.Y(n_211)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_211),
.Y(n_262)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_212),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_137),
.A2(n_42),
.B1(n_40),
.B2(n_33),
.Y(n_213)
);

AOI32xp33_ASAP7_75t_L g245 ( 
.A1(n_213),
.A2(n_218),
.A3(n_117),
.B1(n_124),
.B2(n_147),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_135),
.B(n_78),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_215),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_135),
.B(n_42),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_141),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_217),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_116),
.B(n_40),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_137),
.A2(n_40),
.B1(n_33),
.B2(n_72),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_136),
.B(n_33),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_124),
.Y(n_240)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_166),
.B(n_147),
.C(n_126),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_174),
.C(n_168),
.Y(n_268)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_182),
.B(n_148),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_231),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_233),
.A2(n_239),
.B1(n_209),
.B2(n_213),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_240),
.B(n_260),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_177),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_242),
.B(n_202),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_169),
.A2(n_152),
.B1(n_117),
.B2(n_161),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_244),
.A2(n_255),
.B1(n_134),
.B2(n_130),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_245),
.A2(n_191),
.B1(n_165),
.B2(n_188),
.Y(n_301)
);

OAI32xp33_ASAP7_75t_L g254 ( 
.A1(n_210),
.A2(n_33),
.A3(n_147),
.B1(n_114),
.B2(n_155),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_175),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_186),
.B(n_158),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_259),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_198),
.B(n_145),
.Y(n_259)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_265),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_266),
.A2(n_274),
.B1(n_282),
.B2(n_239),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_268),
.B(n_260),
.Y(n_317)
);

OAI22x1_ASAP7_75t_L g269 ( 
.A1(n_224),
.A2(n_218),
.B1(n_185),
.B2(n_187),
.Y(n_269)
);

OA21x2_ASAP7_75t_L g325 ( 
.A1(n_269),
.A2(n_270),
.B(n_241),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g270 ( 
.A1(n_224),
.A2(n_189),
.B(n_192),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_219),
.C(n_189),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_271),
.B(n_284),
.C(n_226),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_206),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_286),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_236),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_280),
.Y(n_324)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_230),
.Y(n_276)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_276),
.Y(n_311)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

BUFx6f_ASAP7_75t_SL g278 ( 
.A(n_252),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_278),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_279),
.B(n_291),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_208),
.Y(n_280)
);

INVx13_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_281),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_L g282 ( 
.A1(n_240),
.A2(n_134),
.B1(n_130),
.B2(n_145),
.Y(n_282)
);

BUFx8_ASAP7_75t_L g283 ( 
.A(n_235),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_283),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_227),
.B(n_172),
.C(n_167),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_285),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_225),
.B(n_184),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_225),
.B(n_176),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_290),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_250),
.Y(n_288)
);

NOR3xp33_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_292),
.C(n_293),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_255),
.A2(n_192),
.B1(n_200),
.B2(n_181),
.Y(n_289)
);

OAI21xp33_ASAP7_75t_SL g302 ( 
.A1(n_289),
.A2(n_301),
.B(n_245),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_253),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_229),
.B(n_208),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_251),
.Y(n_292)
);

AND2x6_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_178),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_230),
.Y(n_294)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_294),
.Y(n_327)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_220),
.Y(n_295)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_295),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_231),
.A2(n_181),
.B(n_183),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_296),
.A2(n_297),
.B(n_237),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_226),
.A2(n_183),
.B(n_178),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_298),
.A2(n_179),
.B1(n_164),
.B2(n_222),
.Y(n_328)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_237),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_299),
.B(n_300),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_234),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_302),
.A2(n_328),
.B1(n_285),
.B2(n_216),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_305),
.B(n_316),
.C(n_323),
.Y(n_346)
);

OAI21xp33_ASAP7_75t_SL g307 ( 
.A1(n_269),
.A2(n_231),
.B(n_233),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_SL g351 ( 
.A(n_307),
.B(n_283),
.C(n_281),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_308),
.A2(n_319),
.B(n_270),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_310),
.A2(n_312),
.B1(n_314),
.B2(n_330),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_274),
.A2(n_257),
.B1(n_262),
.B2(n_263),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_298),
.A2(n_257),
.B1(n_223),
.B2(n_161),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_272),
.B(n_263),
.C(n_262),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_317),
.B(n_333),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_288),
.B(n_232),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_318),
.B(n_279),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_296),
.A2(n_222),
.B(n_248),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_272),
.B(n_234),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_320),
.B(n_322),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_273),
.B(n_287),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_284),
.B(n_241),
.C(n_238),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_301),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_282),
.A2(n_223),
.B1(n_238),
.B2(n_249),
.Y(n_330)
);

MAJx2_ASAP7_75t_L g333 ( 
.A(n_268),
.B(n_248),
.C(n_232),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_325),
.A2(n_264),
.B(n_267),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_335),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_355),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_271),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_327),
.C(n_309),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_338),
.A2(n_345),
.B(n_352),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_300),
.Y(n_339)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_339),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_340),
.B(n_347),
.Y(n_386)
);

A2O1A1Ixp33_ASAP7_75t_L g341 ( 
.A1(n_303),
.A2(n_297),
.B(n_286),
.C(n_264),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_341),
.B(n_349),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_332),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_342),
.B(n_348),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_292),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_343),
.Y(n_394)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_332),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_344),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_308),
.A2(n_270),
.B(n_290),
.Y(n_345)
);

O2A1O1Ixp33_ASAP7_75t_L g347 ( 
.A1(n_319),
.A2(n_293),
.B(n_289),
.C(n_278),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_324),
.Y(n_348)
);

FAx1_ASAP7_75t_SL g349 ( 
.A(n_303),
.B(n_267),
.CI(n_279),
.CON(n_349),
.SN(n_349)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_350),
.A2(n_334),
.B1(n_249),
.B2(n_261),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_351),
.A2(n_334),
.B1(n_235),
.B2(n_331),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_304),
.A2(n_299),
.B(n_276),
.Y(n_352)
);

OR2x2_ASAP7_75t_L g353 ( 
.A(n_306),
.B(n_283),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_353),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_310),
.A2(n_312),
.B1(n_320),
.B2(n_330),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_354),
.A2(n_358),
.B1(n_336),
.B2(n_344),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_283),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_304),
.B(n_294),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_356),
.Y(n_385)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_311),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_357),
.B(n_361),
.Y(n_382)
);

INVx13_ASAP7_75t_L g359 ( 
.A(n_329),
.Y(n_359)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_359),
.Y(n_377)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_313),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_295),
.Y(n_363)
);

NOR2x1_ASAP7_75t_L g384 ( 
.A(n_363),
.B(n_331),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_321),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_364),
.B(n_365),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_322),
.B(n_243),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_316),
.Y(n_370)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_370),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_372),
.A2(n_353),
.B1(n_365),
.B2(n_362),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_374),
.B(n_379),
.Y(n_411)
);

NOR4xp25_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_333),
.C(n_317),
.D(n_323),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_375),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_376),
.B(n_380),
.C(n_393),
.Y(n_399)
);

NAND3xp33_ASAP7_75t_L g379 ( 
.A(n_348),
.B(n_309),
.C(n_326),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_337),
.B(n_327),
.C(n_313),
.Y(n_380)
);

AOI22x1_ASAP7_75t_SL g381 ( 
.A1(n_351),
.A2(n_328),
.B1(n_326),
.B2(n_315),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_381),
.A2(n_390),
.B1(n_199),
.B2(n_258),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_384),
.A2(n_228),
.B(n_221),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_357),
.Y(n_387)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_387),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_388),
.B(n_349),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_364),
.B(n_277),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_389),
.B(n_392),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_265),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_360),
.B(n_258),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_371),
.A2(n_354),
.B1(n_358),
.B2(n_336),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_396),
.A2(n_400),
.B1(n_402),
.B2(n_406),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_386),
.A2(n_355),
.B(n_339),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g423 ( 
.A(n_398),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_371),
.A2(n_355),
.B1(n_342),
.B2(n_338),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_394),
.A2(n_350),
.B1(n_339),
.B2(n_335),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_401),
.A2(n_403),
.B1(n_404),
.B2(n_417),
.Y(n_438)
);

OAI22x1_ASAP7_75t_L g402 ( 
.A1(n_381),
.A2(n_347),
.B1(n_345),
.B2(n_353),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_394),
.A2(n_362),
.B1(n_341),
.B2(n_349),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_405),
.A2(n_416),
.B1(n_390),
.B2(n_366),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_383),
.A2(n_347),
.B1(n_360),
.B2(n_361),
.Y(n_406)
);

XOR2x2_ASAP7_75t_L g407 ( 
.A(n_375),
.B(n_346),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_413),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_385),
.B(n_346),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_408),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_383),
.A2(n_363),
.B1(n_359),
.B2(n_243),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_377),
.Y(n_433)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_377),
.Y(n_412)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_412),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_385),
.B(n_363),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_359),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_414),
.B(n_400),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_372),
.A2(n_228),
.B1(n_221),
.B2(n_220),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_418),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_380),
.C(n_376),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_421),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_399),
.B(n_369),
.C(n_391),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_424),
.A2(n_384),
.B(n_382),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_425),
.B(n_427),
.Y(n_441)
);

INVxp33_ASAP7_75t_SL g426 ( 
.A(n_402),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_426),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_407),
.B(n_369),
.C(n_391),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_405),
.B(n_373),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_428),
.B(n_434),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_388),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_429),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_433),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_386),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_406),
.B(n_366),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_436),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_397),
.B(n_368),
.C(n_373),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_415),
.B(n_368),
.C(n_366),
.Y(n_437)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_437),
.Y(n_440)
);

AOI322xp5_ASAP7_75t_L g439 ( 
.A1(n_426),
.A2(n_415),
.A3(n_395),
.B1(n_367),
.B2(n_382),
.C1(n_378),
.C2(n_416),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_442),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_378),
.Y(n_442)
);

INVx13_ASAP7_75t_L g443 ( 
.A(n_431),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_443),
.B(n_436),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_422),
.A2(n_403),
.B1(n_405),
.B2(n_398),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_445),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_423),
.A2(n_417),
.B1(n_384),
.B2(n_396),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_424),
.A2(n_418),
.B(n_410),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_446),
.A2(n_212),
.B(n_203),
.Y(n_466)
);

OAI22xp33_ASAP7_75t_SL g448 ( 
.A1(n_430),
.A2(n_412),
.B1(n_387),
.B2(n_409),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_448),
.A2(n_437),
.B1(n_428),
.B2(n_196),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_453),
.B(n_435),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_456),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_447),
.B(n_427),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_450),
.B(n_438),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_461),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_459),
.B(n_464),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_440),
.B(n_421),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_419),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_462),
.B(n_463),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_441),
.B(n_434),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_446),
.A2(n_420),
.B1(n_194),
.B2(n_180),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_465),
.B(n_440),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_466),
.A2(n_453),
.B(n_442),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_454),
.B(n_2),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_467),
.B(n_5),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_3),
.C(n_5),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_468),
.B(n_454),
.C(n_451),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_471),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_474),
.B(n_476),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_458),
.A2(n_450),
.B(n_449),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_475),
.A2(n_460),
.B(n_468),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_462),
.B(n_444),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_478),
.B(n_479),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_452),
.C(n_451),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_473),
.C(n_479),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_481),
.B(n_486),
.Y(n_491)
);

OAI21x1_ASAP7_75t_SL g483 ( 
.A1(n_472),
.A2(n_443),
.B(n_465),
.Y(n_483)
);

AOI322xp5_ASAP7_75t_L g488 ( 
.A1(n_483),
.A2(n_485),
.A3(n_487),
.B1(n_477),
.B2(n_445),
.C1(n_7),
.C2(n_8),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_474),
.B(n_478),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_473),
.B(n_459),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_488),
.A2(n_492),
.B(n_9),
.Y(n_495)
);

AOI322xp5_ASAP7_75t_L g489 ( 
.A1(n_487),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_489),
.A2(n_490),
.B(n_482),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_484),
.B(n_6),
.C(n_7),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_480),
.B(n_6),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_493),
.B(n_494),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_491),
.A2(n_7),
.B(n_8),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_495),
.B(n_10),
.C(n_11),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_497),
.A2(n_10),
.B(n_11),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_498),
.B(n_496),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_499),
.A2(n_15),
.B(n_11),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_500),
.B(n_13),
.C(n_15),
.Y(n_501)
);

FAx1_ASAP7_75t_SL g502 ( 
.A(n_501),
.B(n_13),
.CI(n_486),
.CON(n_502),
.SN(n_502)
);


endmodule