module real_jpeg_27543_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_286, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_286;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_249;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_262;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_253;
wire n_273;
wire n_96;
wire n_269;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_SL g64 ( 
.A(n_0),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_1),
.Y(n_91)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_1),
.Y(n_93)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_1),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_4),
.A2(n_19),
.B1(n_20),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_4),
.A2(n_9),
.B1(n_27),
.B2(n_51),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_4),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_4),
.A2(n_42),
.B1(n_44),
.B2(n_51),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_6),
.A2(n_19),
.B1(n_20),
.B2(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_6),
.A2(n_9),
.B1(n_27),
.B2(n_29),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_6),
.A2(n_29),
.B1(n_42),
.B2(n_44),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_6),
.A2(n_29),
.B1(n_62),
.B2(n_63),
.Y(n_201)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_7),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_8),
.A2(n_19),
.B1(n_20),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_8),
.A2(n_9),
.B1(n_27),
.B2(n_36),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_SL g86 ( 
.A1(n_8),
.A2(n_9),
.B(n_25),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_8),
.A2(n_36),
.B1(n_62),
.B2(n_63),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_8),
.A2(n_36),
.B1(n_42),
.B2(n_44),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_8),
.B(n_26),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_SL g139 ( 
.A1(n_8),
.A2(n_10),
.B(n_42),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_8),
.A2(n_59),
.B(n_63),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_8),
.B(n_41),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_9),
.A2(n_10),
.B1(n_27),
.B2(n_43),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_9),
.A2(n_11),
.B1(n_21),
.B2(n_27),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_9),
.A2(n_36),
.B(n_138),
.C(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_10),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_11),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_11),
.A2(n_21),
.B1(n_62),
.B2(n_63),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_11),
.A2(n_21),
.B1(n_42),
.B2(n_44),
.Y(n_222)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

AOI21xp33_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_278),
.B(n_282),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_66),
.B(n_277),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_30),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_16),
.B(n_30),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_16),
.B(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_16),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_22),
.B1(n_26),
.B2(n_28),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_18),
.A2(n_33),
.B(n_34),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_20),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_20),
.A2(n_24),
.B(n_36),
.C(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_22),
.A2(n_26),
.B1(n_35),
.B2(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_22),
.B(n_26),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_26),
.Y(n_22)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_28),
.B(n_281),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_31),
.B(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_31),
.B(n_275),
.Y(n_276)
);

FAx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_37),
.CI(n_47),
.CON(n_31),
.SN(n_31)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_33),
.A2(n_34),
.B(n_50),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_35),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_36),
.A2(n_42),
.B(n_60),
.C(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_36),
.B(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_36),
.B(n_61),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_41),
.B1(n_45),
.B2(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_40),
.B(n_78),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_41),
.A2(n_53),
.B(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_44),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_45),
.B(n_79),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.C(n_54),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_75),
.B1(n_81),
.B2(n_82),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_48),
.B(n_82),
.C(n_83),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_48),
.A2(n_81),
.B1(n_97),
.B2(n_122),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_48),
.B(n_122),
.C(n_217),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_48),
.A2(n_81),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_52),
.A2(n_54),
.B1(n_256),
.B2(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_52),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_54),
.A2(n_253),
.B1(n_254),
.B2(n_256),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_54),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_65),
.Y(n_54)
);

INVxp33_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_61),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_57),
.B(n_102),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_57),
.A2(n_61),
.B1(n_102),
.B2(n_109),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_57),
.A2(n_61),
.B1(n_65),
.B2(n_222),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_61),
.A2(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_62),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_90),
.Y(n_89)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_274),
.B(n_276),
.Y(n_66)
);

OAI321xp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_248),
.A3(n_267),
.B1(n_272),
.B2(n_273),
.C(n_286),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_230),
.B(n_247),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_211),
.B(n_229),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_131),
.B(n_194),
.C(n_210),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_119),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_72),
.B(n_119),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_94),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_73),
.B(n_95),
.C(n_105),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_83),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_75),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_75),
.B(n_128),
.C(n_129),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_75),
.A2(n_82),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_75),
.A2(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_75),
.B(n_236),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_80),
.B(n_98),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_84),
.A2(n_85),
.B1(n_87),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_87),
.A2(n_126),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_87),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_87),
.B(n_178),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_87),
.B(n_153),
.C(n_165),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_88),
.A2(n_93),
.B(n_116),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_89),
.B(n_90),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_89),
.A2(n_93),
.B1(n_115),
.B2(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_104),
.B2(n_105),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.C(n_103),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_99),
.B1(n_100),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_97),
.A2(n_106),
.B1(n_107),
.B2(n_122),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_98),
.Y(n_255)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_103),
.A2(n_123),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_103),
.A2(n_123),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_103),
.A2(n_123),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_103),
.B(n_254),
.C(n_256),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_103),
.B(n_261),
.C(n_266),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_112),
.B2(n_113),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_106),
.A2(n_107),
.B1(n_160),
.B2(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_106),
.B(n_113),
.Y(n_204)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_122),
.C(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_107),
.B(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_110),
.B(n_111),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_111),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B(n_116),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_125),
.C(n_127),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_120),
.B(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_121),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_123),
.B(n_204),
.C(n_206),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_125),
.B(n_127),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_128),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_193),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_188),
.B(n_192),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_156),
.B(n_187),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_144),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_135),
.B(n_144),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_143),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_142),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_150),
.B2(n_151),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_145),
.B(n_153),
.C(n_154),
.Y(n_189)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_147),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_148),
.B(n_169),
.Y(n_180)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_152),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_153),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_155),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_153),
.A2(n_155),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_153),
.B(n_200),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_182),
.B(n_186),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_167),
.B(n_181),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_162),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_160),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_163),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_164),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_171),
.B(n_180),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_177),
.B(n_179),
.Y(n_171)
);

INVx5_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_184),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_190),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_195),
.B(n_196),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_208),
.B2(n_209),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_203),
.C(n_209),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_200),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_208),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_212),
.B(n_213),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_228),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_219),
.B2(n_220),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_220),
.C(n_228),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_221),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_225),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_224),
.A2(n_225),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_225),
.A2(n_239),
.B(n_241),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_232),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_245),
.B2(n_246),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_238),
.C(n_246),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_250),
.C(n_257),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_250),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_244),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_245),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_259),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_259),
.Y(n_273)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_257),
.A2(n_258),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_266),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_270),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_284),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);


endmodule