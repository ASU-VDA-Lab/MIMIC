module fake_jpeg_18423_n_186 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_6),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_38),
.Y(n_56)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_26),
.A2(n_20),
.B1(n_13),
.B2(n_19),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_45),
.B1(n_36),
.B2(n_20),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_23),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_59),
.B1(n_42),
.B2(n_33),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_12),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_58),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_61),
.B(n_15),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_19),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_13),
.B1(n_20),
.B2(n_18),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_22),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_47),
.B1(n_42),
.B2(n_51),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_65),
.Y(n_94)
);

OR2x4_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_44),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_72),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_33),
.B1(n_13),
.B2(n_42),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_33),
.B1(n_55),
.B2(n_51),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_44),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_46),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_77),
.C(n_61),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_47),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_17),
.B(n_18),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_0),
.B(n_1),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_59),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_93),
.B(n_15),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_82),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_76),
.B(n_17),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_40),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_40),
.Y(n_110)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_88),
.Y(n_98)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_76),
.B(n_11),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_67),
.B(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_103),
.Y(n_111)
);

AOI322xp5_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_74),
.A3(n_64),
.B1(n_78),
.B2(n_77),
.C1(n_68),
.C2(n_73),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_96),
.B(n_105),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_63),
.B1(n_64),
.B2(n_68),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_84),
.B1(n_91),
.B2(n_90),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_72),
.C(n_71),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_80),
.C(n_81),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_73),
.B(n_71),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_72),
.A3(n_62),
.B1(n_75),
.B2(n_14),
.C1(n_16),
.C2(n_38),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_108),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_14),
.B(n_1),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_110),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_101),
.C(n_99),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_115),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_82),
.B1(n_93),
.B2(n_86),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_0),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_86),
.B1(n_66),
.B2(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_84),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_124),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_39),
.B1(n_60),
.B2(n_44),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_100),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_14),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_106),
.B(n_7),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_130),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_95),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_107),
.B1(n_110),
.B2(n_103),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_134),
.Y(n_147)
);

AOI322xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_107),
.A3(n_108),
.B1(n_62),
.B2(n_98),
.C1(n_16),
.C2(n_6),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_133),
.B(n_135),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_16),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_119),
.B1(n_113),
.B2(n_3),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_139),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_132),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_145),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_123),
.B(n_111),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_142),
.A2(n_149),
.B(n_147),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_151),
.B1(n_114),
.B2(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_136),
.A2(n_111),
.B(n_113),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_129),
.C(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_154),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_114),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_7),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_149),
.C(n_147),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_160),
.C(n_140),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_142),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_140),
.C(n_124),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_164),
.B(n_5),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_163),
.C(n_165),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_157),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_145),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_6),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_158),
.B(n_7),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_168),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_5),
.Y(n_169)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_172),
.Y(n_178)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_8),
.B(n_9),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_166),
.A2(n_9),
.B(n_11),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_174),
.A2(n_9),
.B(n_11),
.Y(n_175)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_0),
.C(n_2),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_179),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_170),
.C(n_2),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g182 ( 
.A(n_177),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_182),
.A2(n_178),
.B(n_2),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_184),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_181),
.A2(n_3),
.B(n_180),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_3),
.Y(n_186)
);


endmodule