module real_jpeg_19290_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_11;
wire n_14;
wire n_7;
wire n_22;
wire n_18;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

AOI332xp33_ASAP7_75t_L g6 ( 
.A1(n_0),
.A2(n_2),
.A3(n_7),
.B1(n_13),
.B2(n_14),
.B3(n_17),
.C1(n_20),
.C2(n_22),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_1),
.A2(n_3),
.B1(n_11),
.B2(n_19),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

AO21x1_ASAP7_75t_L g14 ( 
.A1(n_2),
.A2(n_15),
.B(n_16),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_2),
.B(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

OAI21xp5_ASAP7_75t_SL g10 ( 
.A1(n_4),
.A2(n_11),
.B(n_12),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_4),
.B(n_11),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_8),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_10),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_9),
.B(n_10),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_18),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);


endmodule