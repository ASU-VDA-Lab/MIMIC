module real_jpeg_22587_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_0),
.A2(n_63),
.B1(n_64),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_0),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_0),
.A2(n_58),
.B1(n_67),
.B2(n_81),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_0),
.A2(n_36),
.B1(n_38),
.B2(n_81),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_0),
.A2(n_26),
.B1(n_28),
.B2(n_81),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_1),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_1),
.A2(n_26),
.B1(n_28),
.B2(n_37),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_2),
.A2(n_36),
.B1(n_38),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_2),
.A2(n_26),
.B1(n_28),
.B2(n_46),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_26),
.B1(n_28),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_4),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_4),
.A2(n_26),
.B1(n_28),
.B2(n_84),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_4),
.A2(n_36),
.B1(n_38),
.B2(n_84),
.Y(n_174)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_6),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_6),
.B(n_143),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_6),
.A2(n_160),
.B(n_184),
.Y(n_183)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_8),
.A2(n_36),
.B1(n_38),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_8),
.A2(n_54),
.B1(n_58),
.B2(n_67),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_8),
.A2(n_54),
.B1(n_63),
.B2(n_64),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_8),
.A2(n_26),
.B1(n_28),
.B2(n_54),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_10),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_11),
.A2(n_58),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_11),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_11),
.A2(n_62),
.B(n_64),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_11),
.B(n_70),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_11),
.A2(n_36),
.B(n_40),
.C(n_127),
.D(n_128),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_11),
.B(n_36),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_11),
.B(n_78),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_11),
.A2(n_24),
.B(n_142),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g175 ( 
.A1(n_11),
.A2(n_63),
.B(n_75),
.C(n_93),
.D(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_11),
.B(n_63),
.Y(n_176)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_12),
.Y(n_76)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_15),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_120),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_118),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_102),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_20),
.B(n_102),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_85),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_48),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B1(n_30),
.B2(n_32),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_24),
.A2(n_25),
.B1(n_27),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_24),
.A2(n_101),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_24),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_24),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_24),
.B(n_144),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_25),
.A2(n_149),
.B(n_159),
.Y(n_158)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_28),
.B1(n_41),
.B2(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_26),
.A2(n_42),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_28),
.B(n_41),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_28),
.B(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_45),
.B2(n_47),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_47),
.B(n_51),
.Y(n_50)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_36),
.A2(n_38),
.B1(n_76),
.B2(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_36),
.A2(n_176),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_41),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_38),
.B(n_79),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_39),
.A2(n_47),
.B1(n_139),
.B2(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_39),
.A2(n_174),
.B(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_52),
.Y(n_51)
);

CKINVDCx9p33_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_47),
.B(n_53),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_47),
.A2(n_51),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_47),
.B(n_66),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.C(n_72),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_49),
.A2(n_50),
.B1(n_72),
.B2(n_73),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_65),
.B(n_68),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_59),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_59),
.B(n_66),
.C(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_76),
.B(n_77),
.C(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_66),
.B(n_117),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_83),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_112),
.Y(n_111)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_77),
.Y(n_182)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_82),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_96),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_90),
.B1(n_91),
.B2(n_95),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_100),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.C(n_107),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_103),
.B(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_105),
.A2(n_107),
.B1(n_108),
.B2(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_105),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.C(n_114),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_109),
.A2(n_110),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_113),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_199),
.B(n_204),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_187),
.B(n_198),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_168),
.B(n_186),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_145),
.B(n_167),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_133),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_125),
.B(n_133),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_129),
.B1(n_130),
.B2(n_154),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_128),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_140),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_138),
.C(n_140),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_141),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_155),
.B(n_166),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_153),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_147),
.B(n_153),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_161),
.B(n_165),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_157),
.B(n_158),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_169),
.B(n_170),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_179),
.B2(n_185),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_173),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_175),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_178),
.C(n_185),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_179),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_183),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_188),
.B(n_189),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_195),
.C(n_196),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_191),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_200),
.B(n_201),
.Y(n_204)
);


endmodule