module real_jpeg_23181_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_3),
.A2(n_34),
.B1(n_45),
.B2(n_46),
.Y(n_100)
);

INVx8_ASAP7_75t_SL g61 ( 
.A(n_4),
.Y(n_61)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_5),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_5),
.B(n_120),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_110),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_5),
.A2(n_28),
.B(n_41),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_5),
.B(n_88),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_5),
.A2(n_25),
.B1(n_216),
.B2(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_5),
.A2(n_62),
.B(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_6),
.A2(n_67),
.B1(n_70),
.B2(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_6),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_6),
.A2(n_62),
.B1(n_63),
.B2(n_118),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_118),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_118),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_7),
.A2(n_38),
.B1(n_45),
.B2(n_46),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_7),
.A2(n_38),
.B1(n_62),
.B2(n_63),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_8),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_8),
.A2(n_62),
.B1(n_63),
.B2(n_74),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_74),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_74),
.Y(n_208)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_10),
.A2(n_67),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_77),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_77),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_77),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_48),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_13),
.A2(n_48),
.B1(n_62),
.B2(n_63),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_14),
.A2(n_62),
.B1(n_63),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_14),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_86),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_14),
.A2(n_86),
.B1(n_109),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_86),
.Y(n_156)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_15),
.Y(n_97)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_15),
.Y(n_125)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_15),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_146),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_145),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_122),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_20),
.B(n_122),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_21),
.B(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_21),
.B(n_150),
.Y(n_179)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_91),
.CI(n_101),
.CON(n_21),
.SN(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_54),
.B1(n_55),
.B2(n_90),
.Y(n_22)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_24),
.B(n_39),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_35),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_25),
.A2(n_125),
.B(n_126),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_25),
.A2(n_94),
.B(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_25),
.A2(n_97),
.B1(n_208),
.B2(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_25),
.A2(n_35),
.B(n_126),
.Y(n_244)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_26),
.B(n_37),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_26),
.A2(n_33),
.B1(n_96),
.B2(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_26),
.A2(n_36),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_28),
.B1(n_41),
.B2(n_43),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_27),
.B(n_223),
.Y(n_222)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_31),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_31),
.A2(n_93),
.B(n_115),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_44),
.B(n_49),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_40),
.A2(n_44),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_40),
.B(n_51),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_40),
.A2(n_99),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_40),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_40),
.B(n_110),
.Y(n_214)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_SL g192 ( 
.A1(n_43),
.A2(n_46),
.B(n_110),
.C(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_46),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_45),
.B(n_83),
.Y(n_243)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g242 ( 
.A1(n_46),
.A2(n_62),
.A3(n_82),
.B1(n_236),
.B2(n_243),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_52),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_52),
.A2(n_130),
.B(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_52),
.A2(n_191),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_52),
.A2(n_199),
.B1(n_200),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_78),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_56),
.B(n_78),
.C(n_90),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_71),
.B2(n_75),
.Y(n_56)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_57),
.A2(n_75),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_66),
.Y(n_57)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_70),
.Y(n_66)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_59),
.A2(n_63),
.A3(n_107),
.B1(n_108),
.B2(n_111),
.Y(n_106)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_62),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_63),
.B1(n_82),
.B2(n_83),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_63),
.B(n_110),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_70),
.A2(n_108),
.B(n_110),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_85),
.B(n_87),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_79),
.A2(n_81),
.B1(n_175),
.B2(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_80),
.B(n_89),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_80),
.A2(n_88),
.B1(n_103),
.B2(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_80),
.A2(n_88),
.B1(n_160),
.B2(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_85),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_81),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_98),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_98),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_95),
.Y(n_126)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_100),
.B(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_99),
.A2(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.C(n_116),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_116),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_105),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_112),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_106),
.A2(n_112),
.B1(n_113),
.B2(n_170),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_106),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_110),
.B(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_117),
.A2(n_119),
.B1(n_120),
.B2(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_138),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_122),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_132),
.CI(n_144),
.CON(n_122),
.SN(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_127),
.B1(n_128),
.B2(n_131),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_124),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_143),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_180),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_162),
.B(n_179),
.Y(n_148)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_149),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.C(n_161),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_152),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_154),
.B(n_161),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.C(n_159),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_159),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_156),
.B(n_199),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_168),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_163),
.B(n_166),
.Y(n_271)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.C(n_171),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_167),
.B(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_169),
.A2(n_171),
.B1(n_172),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_169),
.Y(n_268)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.C(n_177),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_173),
.B(n_253),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_254),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_176),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_270),
.C(n_271),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_264),
.B(n_269),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_248),
.B(n_263),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_229),
.B(n_247),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_204),
.B(n_228),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_194),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_186),
.B(n_194),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_192),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_187),
.A2(n_188),
.B1(n_192),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_192),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_202),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_201),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_201),
.C(n_202),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_203),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_212),
.B(n_227),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_206),
.B(n_210),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_217),
.B(n_226),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_214),
.B(n_215),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_221),
.Y(n_225)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_230),
.B(n_231),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_241),
.B1(n_245),
.B2(n_246),
.Y(n_231)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_232)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_237),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_240),
.C(n_245),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_238),
.Y(n_259)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_244),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_249),
.B(n_250),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_255),
.B2(n_256),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_258),
.C(n_261),
.Y(n_265)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_261),
.B2(n_262),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_257),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_258),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);


endmodule