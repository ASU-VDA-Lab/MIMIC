module fake_jpeg_31484_n_101 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_33),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_0),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_29),
.Y(n_51)
);

OR2x2_ASAP7_75t_SL g29 ( 
.A(n_18),
.B(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_2),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_32),
.Y(n_53)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_11),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_5),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_22),
.B(n_5),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_46),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_44),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_16),
.C(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_24),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_52),
.B(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_57),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_31),
.B1(n_34),
.B2(n_24),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_62),
.B(n_64),
.Y(n_74)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_49),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_53),
.B(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_42),
.B1(n_47),
.B2(n_26),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_39),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_26),
.B1(n_25),
.B2(n_10),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_44),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_51),
.C(n_53),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_72),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_70),
.A2(n_60),
.B1(n_64),
.B2(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_71),
.B(n_65),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_52),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_76),
.B(n_71),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_77),
.A2(n_70),
.B1(n_73),
.B2(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_81),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_57),
.B(n_45),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_43),
.B(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_84),
.B(n_86),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_85),
.A2(n_80),
.B1(n_9),
.B2(n_10),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_79),
.B(n_80),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_72),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_87),
.C(n_91),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_94),
.Y(n_98)
);

INVxp67_ASAP7_75t_SL g99 ( 
.A(n_98),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_96),
.B(n_7),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_9),
.Y(n_101)
);


endmodule