module fake_jpeg_7258_n_313 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_2),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_42),
.Y(n_50)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_16),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_25),
.B1(n_18),
.B2(n_23),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_47),
.A2(n_42),
.B1(n_38),
.B2(n_29),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_48),
.B(n_21),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_54),
.B(n_17),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_46),
.B1(n_25),
.B2(n_18),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_21),
.B1(n_19),
.B2(n_36),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_25),
.B(n_34),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_27),
.B(n_19),
.C(n_30),
.Y(n_91)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx2_ASAP7_75t_SL g100 ( 
.A(n_58),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_25),
.B1(n_33),
.B2(n_23),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_59),
.A2(n_60),
.B1(n_66),
.B2(n_70),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_23),
.B1(n_35),
.B2(n_34),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_62),
.Y(n_76)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_35),
.B1(n_28),
.B2(n_17),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_28),
.B1(n_35),
.B2(n_38),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_28),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_40),
.A2(n_35),
.B1(n_36),
.B2(n_34),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_72),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_17),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_74),
.B(n_83),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_32),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_91),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_28),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_SL g127 ( 
.A(n_84),
.B(n_109),
.C(n_27),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_95),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_48),
.B(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_93),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_92),
.B1(n_94),
.B2(n_51),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_29),
.B1(n_26),
.B2(n_36),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_65),
.Y(n_90)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_19),
.B1(n_26),
.B2(n_30),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_42),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_30),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_104),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_47),
.A2(n_68),
.B1(n_55),
.B2(n_72),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_103),
.B1(n_67),
.B2(n_27),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_51),
.A2(n_29),
.B1(n_26),
.B2(n_32),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_107),
.Y(n_139)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_1),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_3),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_110),
.B(n_49),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_3),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_112),
.B(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_118),
.B1(n_121),
.B2(n_124),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_32),
.B1(n_24),
.B2(n_27),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_24),
.B1(n_27),
.B2(n_6),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_127),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_24),
.B1(n_27),
.B2(n_6),
.Y(n_124)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_137),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_84),
.A2(n_16),
.B(n_5),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_131),
.A2(n_5),
.B(n_6),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_73),
.B(n_4),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_84),
.B(n_4),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_136),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_75),
.B(n_5),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_76),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_117),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_102),
.B1(n_98),
.B2(n_92),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_142),
.A2(n_149),
.B1(n_155),
.B2(n_132),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_139),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_143),
.B(n_144),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_139),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_120),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_145),
.Y(n_198)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_147),
.Y(n_177)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_99),
.B(n_88),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_148),
.A2(n_150),
.B(n_128),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_109),
.B1(n_95),
.B2(n_79),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_79),
.B(n_107),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_115),
.A2(n_87),
.B1(n_110),
.B2(n_80),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_151),
.A2(n_153),
.B1(n_10),
.B2(n_12),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_121),
.A2(n_87),
.B1(n_80),
.B2(n_103),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_112),
.A2(n_97),
.B1(n_77),
.B2(n_90),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_164),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_136),
.C(n_125),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_166),
.C(n_123),
.Y(n_174)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_158),
.A2(n_116),
.B1(n_105),
.B2(n_81),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_125),
.B(n_77),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_162),
.B(n_123),
.Y(n_176)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_161),
.Y(n_199)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_113),
.B(n_8),
.Y(n_166)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_172),
.Y(n_183)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_170),
.Y(n_200)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_173),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_188),
.Y(n_215)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_175),
.B(n_179),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_176),
.A2(n_178),
.B(n_184),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_118),
.B(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_159),
.A2(n_172),
.B1(n_142),
.B2(n_152),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_186),
.A2(n_189),
.B1(n_195),
.B2(n_201),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_132),
.C(n_128),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_192),
.C(n_162),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_149),
.B1(n_141),
.B2(n_148),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_8),
.Y(n_190)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_105),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_202),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_141),
.A2(n_116),
.B1(n_9),
.B2(n_10),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_146),
.A2(n_8),
.B(n_9),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_15),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_165),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_153),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_203),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_182),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_204),
.B(n_208),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_219),
.C(n_188),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_173),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_196),
.B(n_164),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_209),
.B(n_216),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_161),
.Y(n_211)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_171),
.Y(n_212)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_182),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_221),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_191),
.B(n_147),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_156),
.C(n_158),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_179),
.B(n_193),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_183),
.B(n_185),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_177),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_197),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_181),
.Y(n_225)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_226),
.A2(n_195),
.B1(n_186),
.B2(n_189),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_180),
.B(n_15),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_227),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_175),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_217),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_237),
.Y(n_261)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_232),
.A2(n_213),
.B(n_220),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_241),
.C(n_242),
.Y(n_251)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_207),
.A2(n_183),
.B1(n_201),
.B2(n_178),
.Y(n_239)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_223),
.A2(n_184),
.B1(n_207),
.B2(n_221),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_231),
.B1(n_229),
.B2(n_237),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_192),
.C(n_174),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_176),
.C(n_202),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_205),
.C(n_224),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_220),
.Y(n_248)
);

NAND4xp25_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_240),
.C(n_239),
.D(n_208),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_247),
.Y(n_252)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_241),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_232),
.B(n_224),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_255),
.B(n_257),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_230),
.B(n_177),
.CI(n_219),
.CON(n_256),
.SN(n_256)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_256),
.Y(n_271)
);

AOI322xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_223),
.A3(n_214),
.B1(n_204),
.B2(n_222),
.C1(n_210),
.C2(n_203),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_250),
.C(n_259),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_210),
.B1(n_214),
.B2(n_234),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_265),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_230),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_233),
.B1(n_236),
.B2(n_235),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_242),
.C(n_246),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_274),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_253),
.B(n_261),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_206),
.C(n_190),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_262),
.A2(n_226),
.B1(n_243),
.B2(n_238),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_275),
.A2(n_260),
.B1(n_266),
.B2(n_264),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_277),
.B(n_280),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_255),
.B(n_257),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_261),
.C(n_250),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_283),
.A2(n_291),
.B1(n_289),
.B2(n_290),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_284),
.A2(n_263),
.B1(n_272),
.B2(n_286),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_276),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_287),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_280),
.Y(n_287)
);

NOR3xp33_ASAP7_75t_SL g289 ( 
.A(n_271),
.B(n_256),
.C(n_252),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_278),
.B(n_273),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_256),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_279),
.C(n_272),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_291),
.A2(n_263),
.B(n_288),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_269),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_296),
.Y(n_303)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_282),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_297),
.A2(n_282),
.B1(n_294),
.B2(n_295),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_299),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_302),
.Y(n_308)
);

BUFx5_ASAP7_75t_L g302 ( 
.A(n_296),
.Y(n_302)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_302),
.B(n_303),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_300),
.B(n_308),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_305),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g309 ( 
.A(n_307),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_310),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_309),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_312),
.Y(n_313)
);


endmodule