module fake_jpeg_10225_n_261 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_261);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVxp67_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_23),
.Y(n_32)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_37),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_47),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_50),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_31),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_27),
.B1(n_14),
.B2(n_22),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_56),
.B1(n_68),
.B2(n_72),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_14),
.B1(n_37),
.B2(n_23),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_30),
.C(n_35),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_63),
.C(n_69),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_61),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_28),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_37),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_32),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_71),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_39),
.A2(n_14),
.B1(n_22),
.B2(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_37),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_32),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_39),
.A2(n_22),
.B1(n_35),
.B2(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_66),
.B(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_78),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_20),
.C(n_32),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_86),
.C(n_87),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_44),
.B1(n_32),
.B2(n_41),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_67),
.Y(n_101)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_83),
.Y(n_98)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

AOI22x1_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_91),
.B1(n_92),
.B2(n_43),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_41),
.C(n_44),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_20),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_57),
.A2(n_36),
.B1(n_34),
.B2(n_29),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_43),
.B1(n_46),
.B2(n_51),
.Y(n_97)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_70),
.A2(n_25),
.B1(n_26),
.B2(n_18),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_71),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_111),
.B1(n_109),
.B2(n_105),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_99),
.B1(n_113),
.B2(n_51),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_57),
.B1(n_65),
.B2(n_73),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_63),
.C(n_69),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_106),
.C(n_26),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_112),
.B(n_114),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_73),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_67),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_109),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_71),
.C(n_64),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_71),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_108),
.Y(n_130)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_41),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_70),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_88),
.A2(n_70),
.B1(n_34),
.B2(n_36),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_77),
.B(n_31),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_115),
.B(n_117),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_81),
.A3(n_88),
.B1(n_79),
.B2(n_76),
.Y(n_116)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_0),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_120),
.B(n_13),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_95),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_104),
.A2(n_85),
.B(n_82),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_125),
.B1(n_134),
.B2(n_31),
.Y(n_151)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_0),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_110),
.A2(n_91),
.B1(n_83),
.B2(n_18),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_129),
.B(n_136),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_46),
.B1(n_36),
.B2(n_34),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_132),
.B1(n_36),
.B2(n_34),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_112),
.B1(n_99),
.B2(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_29),
.Y(n_147)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_31),
.B(n_29),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_135),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_137),
.B(n_152),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_119),
.C(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_95),
.Y(n_141)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_145),
.Y(n_165)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_151),
.B1(n_156),
.B2(n_121),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_134),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_150),
.B(n_153),
.Y(n_173)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_134),
.Y(n_153)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_155),
.Y(n_161)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_21),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_157),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_15),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_124),
.B(n_31),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_154),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_29),
.C(n_4),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_130),
.B1(n_133),
.B2(n_116),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_163),
.A2(n_167),
.B1(n_168),
.B2(n_170),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_123),
.B1(n_118),
.B2(n_15),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_19),
.B1(n_21),
.B2(n_17),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_152),
.B(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_174),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_8),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_175),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_20),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_148),
.Y(n_183)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_180),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_143),
.A2(n_21),
.B1(n_0),
.B2(n_2),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_143),
.B1(n_147),
.B2(n_21),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_1),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_161),
.A2(n_156),
.B(n_139),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_181),
.A2(n_179),
.B(n_169),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_163),
.B(n_157),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_182),
.B(n_189),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_184),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_144),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_159),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_190),
.C(n_194),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_177),
.B1(n_169),
.B2(n_160),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_SL g189 ( 
.A(n_171),
.B(n_2),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_3),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_168),
.B(n_4),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_195),
.B(n_170),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_5),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_196),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_6),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_204),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_164),
.C(n_165),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_194),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_205),
.B(n_210),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_191),
.A2(n_179),
.B(n_171),
.Y(n_206)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_192),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_195),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_7),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_212),
.Y(n_218)
);

XOR2x2_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_182),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_213),
.A2(n_215),
.B(n_222),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_214),
.B(n_223),
.Y(n_231)
);

XOR2x2_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_183),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_188),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_8),
.B(n_9),
.Y(n_236)
);

NAND2x1_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_172),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_211),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_230),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_199),
.Y(n_228)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_207),
.C(n_200),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_235),
.C(n_9),
.Y(n_243)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_222),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_217),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_234),
.Y(n_239)
);

NOR2xp67_ASAP7_75t_SL g233 ( 
.A(n_215),
.B(n_213),
.Y(n_233)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_219),
.B(n_201),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_225),
.A2(n_200),
.B1(n_172),
.B2(n_207),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_236),
.B(n_216),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_237),
.B(n_242),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_236),
.B(n_221),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_10),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_10),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_244),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_239),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_246),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_240),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_247),
.B(n_250),
.Y(n_251)
);

BUFx24_ASAP7_75t_SL g252 ( 
.A(n_249),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_252),
.B(n_248),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_241),
.C(n_253),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_254),
.A2(n_255),
.B(n_238),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_256),
.A2(n_227),
.B(n_231),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_257),
.A2(n_10),
.B(n_11),
.Y(n_258)
);

OAI21x1_ASAP7_75t_L g259 ( 
.A1(n_258),
.A2(n_11),
.B(n_12),
.Y(n_259)
);

XNOR2x2_ASAP7_75t_SL g260 ( 
.A(n_259),
.B(n_11),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_29),
.Y(n_261)
);


endmodule