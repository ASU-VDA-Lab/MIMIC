module fake_netlist_6_3043_n_2778 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_762, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_783, n_106, n_725, n_358, n_160, n_751, n_449, n_131, n_749, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_442, n_480, n_142, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_739, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_768, n_38, n_471, n_289, n_421, n_781, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_727, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_748, n_506, n_56, n_763, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_666, n_371, n_770, n_567, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_752, n_112, n_172, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_734, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_779, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_366, n_777, n_407, n_450, n_103, n_272, n_526, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_745, n_654, n_323, n_606, n_393, n_411, n_503, n_716, n_152, n_623, n_92, n_599, n_513, n_776, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_731, n_406, n_483, n_735, n_102, n_204, n_482, n_755, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_714, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_767, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_775, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_759, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_85, n_99, n_257, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_743, n_766, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_728, n_681, n_729, n_110, n_151, n_774, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_722, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_736, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_778, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_2778);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_762;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_783;
input n_106;
input n_725;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_768;
input n_38;
input n_471;
input n_289;
input n_421;
input n_781;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_727;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_666;
input n_371;
input n_770;
input n_567;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_112;
input n_172;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_734;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_779;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_366;
input n_777;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_745;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_731;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_755;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_767;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_775;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_85;
input n_99;
input n_257;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_722;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_778;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_2778;

wire n_992;
wire n_2542;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_1027;
wire n_1351;
wire n_1189;
wire n_1212;
wire n_2157;
wire n_2332;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_822;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_1591;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_940;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_2603;
wire n_2660;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_1986;
wire n_2300;
wire n_2397;
wire n_824;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_966;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2009;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_2641;
wire n_1165;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_1214;
wire n_928;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2319;
wire n_2519;
wire n_825;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_890;
wire n_2377;
wire n_2178;
wire n_950;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_794;
wire n_2767;
wire n_894;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_2707;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_1139;
wire n_872;
wire n_1714;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_797;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2675;
wire n_1426;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_1992;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_1299;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_1475;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_931;
wire n_1021;
wire n_811;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_1314;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2596;
wire n_2274;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_2732;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_856;
wire n_2100;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_1129;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_1593;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_999;
wire n_1254;
wire n_2420;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_901;
wire n_1499;
wire n_2755;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_2154;
wire n_2727;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_1045;
wire n_1650;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_2671;
wire n_2761;
wire n_2715;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_2054;
wire n_876;
wire n_1337;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_1542;
wire n_2587;
wire n_875;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_933;
wire n_978;
wire n_2752;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_1379;
wire n_2528;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_2380;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_814;
wire n_2746;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_1461;
wire n_2076;
wire n_2736;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_971;
wire n_2702;
wire n_946;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_2743;
wire n_1973;
wire n_2267;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_1753;
wire n_2471;
wire n_2540;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_1170;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_2774;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_411),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_311),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_779),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_678),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_63),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_368),
.Y(n_792)
);

CKINVDCx14_ASAP7_75t_R g793 ( 
.A(n_160),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_442),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_328),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_786),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_752),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_749),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_103),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_81),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_775),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_491),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_469),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_195),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_573),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_680),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_760),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_776),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_220),
.Y(n_809)
);

BUFx10_ASAP7_75t_L g810 ( 
.A(n_210),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_579),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_780),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_683),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_355),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_369),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_371),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_269),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_728),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_295),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_710),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_662),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_422),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_707),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_151),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_305),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_54),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_105),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_709),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_515),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_552),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_150),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_50),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_663),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_222),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_697),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_571),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_374),
.Y(n_837)
);

BUFx10_ASAP7_75t_L g838 ( 
.A(n_536),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_670),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_411),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_51),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_14),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_730),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_320),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_260),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_647),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_119),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_484),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_783),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_785),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_283),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_368),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_684),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_67),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_690),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_674),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_10),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_691),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_657),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_425),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_638),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_774),
.Y(n_862)
);

CKINVDCx16_ASAP7_75t_R g863 ( 
.A(n_569),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_438),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_424),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_337),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_268),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_164),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_433),
.Y(n_869)
);

BUFx10_ASAP7_75t_L g870 ( 
.A(n_430),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_708),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_689),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_763),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_687),
.Y(n_874)
);

BUFx10_ASAP7_75t_L g875 ( 
.A(n_714),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_129),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_220),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_341),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_30),
.Y(n_879)
);

INVxp67_ASAP7_75t_SL g880 ( 
.A(n_751),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_331),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_527),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_19),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_38),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_68),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_174),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_267),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_623),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_731),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_247),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_711),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_727),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_695),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_765),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_77),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_692),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_437),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_729),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_90),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_773),
.Y(n_900)
);

BUFx8_ASAP7_75t_SL g901 ( 
.A(n_718),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_734),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_675),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_422),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_123),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_755),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_685),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_417),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_209),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_408),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_761),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_772),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_722),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_1),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_564),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_738),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_456),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_237),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_724),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_676),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_742),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_635),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_725),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_457),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_616),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_13),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_420),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_357),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_777),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_693),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_703),
.Y(n_931)
);

INVx1_ASAP7_75t_SL g932 ( 
.A(n_603),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_679),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_726),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_611),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_771),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_0),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_240),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_184),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_531),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_516),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_181),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_688),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_621),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_64),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_778),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_26),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_648),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_782),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_366),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_524),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_407),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_325),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_630),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_723),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_764),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_756),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_217),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_120),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_716),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_747),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_319),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_478),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_699),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_741),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_233),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_642),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_79),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_655),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_673),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_721),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_113),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_593),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_517),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_615),
.Y(n_975)
);

INVxp67_ASAP7_75t_SL g976 ( 
.A(n_211),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_32),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_404),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_104),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_694),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_658),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_704),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_720),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_318),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_125),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_715),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_509),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_353),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_496),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_372),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_219),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_767),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_768),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_245),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_543),
.Y(n_995)
);

BUFx5_ASAP7_75t_L g996 ( 
.A(n_370),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_576),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_712),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_705),
.Y(n_999)
);

BUFx2_ASAP7_75t_SL g1000 ( 
.A(n_654),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_348),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_757),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_417),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_125),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_682),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_745),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_748),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_563),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_386),
.Y(n_1009)
);

BUFx10_ASAP7_75t_L g1010 ( 
.A(n_733),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_78),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_39),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_633),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_73),
.Y(n_1014)
);

CKINVDCx14_ASAP7_75t_R g1015 ( 
.A(n_173),
.Y(n_1015)
);

BUFx8_ASAP7_75t_SL g1016 ( 
.A(n_567),
.Y(n_1016)
);

BUFx10_ASAP7_75t_L g1017 ( 
.A(n_604),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_440),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_744),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_58),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_278),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_739),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_617),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_459),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_48),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_753),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_681),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_736),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_637),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_396),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_408),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_354),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_737),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_732),
.Y(n_1034)
);

BUFx10_ASAP7_75t_L g1035 ( 
.A(n_784),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_6),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_341),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_455),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_769),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_672),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_696),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_627),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_700),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_388),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_319),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_762),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_15),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_750),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_698),
.Y(n_1049)
);

BUFx10_ASAP7_75t_L g1050 ( 
.A(n_465),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_601),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_110),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_701),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_420),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_754),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_187),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_646),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_781),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_81),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_493),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_520),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_252),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_544),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_702),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_48),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_76),
.Y(n_1066)
);

BUFx8_ASAP7_75t_SL g1067 ( 
.A(n_242),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_599),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_130),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_124),
.Y(n_1070)
);

CKINVDCx16_ASAP7_75t_R g1071 ( 
.A(n_127),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_429),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_713),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_61),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_528),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_126),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_468),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_581),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_300),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_62),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_447),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_758),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_717),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_759),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_329),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_525),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_37),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_106),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_155),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_212),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_176),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_719),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_36),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_0),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_59),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_511),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_746),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_735),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_743),
.Y(n_1099)
);

CKINVDCx14_ASAP7_75t_R g1100 ( 
.A(n_613),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_9),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_770),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_522),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_686),
.Y(n_1104)
);

INVx2_ASAP7_75t_SL g1105 ( 
.A(n_706),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_375),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_324),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_18),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_259),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_261),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_766),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_740),
.Y(n_1112)
);

CKINVDCx16_ASAP7_75t_R g1113 ( 
.A(n_677),
.Y(n_1113)
);

INVxp67_ASAP7_75t_SL g1114 ( 
.A(n_1110),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_901),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_996),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_798),
.Y(n_1117)
);

INVxp67_ASAP7_75t_SL g1118 ( 
.A(n_915),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_996),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_801),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_996),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_1016),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_1071),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_818),
.Y(n_1124)
);

INVxp33_ASAP7_75t_SL g1125 ( 
.A(n_787),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_850),
.Y(n_1126)
);

INVxp67_ASAP7_75t_SL g1127 ( 
.A(n_920),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_996),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_996),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_866),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_893),
.B(n_2),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_911),
.B(n_2),
.Y(n_1132)
);

INVxp67_ASAP7_75t_SL g1133 ( 
.A(n_943),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1110),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1110),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_892),
.Y(n_1136)
);

CKINVDCx16_ASAP7_75t_R g1137 ( 
.A(n_863),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1067),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_793),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_841),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_906),
.Y(n_1141)
);

CKINVDCx16_ASAP7_75t_R g1142 ( 
.A(n_1113),
.Y(n_1142)
);

INVxp67_ASAP7_75t_SL g1143 ( 
.A(n_944),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_1039),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_857),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_947),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_805),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1046),
.B(n_1015),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_917),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1012),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1101),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_791),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_804),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_838),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_814),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_817),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_806),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_825),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_807),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_907),
.Y(n_1160)
);

INVxp67_ASAP7_75t_SL g1161 ( 
.A(n_1043),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_821),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_827),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_828),
.Y(n_1164)
);

NOR2xp67_ASAP7_75t_L g1165 ( 
.A(n_840),
.B(n_1),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_1134),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_1135),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1114),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1147),
.B(n_1100),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1128),
.Y(n_1170)
);

OAI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1123),
.A2(n_937),
.B1(n_991),
.B2(n_881),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1116),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1114),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1119),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1139),
.B(n_1098),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1157),
.B(n_829),
.Y(n_1176)
);

AND3x2_ASAP7_75t_L g1177 ( 
.A(n_1148),
.B(n_976),
.C(n_951),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1152),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1121),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1153),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1154),
.B(n_932),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1129),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1159),
.B(n_1162),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1155),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1160),
.B(n_1034),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1156),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1158),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1164),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1140),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1163),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1145),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1146),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_1150),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_1151),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_1170),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1168),
.A2(n_1127),
.B1(n_1133),
.B2(n_1118),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1185),
.B(n_1161),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1174),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1173),
.B(n_1165),
.Y(n_1199)
);

BUFx4f_ASAP7_75t_L g1200 ( 
.A(n_1178),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1191),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1186),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1170),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1169),
.B(n_1176),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1191),
.Y(n_1205)
);

INVxp33_ASAP7_75t_L g1206 ( 
.A(n_1181),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1187),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1166),
.Y(n_1208)
);

CKINVDCx6p67_ASAP7_75t_R g1209 ( 
.A(n_1188),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1166),
.Y(n_1210)
);

INVx6_ASAP7_75t_L g1211 ( 
.A(n_1192),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1192),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1175),
.B(n_1137),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1172),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1179),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1182),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1178),
.Y(n_1217)
);

OR2x6_ASAP7_75t_L g1218 ( 
.A(n_1183),
.B(n_1130),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1171),
.B(n_1142),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1180),
.B(n_1125),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1193),
.B(n_1143),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1180),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1194),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1184),
.A2(n_1144),
.B1(n_1132),
.B2(n_1131),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1194),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1184),
.B(n_1115),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1190),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1190),
.B(n_1122),
.Y(n_1228)
);

NAND2xp33_ASAP7_75t_L g1229 ( 
.A(n_1189),
.B(n_803),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1177),
.A2(n_845),
.B1(n_847),
.B2(n_842),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1167),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1193),
.Y(n_1232)
);

INVx5_ASAP7_75t_L g1233 ( 
.A(n_1178),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1176),
.B(n_1138),
.Y(n_1234)
);

BUFx10_ASAP7_75t_L g1235 ( 
.A(n_1181),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1168),
.A2(n_868),
.B1(n_876),
.B2(n_867),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1181),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1181),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1168),
.B(n_1028),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1170),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1214),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1235),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1204),
.A2(n_1117),
.B1(n_1124),
.B2(n_1120),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1206),
.B(n_1237),
.Y(n_1244)
);

AND2x6_ASAP7_75t_SL g1245 ( 
.A(n_1218),
.B(n_1234),
.Y(n_1245)
);

AND2x2_ASAP7_75t_SL g1246 ( 
.A(n_1213),
.B(n_1126),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1197),
.B(n_1238),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1239),
.A2(n_1136),
.B1(n_1149),
.B2(n_1141),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1198),
.B(n_913),
.Y(n_1249)
);

INVx4_ASAP7_75t_L g1250 ( 
.A(n_1233),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1217),
.B(n_790),
.Y(n_1251)
);

INVxp33_ASAP7_75t_L g1252 ( 
.A(n_1219),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1216),
.Y(n_1253)
);

INVxp67_ASAP7_75t_L g1254 ( 
.A(n_1221),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1198),
.B(n_1215),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1215),
.B(n_1007),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1221),
.B(n_1064),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1202),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1199),
.B(n_1105),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1199),
.B(n_880),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1239),
.A2(n_1073),
.B1(n_1081),
.B2(n_1068),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1207),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1203),
.B(n_794),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1224),
.B(n_796),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1240),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1196),
.B(n_797),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1200),
.B(n_1103),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1233),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1218),
.B(n_802),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1240),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1236),
.A2(n_789),
.B1(n_830),
.B2(n_812),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1222),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1220),
.B(n_1030),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1195),
.B(n_808),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1233),
.B(n_1112),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1232),
.B(n_1059),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1208),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1227),
.B(n_788),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1231),
.B(n_811),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1209),
.B(n_1130),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1230),
.A2(n_916),
.B1(n_929),
.B2(n_882),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1210),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1201),
.B(n_810),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1223),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1225),
.B(n_820),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1205),
.B(n_1212),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1211),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1226),
.B(n_1099),
.Y(n_1288)
);

NOR3xp33_ASAP7_75t_L g1289 ( 
.A(n_1228),
.B(n_795),
.C(n_792),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1211),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1229),
.B(n_1104),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1202),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1211),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1204),
.B(n_823),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1202),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1202),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1204),
.A2(n_836),
.B(n_839),
.C(n_833),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1214),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1204),
.A2(n_890),
.B(n_897),
.C(n_887),
.Y(n_1299)
);

INVx4_ASAP7_75t_L g1300 ( 
.A(n_1233),
.Y(n_1300)
);

NAND2xp33_ASAP7_75t_L g1301 ( 
.A(n_1204),
.B(n_835),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1214),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1202),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_SL g1304 ( 
.A1(n_1206),
.A2(n_826),
.B1(n_844),
.B2(n_799),
.Y(n_1304)
);

AND2x6_ASAP7_75t_SL g1305 ( 
.A(n_1218),
.B(n_909),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1237),
.B(n_800),
.Y(n_1306)
);

INVxp67_ASAP7_75t_L g1307 ( 
.A(n_1237),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_1240),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1204),
.B(n_856),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1214),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1204),
.B(n_858),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1204),
.B(n_871),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1204),
.B(n_889),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1214),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1204),
.A2(n_846),
.B1(n_848),
.B2(n_843),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1204),
.B(n_896),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1204),
.B(n_809),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1204),
.B(n_900),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1214),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1235),
.Y(n_1320)
);

OAI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1204),
.A2(n_992),
.B1(n_1082),
.B2(n_974),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1204),
.B(n_903),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1214),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1204),
.B(n_815),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1202),
.Y(n_1325)
);

AOI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1204),
.A2(n_853),
.B1(n_855),
.B2(n_849),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1237),
.B(n_1102),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1206),
.B(n_810),
.Y(n_1328)
);

AO22x2_ASAP7_75t_L g1329 ( 
.A1(n_1219),
.A2(n_942),
.B1(n_958),
.B2(n_945),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1240),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1202),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1204),
.B(n_816),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1204),
.B(n_933),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1204),
.B(n_819),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1240),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1204),
.A2(n_956),
.B1(n_965),
.B2(n_946),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1204),
.B(n_822),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1237),
.B(n_1096),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1202),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1204),
.B(n_960),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1206),
.B(n_870),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1202),
.Y(n_1342)
);

INVx4_ASAP7_75t_L g1343 ( 
.A(n_1233),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1255),
.A2(n_975),
.B(n_969),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1336),
.A2(n_1266),
.B(n_1309),
.C(n_1294),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1317),
.B(n_1337),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1324),
.A2(n_1002),
.B1(n_1006),
.B2(n_989),
.Y(n_1347)
);

OAI321xp33_ASAP7_75t_L g1348 ( 
.A1(n_1321),
.A2(n_1334),
.A3(n_1332),
.B1(n_1264),
.B2(n_1273),
.C(n_1261),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1330),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1258),
.Y(n_1350)
);

O2A1O1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1311),
.A2(n_1022),
.B(n_1023),
.C(n_1019),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1260),
.A2(n_1029),
.B(n_1027),
.Y(n_1352)
);

OAI21xp33_ASAP7_75t_L g1353 ( 
.A1(n_1247),
.A2(n_831),
.B(n_824),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1280),
.B(n_870),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1312),
.A2(n_1061),
.B(n_1053),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1329),
.A2(n_1340),
.B1(n_1333),
.B2(n_1316),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1313),
.B(n_1075),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1318),
.A2(n_1083),
.B(n_1077),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1241),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1322),
.B(n_1092),
.Y(n_1360)
);

NOR2xp67_ASAP7_75t_L g1361 ( 
.A(n_1307),
.B(n_859),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1262),
.B(n_1097),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1252),
.B(n_854),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1292),
.B(n_861),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1259),
.A2(n_813),
.B(n_803),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1254),
.B(n_862),
.Y(n_1366)
);

AOI21xp33_ASAP7_75t_L g1367 ( 
.A1(n_1301),
.A2(n_834),
.B(n_832),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1257),
.A2(n_1342),
.B(n_1296),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1295),
.B(n_872),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1330),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1315),
.B(n_1326),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1297),
.A2(n_962),
.B(n_1018),
.C(n_959),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1253),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1303),
.A2(n_813),
.B(n_803),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1325),
.B(n_873),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1331),
.B(n_874),
.Y(n_1376)
);

NAND2x1p5_ASAP7_75t_L g1377 ( 
.A(n_1335),
.B(n_813),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1339),
.Y(n_1378)
);

AOI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1249),
.A2(n_1044),
.B(n_1032),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1286),
.A2(n_1078),
.B(n_999),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1276),
.B(n_888),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1298),
.B(n_891),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1302),
.B(n_894),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1310),
.A2(n_1078),
.B(n_999),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1314),
.A2(n_1078),
.B(n_999),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1319),
.A2(n_902),
.B(n_898),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1323),
.B(n_1256),
.Y(n_1387)
);

AOI21xp33_ASAP7_75t_L g1388 ( 
.A1(n_1306),
.A2(n_851),
.B(n_837),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1279),
.B(n_1244),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1251),
.Y(n_1390)
);

A2O1A1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1299),
.A2(n_1047),
.B(n_1062),
.C(n_1045),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1272),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1327),
.A2(n_919),
.B(n_912),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1251),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1338),
.A2(n_922),
.B(n_921),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1329),
.B(n_923),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1277),
.A2(n_925),
.B(n_924),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1274),
.A2(n_931),
.B(n_930),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1285),
.A2(n_935),
.B(n_934),
.Y(n_1399)
);

INVx4_ASAP7_75t_L g1400 ( 
.A(n_1335),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1282),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1246),
.B(n_1243),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1328),
.B(n_852),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1263),
.A2(n_940),
.B(n_936),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1341),
.B(n_941),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_SL g1406 ( 
.A(n_1284),
.B(n_948),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_1248),
.B(n_949),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1308),
.A2(n_955),
.B(n_954),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1265),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1269),
.B(n_957),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1304),
.B(n_879),
.Y(n_1411)
);

A2O1A1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1278),
.A2(n_1085),
.B(n_1088),
.C(n_1079),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1288),
.A2(n_1094),
.B(n_1095),
.C(n_1091),
.Y(n_1413)
);

INVx2_ASAP7_75t_SL g1414 ( 
.A(n_1283),
.Y(n_1414)
);

OR2x6_ASAP7_75t_L g1415 ( 
.A(n_1242),
.B(n_1000),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1270),
.Y(n_1416)
);

AO21x1_ASAP7_75t_L g1417 ( 
.A1(n_1267),
.A2(n_1107),
.B(n_3),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1320),
.B(n_860),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1287),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1289),
.B(n_961),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1281),
.A2(n_1271),
.B(n_1275),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1290),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1250),
.B(n_963),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1291),
.A2(n_967),
.B(n_964),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1293),
.A2(n_971),
.B1(n_973),
.B2(n_970),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1268),
.Y(n_1426)
);

AO21x1_ASAP7_75t_L g1427 ( 
.A1(n_1300),
.A2(n_3),
.B(n_4),
.Y(n_1427)
);

CKINVDCx10_ASAP7_75t_R g1428 ( 
.A(n_1305),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1343),
.B(n_980),
.Y(n_1429)
);

NOR2x2_ASAP7_75t_L g1430 ( 
.A(n_1245),
.B(n_905),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1317),
.B(n_981),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1317),
.B(n_982),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1317),
.B(n_983),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1255),
.A2(n_987),
.B(n_986),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1317),
.B(n_950),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1255),
.A2(n_995),
.B(n_993),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1255),
.A2(n_998),
.B(n_997),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1241),
.Y(n_1438)
);

OAI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1294),
.A2(n_1008),
.B(n_1005),
.Y(n_1439)
);

INVxp67_ASAP7_75t_L g1440 ( 
.A(n_1276),
.Y(n_1440)
);

INVx4_ASAP7_75t_L g1441 ( 
.A(n_1330),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1317),
.B(n_984),
.Y(n_1442)
);

A2O1A1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1317),
.A2(n_1024),
.B(n_1026),
.C(n_1013),
.Y(n_1443)
);

AOI21xp33_ASAP7_75t_L g1444 ( 
.A1(n_1317),
.A2(n_865),
.B(n_864),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1317),
.B(n_1033),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1258),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1294),
.A2(n_1040),
.B(n_1038),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1317),
.B(n_1041),
.Y(n_1448)
);

AOI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1255),
.A2(n_1048),
.B(n_1042),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1241),
.Y(n_1450)
);

BUFx10_ASAP7_75t_L g1451 ( 
.A(n_1245),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1258),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1317),
.B(n_1049),
.Y(n_1453)
);

NOR2x1_ASAP7_75t_R g1454 ( 
.A(n_1280),
.B(n_869),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1317),
.B(n_1051),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1255),
.A2(n_1057),
.B(n_1055),
.Y(n_1456)
);

O2A1O1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1336),
.A2(n_1021),
.B(n_1056),
.C(n_985),
.Y(n_1457)
);

BUFx4f_ASAP7_75t_L g1458 ( 
.A(n_1330),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1258),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1258),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1241),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1254),
.B(n_1058),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1276),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1317),
.B(n_1060),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1255),
.A2(n_1084),
.B(n_1063),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1317),
.B(n_1086),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1255),
.A2(n_1111),
.B(n_878),
.Y(n_1467)
);

AO21x1_ASAP7_75t_L g1468 ( 
.A1(n_1336),
.A2(n_4),
.B(n_5),
.Y(n_1468)
);

AO21x2_ASAP7_75t_L g1469 ( 
.A1(n_1294),
.A2(n_443),
.B(n_441),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1276),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1317),
.B(n_877),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1255),
.A2(n_884),
.B(n_883),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1258),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1294),
.A2(n_1108),
.B(n_1106),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1255),
.A2(n_886),
.B(n_885),
.Y(n_1475)
);

OAI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1294),
.A2(n_1054),
.B(n_1052),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1255),
.A2(n_899),
.B(n_895),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1258),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1317),
.B(n_904),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1258),
.Y(n_1480)
);

AO21x1_ASAP7_75t_L g1481 ( 
.A1(n_1336),
.A2(n_5),
.B(n_6),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1317),
.A2(n_875),
.B1(n_1010),
.B2(n_838),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1330),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1294),
.A2(n_1080),
.B(n_1076),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1258),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1280),
.Y(n_1486)
);

BUFx12f_ASAP7_75t_L g1487 ( 
.A(n_1305),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1254),
.Y(n_1488)
);

BUFx4f_ASAP7_75t_SL g1489 ( 
.A(n_1246),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1255),
.A2(n_910),
.B(n_908),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1254),
.B(n_875),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1317),
.B(n_914),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1330),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1258),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1255),
.A2(n_926),
.B(n_918),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1346),
.B(n_927),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1345),
.A2(n_445),
.B(n_444),
.Y(n_1497)
);

A2O1A1Ixp33_ASAP7_75t_L g1498 ( 
.A1(n_1435),
.A2(n_938),
.B(n_939),
.C(n_928),
.Y(n_1498)
);

NOR3xp33_ASAP7_75t_L g1499 ( 
.A(n_1442),
.B(n_953),
.C(n_952),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1349),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1359),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1371),
.A2(n_448),
.B(n_446),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1356),
.A2(n_1432),
.B1(n_1433),
.B2(n_1431),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1350),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1373),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1387),
.A2(n_450),
.B(n_449),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1378),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1348),
.B(n_1010),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1400),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1411),
.A2(n_1035),
.B1(n_1050),
.B2(n_1017),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1445),
.A2(n_968),
.B1(n_972),
.B2(n_966),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1489),
.Y(n_1512)
);

NAND2xp33_ASAP7_75t_SL g1513 ( 
.A(n_1349),
.B(n_977),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1458),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1446),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1449),
.A2(n_1368),
.B(n_1362),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1389),
.A2(n_452),
.B(n_451),
.Y(n_1517)
);

O2A1O1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1444),
.A2(n_1035),
.B(n_1050),
.C(n_1017),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1349),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1448),
.A2(n_1455),
.B(n_1453),
.Y(n_1520)
);

O2A1O1Ixp5_ASAP7_75t_L g1521 ( 
.A1(n_1464),
.A2(n_454),
.B(n_458),
.C(n_453),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1440),
.B(n_978),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1466),
.A2(n_1421),
.B(n_1366),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1462),
.A2(n_461),
.B(n_460),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_SL g1525 ( 
.A1(n_1474),
.A2(n_1484),
.B(n_1476),
.C(n_1479),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1370),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1463),
.B(n_979),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1382),
.A2(n_1383),
.B(n_1360),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1470),
.B(n_988),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1452),
.A2(n_994),
.B1(n_1001),
.B2(n_990),
.Y(n_1530)
);

AOI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1402),
.A2(n_1004),
.B1(n_1009),
.B2(n_1003),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1357),
.A2(n_463),
.B(n_462),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1471),
.B(n_1011),
.Y(n_1533)
);

O2A1O1Ixp33_ASAP7_75t_SL g1534 ( 
.A1(n_1443),
.A2(n_466),
.B(n_467),
.C(n_464),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1441),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1414),
.B(n_1014),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1492),
.B(n_1020),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1459),
.B(n_1025),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1364),
.A2(n_471),
.B(n_470),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1438),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1460),
.B(n_1031),
.Y(n_1541)
);

A2O1A1Ixp33_ASAP7_75t_L g1542 ( 
.A1(n_1457),
.A2(n_1037),
.B(n_1065),
.C(n_1036),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1473),
.A2(n_1069),
.B1(n_1070),
.B2(n_1066),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1363),
.B(n_1072),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1441),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1478),
.A2(n_1087),
.B1(n_1089),
.B2(n_1074),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1369),
.A2(n_1376),
.B(n_1375),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1480),
.A2(n_1093),
.B1(n_1109),
.B2(n_1090),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1450),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_SL g1550 ( 
.A(n_1486),
.B(n_472),
.Y(n_1550)
);

CKINVDCx6p67_ASAP7_75t_R g1551 ( 
.A(n_1415),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1485),
.B(n_1494),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1403),
.B(n_7),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1405),
.B(n_7),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1488),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1461),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1483),
.Y(n_1557)
);

O2A1O1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1367),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_1558)
);

AO32x1_ASAP7_75t_L g1559 ( 
.A1(n_1401),
.A2(n_12),
.A3(n_8),
.B1(n_11),
.B2(n_13),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1493),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1392),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1381),
.B(n_11),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1416),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1353),
.B(n_12),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1390),
.A2(n_474),
.B(n_473),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1394),
.A2(n_476),
.B(n_475),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1409),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1439),
.B(n_14),
.Y(n_1568)
);

OAI22x1_ASAP7_75t_L g1569 ( 
.A1(n_1491),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1569)
);

AOI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1344),
.A2(n_479),
.B(n_477),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1419),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1422),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1347),
.A2(n_481),
.B1(n_482),
.B2(n_480),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1410),
.A2(n_485),
.B1(n_486),
.B2(n_483),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1447),
.B(n_16),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1482),
.A2(n_1396),
.B1(n_1361),
.B2(n_1426),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1379),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1352),
.A2(n_488),
.B(n_487),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1469),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1354),
.B(n_17),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1495),
.B(n_18),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1472),
.B(n_19),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1388),
.B(n_20),
.Y(n_1583)
);

BUFx4f_ASAP7_75t_L g1584 ( 
.A(n_1487),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1407),
.B(n_20),
.Y(n_1585)
);

INVx5_ASAP7_75t_L g1586 ( 
.A(n_1415),
.Y(n_1586)
);

O2A1O1Ixp33_ASAP7_75t_L g1587 ( 
.A1(n_1412),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_1587)
);

AOI222xp33_ASAP7_75t_L g1588 ( 
.A1(n_1454),
.A2(n_23),
.B1(n_25),
.B2(n_21),
.C1(n_22),
.C2(n_24),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1467),
.B(n_1475),
.Y(n_1589)
);

BUFx4f_ASAP7_75t_SL g1590 ( 
.A(n_1451),
.Y(n_1590)
);

A2O1A1Ixp33_ASAP7_75t_L g1591 ( 
.A1(n_1477),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1418),
.B(n_27),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1490),
.B(n_27),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1406),
.A2(n_490),
.B(n_489),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1417),
.Y(n_1595)
);

O2A1O1Ixp5_ASAP7_75t_SL g1596 ( 
.A1(n_1420),
.A2(n_1429),
.B(n_1481),
.C(n_1468),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1434),
.B(n_28),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1436),
.B(n_28),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1423),
.A2(n_494),
.B1(n_495),
.B2(n_492),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1437),
.B(n_29),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1377),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1456),
.B(n_29),
.Y(n_1602)
);

A2O1A1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1355),
.A2(n_1358),
.B(n_1413),
.C(n_1351),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1425),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1430),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1427),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1386),
.A2(n_498),
.B(n_497),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1391),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_L g1609 ( 
.A(n_1451),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1372),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1465),
.B(n_30),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1365),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1408),
.A2(n_500),
.B1(n_501),
.B2(n_499),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1398),
.B(n_31),
.Y(n_1614)
);

AO31x2_ASAP7_75t_L g1615 ( 
.A1(n_1579),
.A2(n_1380),
.A3(n_1374),
.B(n_1384),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1552),
.A2(n_1393),
.B1(n_1395),
.B2(n_1399),
.Y(n_1616)
);

NAND3xp33_ASAP7_75t_SL g1617 ( 
.A(n_1510),
.B(n_1404),
.C(n_1424),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1514),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1555),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1504),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1496),
.B(n_1397),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1507),
.Y(n_1622)
);

NAND3xp33_ASAP7_75t_SL g1623 ( 
.A(n_1499),
.B(n_1428),
.C(n_1385),
.Y(n_1623)
);

A2O1A1Ixp33_ASAP7_75t_L g1624 ( 
.A1(n_1525),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1544),
.B(n_33),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1519),
.Y(n_1626)
);

A2O1A1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1583),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1503),
.A2(n_503),
.B(n_502),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1533),
.B(n_34),
.Y(n_1629)
);

OAI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1523),
.A2(n_505),
.B(n_504),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1537),
.B(n_1515),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1529),
.B(n_35),
.Y(n_1632)
);

INVxp67_ASAP7_75t_SL g1633 ( 
.A(n_1560),
.Y(n_1633)
);

AO31x2_ASAP7_75t_L g1634 ( 
.A1(n_1497),
.A2(n_507),
.A3(n_508),
.B(n_506),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1500),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1520),
.A2(n_512),
.B(n_510),
.Y(n_1636)
);

A2O1A1Ixp33_ASAP7_75t_L g1637 ( 
.A1(n_1568),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1547),
.A2(n_514),
.B(n_513),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1526),
.Y(n_1639)
);

AOI211x1_ASAP7_75t_L g1640 ( 
.A1(n_1575),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_1640)
);

INVx2_ASAP7_75t_SL g1641 ( 
.A(n_1557),
.Y(n_1641)
);

A2O1A1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1585),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_1642)
);

AOI221xp5_ASAP7_75t_SL g1643 ( 
.A1(n_1518),
.A2(n_1542),
.B1(n_1508),
.B2(n_1498),
.C(n_1511),
.Y(n_1643)
);

O2A1O1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1592),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1528),
.A2(n_519),
.B(n_518),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1527),
.B(n_43),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_1557),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1572),
.Y(n_1648)
);

OAI21x1_ASAP7_75t_L g1649 ( 
.A1(n_1516),
.A2(n_523),
.B(n_521),
.Y(n_1649)
);

NOR2x1_ASAP7_75t_R g1650 ( 
.A(n_1586),
.B(n_526),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1589),
.A2(n_530),
.B(n_529),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1554),
.B(n_1553),
.Y(n_1652)
);

O2A1O1Ixp33_ASAP7_75t_L g1653 ( 
.A1(n_1580),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1501),
.Y(n_1654)
);

OAI21x1_ASAP7_75t_L g1655 ( 
.A1(n_1612),
.A2(n_533),
.B(n_532),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1604),
.B(n_46),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1578),
.A2(n_535),
.B(n_534),
.Y(n_1657)
);

OAI22x1_ASAP7_75t_L g1658 ( 
.A1(n_1606),
.A2(n_50),
.B1(n_51),
.B2(n_49),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1500),
.Y(n_1659)
);

OAI21xp33_ASAP7_75t_L g1660 ( 
.A1(n_1531),
.A2(n_47),
.B(n_49),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1567),
.Y(n_1661)
);

OR2x6_ASAP7_75t_L g1662 ( 
.A(n_1535),
.B(n_537),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1505),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1603),
.A2(n_539),
.B(n_538),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1540),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1538),
.B(n_47),
.Y(n_1666)
);

AOI211x1_ASAP7_75t_L g1667 ( 
.A1(n_1564),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1549),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1576),
.A2(n_541),
.B(n_540),
.Y(n_1669)
);

OAI21x1_ASAP7_75t_L g1670 ( 
.A1(n_1570),
.A2(n_545),
.B(n_542),
.Y(n_1670)
);

AO31x2_ASAP7_75t_L g1671 ( 
.A1(n_1577),
.A2(n_547),
.A3(n_548),
.B(n_546),
.Y(n_1671)
);

AO31x2_ASAP7_75t_L g1672 ( 
.A1(n_1595),
.A2(n_550),
.A3(n_551),
.B(n_549),
.Y(n_1672)
);

CKINVDCx11_ASAP7_75t_R g1673 ( 
.A(n_1609),
.Y(n_1673)
);

CKINVDCx20_ASAP7_75t_R g1674 ( 
.A(n_1512),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1556),
.B(n_52),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1561),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1593),
.A2(n_56),
.B1(n_53),
.B2(n_55),
.Y(n_1677)
);

OAI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1596),
.A2(n_554),
.B(n_553),
.Y(n_1678)
);

NOR4xp25_ASAP7_75t_L g1679 ( 
.A(n_1558),
.B(n_57),
.C(n_55),
.D(n_56),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1545),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1541),
.B(n_57),
.Y(n_1681)
);

AOI221xp5_ASAP7_75t_SL g1682 ( 
.A1(n_1569),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.C(n_61),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1571),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1502),
.A2(n_556),
.B(n_555),
.Y(n_1684)
);

A2O1A1Ixp33_ASAP7_75t_L g1685 ( 
.A1(n_1562),
.A2(n_63),
.B(n_60),
.C(n_62),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1522),
.B(n_64),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1509),
.B(n_557),
.Y(n_1687)
);

NAND2xp33_ASAP7_75t_SL g1688 ( 
.A(n_1609),
.B(n_65),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1563),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1689)
);

NOR2xp67_ASAP7_75t_L g1690 ( 
.A(n_1586),
.B(n_558),
.Y(n_1690)
);

O2A1O1Ixp33_ASAP7_75t_SL g1691 ( 
.A1(n_1591),
.A2(n_560),
.B(n_561),
.C(n_559),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1607),
.A2(n_565),
.B(n_562),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1608),
.A2(n_69),
.B1(n_66),
.B2(n_68),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1517),
.A2(n_568),
.B(n_566),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1610),
.Y(n_1695)
);

INVx5_ASAP7_75t_L g1696 ( 
.A(n_1609),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_1586),
.Y(n_1697)
);

CKINVDCx20_ASAP7_75t_R g1698 ( 
.A(n_1590),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1536),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1581),
.B(n_70),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1539),
.A2(n_1506),
.B(n_1534),
.Y(n_1701)
);

OR2x6_ASAP7_75t_L g1702 ( 
.A(n_1605),
.B(n_570),
.Y(n_1702)
);

NOR2xp67_ASAP7_75t_L g1703 ( 
.A(n_1601),
.B(n_572),
.Y(n_1703)
);

O2A1O1Ixp33_ASAP7_75t_SL g1704 ( 
.A1(n_1597),
.A2(n_575),
.B(n_577),
.C(n_574),
.Y(n_1704)
);

AO31x2_ASAP7_75t_L g1705 ( 
.A1(n_1599),
.A2(n_580),
.A3(n_582),
.B(n_578),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1582),
.B(n_583),
.Y(n_1706)
);

INVx4_ASAP7_75t_L g1707 ( 
.A(n_1551),
.Y(n_1707)
);

AO21x1_ASAP7_75t_L g1708 ( 
.A1(n_1598),
.A2(n_73),
.B(n_72),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1600),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1602),
.A2(n_74),
.B1(n_71),
.B2(n_72),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1588),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1611),
.Y(n_1712)
);

AO32x2_ASAP7_75t_L g1713 ( 
.A1(n_1530),
.A2(n_78),
.A3(n_75),
.B1(n_77),
.B2(n_79),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1543),
.B(n_80),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1546),
.B(n_80),
.Y(n_1715)
);

OAI21x1_ASAP7_75t_L g1716 ( 
.A1(n_1521),
.A2(n_585),
.B(n_584),
.Y(n_1716)
);

OAI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1614),
.A2(n_587),
.B(n_586),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1513),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_1718)
);

OAI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1565),
.A2(n_589),
.B(n_588),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1548),
.B(n_82),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1574),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_1721)
);

AOI21x1_ASAP7_75t_L g1722 ( 
.A1(n_1566),
.A2(n_1532),
.B(n_1524),
.Y(n_1722)
);

O2A1O1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1587),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1594),
.A2(n_1613),
.B(n_1573),
.Y(n_1724)
);

BUFx3_ASAP7_75t_L g1725 ( 
.A(n_1584),
.Y(n_1725)
);

AOI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1550),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.C(n_89),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1559),
.A2(n_591),
.B(n_590),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1559),
.A2(n_594),
.B(n_592),
.Y(n_1728)
);

OAI21x1_ASAP7_75t_L g1729 ( 
.A1(n_1516),
.A2(n_596),
.B(n_595),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1496),
.B(n_88),
.Y(n_1730)
);

CKINVDCx8_ASAP7_75t_R g1731 ( 
.A(n_1609),
.Y(n_1731)
);

BUFx2_ASAP7_75t_L g1732 ( 
.A(n_1514),
.Y(n_1732)
);

BUFx10_ASAP7_75t_L g1733 ( 
.A(n_1609),
.Y(n_1733)
);

AOI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1520),
.A2(n_598),
.B(n_597),
.Y(n_1734)
);

OA21x2_ASAP7_75t_L g1735 ( 
.A1(n_1579),
.A2(n_602),
.B(n_600),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1504),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1520),
.A2(n_606),
.B(n_605),
.Y(n_1737)
);

BUFx8_ASAP7_75t_L g1738 ( 
.A(n_1609),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1496),
.B(n_89),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1520),
.A2(n_608),
.B(n_607),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1496),
.B(n_90),
.Y(n_1741)
);

OAI21x1_ASAP7_75t_L g1742 ( 
.A1(n_1516),
.A2(n_610),
.B(n_609),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1544),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_1743)
);

AO31x2_ASAP7_75t_L g1744 ( 
.A1(n_1579),
.A2(n_614),
.A3(n_618),
.B(n_612),
.Y(n_1744)
);

OAI21x1_ASAP7_75t_L g1745 ( 
.A1(n_1516),
.A2(n_620),
.B(n_619),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1504),
.Y(n_1746)
);

BUFx8_ASAP7_75t_L g1747 ( 
.A(n_1609),
.Y(n_1747)
);

OR2x6_ASAP7_75t_L g1748 ( 
.A(n_1514),
.B(n_622),
.Y(n_1748)
);

OAI21x1_ASAP7_75t_L g1749 ( 
.A1(n_1516),
.A2(n_625),
.B(n_624),
.Y(n_1749)
);

AOI221x1_ASAP7_75t_L g1750 ( 
.A1(n_1503),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.C(n_94),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1504),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1555),
.B(n_94),
.Y(n_1752)
);

CKINVDCx11_ASAP7_75t_R g1753 ( 
.A(n_1698),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1711),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_1754)
);

INVx4_ASAP7_75t_L g1755 ( 
.A(n_1696),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1625),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1631),
.B(n_1709),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1652),
.A2(n_1632),
.B1(n_1633),
.B2(n_1712),
.Y(n_1758)
);

INVx4_ASAP7_75t_L g1759 ( 
.A(n_1696),
.Y(n_1759)
);

CKINVDCx11_ASAP7_75t_R g1760 ( 
.A(n_1673),
.Y(n_1760)
);

BUFx4f_ASAP7_75t_SL g1761 ( 
.A(n_1674),
.Y(n_1761)
);

OAI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1743),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1660),
.A2(n_1686),
.B1(n_1721),
.B2(n_1628),
.Y(n_1763)
);

OAI21xp5_ASAP7_75t_SL g1764 ( 
.A1(n_1677),
.A2(n_100),
.B(n_99),
.Y(n_1764)
);

CKINVDCx11_ASAP7_75t_R g1765 ( 
.A(n_1731),
.Y(n_1765)
);

BUFx3_ASAP7_75t_L g1766 ( 
.A(n_1639),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1619),
.A2(n_1695),
.B1(n_1739),
.B2(n_1730),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1746),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1620),
.Y(n_1769)
);

INVx4_ASAP7_75t_L g1770 ( 
.A(n_1635),
.Y(n_1770)
);

BUFx3_ASAP7_75t_L g1771 ( 
.A(n_1618),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1622),
.Y(n_1772)
);

CKINVDCx20_ASAP7_75t_R g1773 ( 
.A(n_1738),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1648),
.Y(n_1774)
);

BUFx2_ASAP7_75t_R g1775 ( 
.A(n_1725),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1747),
.Y(n_1776)
);

NAND2x1p5_ASAP7_75t_L g1777 ( 
.A(n_1680),
.B(n_626),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1720),
.A2(n_102),
.B1(n_98),
.B2(n_101),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1736),
.Y(n_1779)
);

BUFx5_ASAP7_75t_L g1780 ( 
.A(n_1751),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1626),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1654),
.Y(n_1782)
);

OAI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1699),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1732),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1661),
.Y(n_1785)
);

INVx6_ASAP7_75t_L g1786 ( 
.A(n_1733),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1683),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1663),
.Y(n_1788)
);

OAI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1724),
.A2(n_104),
.B(n_105),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1665),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1635),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_1697),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1641),
.Y(n_1793)
);

AOI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1688),
.A2(n_1706),
.B1(n_1741),
.B2(n_1643),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1668),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_SL g1796 ( 
.A1(n_1715),
.A2(n_114),
.B1(n_122),
.B2(n_106),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1647),
.Y(n_1797)
);

INVx4_ASAP7_75t_L g1798 ( 
.A(n_1662),
.Y(n_1798)
);

INVx2_ASAP7_75t_SL g1799 ( 
.A(n_1659),
.Y(n_1799)
);

INVx3_ASAP7_75t_SL g1800 ( 
.A(n_1707),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1662),
.Y(n_1801)
);

BUFx10_ASAP7_75t_L g1802 ( 
.A(n_1687),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1676),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1681),
.B(n_107),
.Y(n_1804)
);

CKINVDCx6p67_ASAP7_75t_R g1805 ( 
.A(n_1748),
.Y(n_1805)
);

CKINVDCx14_ASAP7_75t_R g1806 ( 
.A(n_1752),
.Y(n_1806)
);

OAI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1629),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_1807)
);

INVx4_ASAP7_75t_L g1808 ( 
.A(n_1748),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1656),
.Y(n_1809)
);

BUFx2_ASAP7_75t_SL g1810 ( 
.A(n_1690),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1675),
.Y(n_1811)
);

CKINVDCx11_ASAP7_75t_R g1812 ( 
.A(n_1702),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1646),
.B(n_108),
.Y(n_1813)
);

NAND2x1p5_ASAP7_75t_L g1814 ( 
.A(n_1703),
.B(n_628),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1666),
.B(n_109),
.Y(n_1815)
);

BUFx3_ASAP7_75t_L g1816 ( 
.A(n_1702),
.Y(n_1816)
);

BUFx12f_ASAP7_75t_L g1817 ( 
.A(n_1714),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1700),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1623),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1621),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_1820)
);

NAND2x1p5_ASAP7_75t_L g1821 ( 
.A(n_1651),
.B(n_629),
.Y(n_1821)
);

BUFx4f_ASAP7_75t_L g1822 ( 
.A(n_1735),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1726),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1710),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_1824)
);

INVx5_ASAP7_75t_L g1825 ( 
.A(n_1650),
.Y(n_1825)
);

BUFx3_ASAP7_75t_L g1826 ( 
.A(n_1658),
.Y(n_1826)
);

CKINVDCx20_ASAP7_75t_R g1827 ( 
.A(n_1708),
.Y(n_1827)
);

CKINVDCx20_ASAP7_75t_R g1828 ( 
.A(n_1689),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1657),
.B(n_117),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1713),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1717),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_1831)
);

INVx6_ASAP7_75t_L g1832 ( 
.A(n_1682),
.Y(n_1832)
);

BUFx4f_ASAP7_75t_SL g1833 ( 
.A(n_1704),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1713),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1718),
.A2(n_122),
.B1(n_118),
.B2(n_121),
.Y(n_1835)
);

BUFx2_ASAP7_75t_L g1836 ( 
.A(n_1705),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1669),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1630),
.A2(n_124),
.B1(n_121),
.B2(n_123),
.Y(n_1838)
);

INVx5_ASAP7_75t_L g1839 ( 
.A(n_1750),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1744),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1642),
.B(n_1627),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1617),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_SL g1843 ( 
.A1(n_1693),
.A2(n_136),
.B1(n_144),
.B2(n_128),
.Y(n_1843)
);

INVx6_ASAP7_75t_L g1844 ( 
.A(n_1685),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1616),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1637),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1679),
.B(n_1644),
.Y(n_1847)
);

CKINVDCx6p67_ASAP7_75t_R g1848 ( 
.A(n_1624),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1678),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1744),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_SL g1851 ( 
.A1(n_1664),
.A2(n_140),
.B1(n_148),
.B2(n_132),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1667),
.Y(n_1852)
);

BUFx6f_ASAP7_75t_L g1853 ( 
.A(n_1655),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1671),
.Y(n_1854)
);

CKINVDCx11_ASAP7_75t_R g1855 ( 
.A(n_1640),
.Y(n_1855)
);

INVx6_ASAP7_75t_L g1856 ( 
.A(n_1653),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1636),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1734),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_1858)
);

OAI21xp33_ASAP7_75t_L g1859 ( 
.A1(n_1723),
.A2(n_137),
.B(n_138),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1737),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_L g1861 ( 
.A(n_1719),
.Y(n_1861)
);

OAI22x1_ASAP7_75t_L g1862 ( 
.A1(n_1722),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_1862)
);

AOI21xp33_ASAP7_75t_L g1863 ( 
.A1(n_1701),
.A2(n_141),
.B(n_142),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_SL g1864 ( 
.A1(n_1740),
.A2(n_150),
.B1(n_158),
.B2(n_142),
.Y(n_1864)
);

BUFx6f_ASAP7_75t_L g1865 ( 
.A(n_1649),
.Y(n_1865)
);

BUFx2_ASAP7_75t_SL g1866 ( 
.A(n_1638),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_SL g1867 ( 
.A1(n_1645),
.A2(n_152),
.B1(n_160),
.B2(n_143),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1749),
.Y(n_1868)
);

INVx6_ASAP7_75t_L g1869 ( 
.A(n_1691),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_SL g1870 ( 
.A1(n_1694),
.A2(n_152),
.B1(n_161),
.B2(n_143),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_1684),
.Y(n_1871)
);

BUFx2_ASAP7_75t_L g1872 ( 
.A(n_1705),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1671),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1692),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1672),
.Y(n_1875)
);

INVx1_ASAP7_75t_SL g1876 ( 
.A(n_1727),
.Y(n_1876)
);

BUFx2_ASAP7_75t_SL g1877 ( 
.A(n_1728),
.Y(n_1877)
);

INVx3_ASAP7_75t_SL g1878 ( 
.A(n_1634),
.Y(n_1878)
);

AOI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1716),
.A2(n_1670),
.B1(n_1742),
.B2(n_1729),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1672),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1745),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_1881)
);

AOI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1634),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_1882)
);

BUFx2_ASAP7_75t_L g1883 ( 
.A(n_1615),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_SL g1884 ( 
.A1(n_1615),
.A2(n_159),
.B1(n_168),
.B2(n_149),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1782),
.Y(n_1885)
);

OAI21x1_ASAP7_75t_L g1886 ( 
.A1(n_1879),
.A2(n_632),
.B(n_631),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1790),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1883),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1803),
.Y(n_1889)
);

AO31x2_ASAP7_75t_L g1890 ( 
.A1(n_1875),
.A2(n_636),
.A3(n_639),
.B(n_634),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1768),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_SL g1892 ( 
.A1(n_1827),
.A2(n_154),
.B1(n_151),
.B2(n_153),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1880),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1787),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1763),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1757),
.B(n_156),
.Y(n_1896)
);

CKINVDCx20_ASAP7_75t_R g1897 ( 
.A(n_1753),
.Y(n_1897)
);

BUFx3_ASAP7_75t_L g1898 ( 
.A(n_1766),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1788),
.Y(n_1899)
);

BUFx3_ASAP7_75t_L g1900 ( 
.A(n_1791),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1795),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1769),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1772),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1774),
.Y(n_1904)
);

BUFx2_ASAP7_75t_SL g1905 ( 
.A(n_1808),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1779),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1785),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1781),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1780),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1811),
.B(n_640),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1780),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1780),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1809),
.B(n_156),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1854),
.Y(n_1914)
);

AO21x2_ASAP7_75t_L g1915 ( 
.A1(n_1789),
.A2(n_157),
.B(n_158),
.Y(n_1915)
);

OAI21x1_ASAP7_75t_L g1916 ( 
.A1(n_1868),
.A2(n_643),
.B(n_641),
.Y(n_1916)
);

OAI21x1_ASAP7_75t_L g1917 ( 
.A1(n_1840),
.A2(n_645),
.B(n_644),
.Y(n_1917)
);

CKINVDCx12_ASAP7_75t_R g1918 ( 
.A(n_1815),
.Y(n_1918)
);

BUFx3_ASAP7_75t_L g1919 ( 
.A(n_1791),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1767),
.B(n_157),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1784),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1758),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1780),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1799),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1873),
.Y(n_1925)
);

INVx3_ASAP7_75t_L g1926 ( 
.A(n_1798),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1826),
.B(n_1813),
.Y(n_1927)
);

AOI21x1_ASAP7_75t_L g1928 ( 
.A1(n_1836),
.A2(n_650),
.B(n_649),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1830),
.Y(n_1929)
);

NOR2x1p5_ASAP7_75t_L g1930 ( 
.A(n_1805),
.B(n_651),
.Y(n_1930)
);

OAI21x1_ASAP7_75t_L g1931 ( 
.A1(n_1850),
.A2(n_653),
.B(n_652),
.Y(n_1931)
);

OA21x2_ASAP7_75t_L g1932 ( 
.A1(n_1872),
.A2(n_159),
.B(n_161),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1771),
.Y(n_1933)
);

OAI21x1_ASAP7_75t_L g1934 ( 
.A1(n_1821),
.A2(n_1829),
.B(n_1881),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1834),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1862),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1852),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1832),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1878),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1839),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1841),
.B(n_656),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1839),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1869),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1793),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1847),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1844),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1802),
.Y(n_1947)
);

BUFx2_ASAP7_75t_L g1948 ( 
.A(n_1801),
.Y(n_1948)
);

BUFx3_ASAP7_75t_L g1949 ( 
.A(n_1765),
.Y(n_1949)
);

HB1xp67_ASAP7_75t_L g1950 ( 
.A(n_1856),
.Y(n_1950)
);

AND2x4_ASAP7_75t_L g1951 ( 
.A(n_1816),
.B(n_659),
.Y(n_1951)
);

INVx3_ASAP7_75t_L g1952 ( 
.A(n_1755),
.Y(n_1952)
);

BUFx3_ASAP7_75t_L g1953 ( 
.A(n_1786),
.Y(n_1953)
);

INVx2_ASAP7_75t_SL g1954 ( 
.A(n_1786),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1804),
.B(n_660),
.Y(n_1955)
);

AOI22xp33_ASAP7_75t_L g1956 ( 
.A1(n_1855),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1794),
.B(n_162),
.Y(n_1957)
);

HB1xp67_ASAP7_75t_L g1958 ( 
.A(n_1817),
.Y(n_1958)
);

BUFx6f_ASAP7_75t_L g1959 ( 
.A(n_1797),
.Y(n_1959)
);

OAI21x1_ASAP7_75t_L g1960 ( 
.A1(n_1882),
.A2(n_664),
.B(n_661),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1822),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1814),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1861),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1845),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1848),
.Y(n_1965)
);

BUFx2_ASAP7_75t_L g1966 ( 
.A(n_1792),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1871),
.Y(n_1967)
);

NAND2xp33_ASAP7_75t_R g1968 ( 
.A(n_1938),
.B(n_1819),
.Y(n_1968)
);

INVx3_ASAP7_75t_L g1969 ( 
.A(n_1953),
.Y(n_1969)
);

AO21x2_ASAP7_75t_L g1970 ( 
.A1(n_1928),
.A2(n_1863),
.B(n_1859),
.Y(n_1970)
);

AOI221xp5_ASAP7_75t_L g1971 ( 
.A1(n_1956),
.A2(n_1762),
.B1(n_1783),
.B2(n_1764),
.C(n_1807),
.Y(n_1971)
);

NOR2xp67_ASAP7_75t_L g1972 ( 
.A(n_1967),
.B(n_1950),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1927),
.B(n_1806),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1902),
.Y(n_1974)
);

AOI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1965),
.A2(n_1828),
.B1(n_1846),
.B2(n_1831),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1945),
.B(n_1884),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1898),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1903),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1921),
.B(n_1759),
.Y(n_1979)
);

AOI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1915),
.A2(n_1837),
.B(n_1849),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1904),
.B(n_1907),
.Y(n_1981)
);

NOR2xp33_ASAP7_75t_L g1982 ( 
.A(n_1964),
.B(n_1761),
.Y(n_1982)
);

OAI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1934),
.A2(n_1842),
.B(n_1838),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1906),
.Y(n_1984)
);

INVx5_ASAP7_75t_L g1985 ( 
.A(n_1959),
.Y(n_1985)
);

OAI21xp5_ASAP7_75t_L g1986 ( 
.A1(n_1957),
.A2(n_1867),
.B(n_1864),
.Y(n_1986)
);

OAI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1895),
.A2(n_1870),
.B(n_1874),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1961),
.A2(n_1876),
.B(n_1858),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1922),
.B(n_1908),
.Y(n_1989)
);

OAI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1946),
.A2(n_1823),
.B1(n_1754),
.B2(n_1756),
.Y(n_1990)
);

CKINVDCx5p33_ASAP7_75t_R g1991 ( 
.A(n_1897),
.Y(n_1991)
);

O2A1O1Ixp33_ASAP7_75t_SL g1992 ( 
.A1(n_1920),
.A2(n_1820),
.B(n_1835),
.C(n_1773),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1948),
.B(n_1777),
.Y(n_1993)
);

OAI21xp5_ASAP7_75t_L g1994 ( 
.A1(n_1960),
.A2(n_1851),
.B(n_1857),
.Y(n_1994)
);

AND2x4_ASAP7_75t_L g1995 ( 
.A(n_1933),
.B(n_1770),
.Y(n_1995)
);

OAI211xp5_ASAP7_75t_L g1996 ( 
.A1(n_1892),
.A2(n_1796),
.B(n_1778),
.C(n_1818),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1894),
.B(n_1824),
.Y(n_1997)
);

AO32x2_ASAP7_75t_L g1998 ( 
.A1(n_1929),
.A2(n_1877),
.A3(n_1843),
.B1(n_1833),
.B2(n_1860),
.Y(n_1998)
);

O2A1O1Ixp33_ASAP7_75t_SL g1999 ( 
.A1(n_1943),
.A2(n_1812),
.B(n_1760),
.C(n_1825),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1899),
.B(n_1825),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1891),
.Y(n_2001)
);

INVx5_ASAP7_75t_L g2002 ( 
.A(n_1959),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1901),
.B(n_1810),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1887),
.B(n_1866),
.Y(n_2004)
);

OA21x2_ASAP7_75t_L g2005 ( 
.A1(n_1940),
.A2(n_1865),
.B(n_1853),
.Y(n_2005)
);

AOI22xp5_ASAP7_75t_L g2006 ( 
.A1(n_1962),
.A2(n_1800),
.B1(n_1776),
.B2(n_1861),
.Y(n_2006)
);

AND2x4_ASAP7_75t_L g2007 ( 
.A(n_1961),
.B(n_1853),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1935),
.B(n_1865),
.Y(n_2008)
);

O2A1O1Ixp33_ASAP7_75t_SL g2009 ( 
.A1(n_1958),
.A2(n_1775),
.B(n_172),
.C(n_180),
.Y(n_2009)
);

HB1xp67_ASAP7_75t_L g2010 ( 
.A(n_1942),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1944),
.B(n_1936),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_1918),
.B(n_163),
.Y(n_2012)
);

INVx2_ASAP7_75t_SL g2013 ( 
.A(n_1959),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1889),
.B(n_1939),
.Y(n_2014)
);

BUFx6f_ASAP7_75t_L g2015 ( 
.A(n_1900),
.Y(n_2015)
);

BUFx12f_ASAP7_75t_L g2016 ( 
.A(n_1949),
.Y(n_2016)
);

OAI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_1896),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_2017)
);

OAI21xp5_ASAP7_75t_L g2018 ( 
.A1(n_1955),
.A2(n_666),
.B(n_665),
.Y(n_2018)
);

AOI22xp33_ASAP7_75t_L g2019 ( 
.A1(n_1941),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_2019)
);

OR2x2_ASAP7_75t_L g2020 ( 
.A(n_1888),
.B(n_168),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1939),
.B(n_169),
.Y(n_2021)
);

AOI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1930),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_2022)
);

INVxp67_ASAP7_75t_L g2023 ( 
.A(n_1924),
.Y(n_2023)
);

BUFx3_ASAP7_75t_L g2024 ( 
.A(n_1919),
.Y(n_2024)
);

OAI211xp5_ASAP7_75t_SL g2025 ( 
.A1(n_1913),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_2025)
);

A2O1A1Ixp33_ASAP7_75t_L g2026 ( 
.A1(n_1886),
.A2(n_175),
.B(n_173),
.C(n_174),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1885),
.B(n_175),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1888),
.B(n_176),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1910),
.B(n_177),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1926),
.B(n_177),
.Y(n_2030)
);

OA21x2_ASAP7_75t_L g2031 ( 
.A1(n_1893),
.A2(n_178),
.B(n_179),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1926),
.B(n_178),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_1963),
.B(n_667),
.Y(n_2033)
);

AND2x6_ASAP7_75t_L g2034 ( 
.A(n_1951),
.B(n_1909),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1893),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1911),
.B(n_179),
.Y(n_2036)
);

AOI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_1951),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1912),
.B(n_182),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1914),
.Y(n_2039)
);

NOR2x1_ASAP7_75t_SL g2040 ( 
.A(n_1928),
.B(n_668),
.Y(n_2040)
);

OAI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_1947),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_2041)
);

INVxp67_ASAP7_75t_L g2042 ( 
.A(n_1954),
.Y(n_2042)
);

NOR2xp33_ASAP7_75t_L g2043 ( 
.A(n_1977),
.B(n_1947),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_2014),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1974),
.Y(n_2045)
);

OR2x2_ASAP7_75t_L g2046 ( 
.A(n_1989),
.B(n_1914),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2035),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2039),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_L g2049 ( 
.A(n_1969),
.B(n_1966),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1978),
.Y(n_2050)
);

OAI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_1975),
.A2(n_1905),
.B1(n_1932),
.B2(n_1937),
.Y(n_2051)
);

INVx2_ASAP7_75t_SL g2052 ( 
.A(n_1985),
.Y(n_2052)
);

OR2x2_ASAP7_75t_L g2053 ( 
.A(n_1984),
.B(n_1925),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1973),
.B(n_2011),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_2001),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1981),
.Y(n_2056)
);

INVx2_ASAP7_75t_SL g2057 ( 
.A(n_1985),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_1971),
.A2(n_1905),
.B1(n_1932),
.B2(n_1952),
.Y(n_2058)
);

HB1xp67_ASAP7_75t_L g2059 ( 
.A(n_2010),
.Y(n_2059)
);

INVx2_ASAP7_75t_SL g2060 ( 
.A(n_2002),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1972),
.B(n_1923),
.Y(n_2061)
);

INVx2_ASAP7_75t_SL g2062 ( 
.A(n_2002),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_2003),
.B(n_1890),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1979),
.B(n_1952),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2008),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2004),
.Y(n_2066)
);

AND2x4_ASAP7_75t_L g2067 ( 
.A(n_2007),
.B(n_1890),
.Y(n_2067)
);

NOR2x1_ASAP7_75t_L g2068 ( 
.A(n_2000),
.B(n_2031),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1993),
.B(n_1890),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_2013),
.B(n_1917),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2023),
.B(n_1931),
.Y(n_2071)
);

INVx4_ASAP7_75t_L g2072 ( 
.A(n_1995),
.Y(n_2072)
);

BUFx3_ASAP7_75t_L g2073 ( 
.A(n_2016),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2020),
.Y(n_2074)
);

INVx1_ASAP7_75t_SL g2075 ( 
.A(n_2024),
.Y(n_2075)
);

OR2x2_ASAP7_75t_L g2076 ( 
.A(n_2028),
.B(n_1916),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1976),
.B(n_183),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2021),
.B(n_185),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2027),
.B(n_186),
.Y(n_2079)
);

BUFx3_ASAP7_75t_L g2080 ( 
.A(n_2015),
.Y(n_2080)
);

NOR2x1_ASAP7_75t_SL g2081 ( 
.A(n_1970),
.B(n_187),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_2036),
.B(n_186),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2038),
.B(n_188),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1980),
.B(n_188),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2005),
.Y(n_2085)
);

HB1xp67_ASAP7_75t_L g2086 ( 
.A(n_1997),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_1982),
.B(n_2042),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_R g2088 ( 
.A(n_1991),
.B(n_189),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1988),
.B(n_189),
.Y(n_2089)
);

HB1xp67_ASAP7_75t_L g2090 ( 
.A(n_2030),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2032),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_2015),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2034),
.B(n_190),
.Y(n_2093)
);

OAI22xp5_ASAP7_75t_L g2094 ( 
.A1(n_2022),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2040),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2012),
.B(n_191),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2006),
.B(n_2029),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_2034),
.Y(n_2098)
);

BUFx3_ASAP7_75t_L g2099 ( 
.A(n_2034),
.Y(n_2099)
);

AOI22xp33_ASAP7_75t_L g2100 ( 
.A1(n_1986),
.A2(n_1987),
.B1(n_1983),
.B2(n_1994),
.Y(n_2100)
);

NOR2xp67_ASAP7_75t_L g2101 ( 
.A(n_2017),
.B(n_192),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2033),
.B(n_193),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1998),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_2025),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1998),
.B(n_194),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2018),
.B(n_196),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2026),
.B(n_196),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2037),
.B(n_197),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_L g2109 ( 
.A(n_1968),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2019),
.B(n_197),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_2041),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_1990),
.B(n_198),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_1999),
.B(n_198),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_2009),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1992),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_1996),
.B(n_199),
.Y(n_2116)
);

HB1xp67_ASAP7_75t_L g2117 ( 
.A(n_2010),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1973),
.B(n_199),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_2014),
.Y(n_2119)
);

AND2x2_ASAP7_75t_SL g2120 ( 
.A(n_1976),
.B(n_200),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_1973),
.B(n_200),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2035),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2035),
.Y(n_2123)
);

BUFx2_ASAP7_75t_L g2124 ( 
.A(n_2085),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2086),
.B(n_201),
.Y(n_2125)
);

OAI31xp33_ASAP7_75t_L g2126 ( 
.A1(n_2100),
.A2(n_203),
.A3(n_201),
.B(n_202),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2045),
.Y(n_2127)
);

HB1xp67_ASAP7_75t_L g2128 ( 
.A(n_2059),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2050),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2117),
.Y(n_2130)
);

AO21x2_ASAP7_75t_L g2131 ( 
.A1(n_2084),
.A2(n_202),
.B(n_203),
.Y(n_2131)
);

AO22x1_ASAP7_75t_L g2132 ( 
.A1(n_2109),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_2132)
);

INVx2_ASAP7_75t_SL g2133 ( 
.A(n_2080),
.Y(n_2133)
);

AO221x2_ASAP7_75t_L g2134 ( 
.A1(n_2051),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.C(n_207),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2047),
.Y(n_2135)
);

AOI22xp33_ASAP7_75t_L g2136 ( 
.A1(n_2120),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2065),
.B(n_208),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2048),
.Y(n_2138)
);

AOI21x1_ASAP7_75t_L g2139 ( 
.A1(n_2089),
.A2(n_210),
.B(n_211),
.Y(n_2139)
);

OR2x2_ASAP7_75t_L g2140 ( 
.A(n_2046),
.B(n_212),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2055),
.Y(n_2141)
);

INVx1_ASAP7_75t_SL g2142 ( 
.A(n_2075),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2122),
.Y(n_2143)
);

INVx3_ASAP7_75t_L g2144 ( 
.A(n_2072),
.Y(n_2144)
);

BUFx2_ASAP7_75t_L g2145 ( 
.A(n_2099),
.Y(n_2145)
);

NOR3xp33_ASAP7_75t_SL g2146 ( 
.A(n_2094),
.B(n_213),
.C(n_214),
.Y(n_2146)
);

INVxp67_ASAP7_75t_L g2147 ( 
.A(n_2090),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_2123),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2044),
.B(n_213),
.Y(n_2149)
);

AOI221x1_ASAP7_75t_L g2150 ( 
.A1(n_2114),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.C(n_217),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2119),
.B(n_215),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2061),
.Y(n_2152)
);

AND2x4_ASAP7_75t_SL g2153 ( 
.A(n_2109),
.B(n_669),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2053),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2056),
.Y(n_2155)
);

BUFx2_ASAP7_75t_L g2156 ( 
.A(n_2072),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2066),
.Y(n_2157)
);

OAI221xp5_ASAP7_75t_L g2158 ( 
.A1(n_2104),
.A2(n_2058),
.B1(n_2112),
.B2(n_2101),
.C(n_2115),
.Y(n_2158)
);

HB1xp67_ASAP7_75t_L g2159 ( 
.A(n_2068),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2074),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2054),
.B(n_2069),
.Y(n_2161)
);

AOI22xp33_ASAP7_75t_L g2162 ( 
.A1(n_2116),
.A2(n_219),
.B1(n_216),
.B2(n_218),
.Y(n_2162)
);

INVxp67_ASAP7_75t_L g2163 ( 
.A(n_2091),
.Y(n_2163)
);

OR2x2_ASAP7_75t_L g2164 ( 
.A(n_2063),
.B(n_218),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2064),
.B(n_221),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2098),
.B(n_221),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2097),
.B(n_222),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2071),
.Y(n_2168)
);

OA21x2_ASAP7_75t_L g2169 ( 
.A1(n_2103),
.A2(n_223),
.B(n_224),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2092),
.B(n_223),
.Y(n_2170)
);

BUFx3_ASAP7_75t_L g2171 ( 
.A(n_2073),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2076),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_2067),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2067),
.Y(n_2174)
);

AOI22xp5_ASAP7_75t_L g2175 ( 
.A1(n_2113),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2087),
.B(n_225),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2095),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2105),
.B(n_226),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2070),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2070),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2043),
.B(n_227),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2049),
.B(n_227),
.Y(n_2182)
);

OAI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_2109),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_2077),
.B(n_228),
.Y(n_2184)
);

AOI22xp33_ASAP7_75t_SL g2185 ( 
.A1(n_2106),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2081),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2093),
.B(n_231),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2052),
.B(n_232),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2057),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2060),
.Y(n_2190)
);

AOI221xp5_ASAP7_75t_L g2191 ( 
.A1(n_2107),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.C(n_235),
.Y(n_2191)
);

AO21x2_ASAP7_75t_L g2192 ( 
.A1(n_2088),
.A2(n_234),
.B(n_235),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2062),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_2118),
.B(n_236),
.Y(n_2194)
);

NAND3xp33_ASAP7_75t_L g2195 ( 
.A(n_2111),
.B(n_236),
.C(n_237),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_2121),
.Y(n_2196)
);

OR2x2_ASAP7_75t_L g2197 ( 
.A(n_2079),
.B(n_238),
.Y(n_2197)
);

BUFx2_ASAP7_75t_L g2198 ( 
.A(n_2113),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2078),
.B(n_238),
.Y(n_2199)
);

INVx5_ASAP7_75t_L g2200 ( 
.A(n_2102),
.Y(n_2200)
);

INVxp67_ASAP7_75t_L g2201 ( 
.A(n_2082),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2096),
.B(n_239),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2083),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2110),
.Y(n_2204)
);

NAND3xp33_ASAP7_75t_SL g2205 ( 
.A(n_2108),
.B(n_239),
.C(n_240),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_2059),
.B(n_241),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2059),
.B(n_241),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2045),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_2059),
.B(n_242),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2047),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2045),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2086),
.B(n_243),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2047),
.Y(n_2213)
);

OAI33xp33_ASAP7_75t_L g2214 ( 
.A1(n_2084),
.A2(n_245),
.A3(n_247),
.B1(n_243),
.B2(n_244),
.B3(n_246),
.Y(n_2214)
);

AO31x2_ASAP7_75t_L g2215 ( 
.A1(n_2085),
.A2(n_248),
.A3(n_244),
.B(n_246),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2047),
.Y(n_2216)
);

AND2x4_ASAP7_75t_L g2217 ( 
.A(n_2098),
.B(n_248),
.Y(n_2217)
);

INVx2_ASAP7_75t_SL g2218 ( 
.A(n_2080),
.Y(n_2218)
);

OAI31xp33_ASAP7_75t_SL g2219 ( 
.A1(n_2051),
.A2(n_251),
.A3(n_249),
.B(n_250),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2059),
.B(n_249),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2045),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2047),
.Y(n_2222)
);

OR2x2_ASAP7_75t_L g2223 ( 
.A(n_2172),
.B(n_250),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2135),
.Y(n_2224)
);

INVx1_ASAP7_75t_SL g2225 ( 
.A(n_2142),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2156),
.B(n_2161),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2177),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2138),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2128),
.B(n_251),
.Y(n_2229)
);

OR2x2_ASAP7_75t_L g2230 ( 
.A(n_2147),
.B(n_252),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2143),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2130),
.B(n_253),
.Y(n_2232)
);

INVxp67_ASAP7_75t_L g2233 ( 
.A(n_2192),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2168),
.B(n_253),
.Y(n_2234)
);

BUFx2_ASAP7_75t_L g2235 ( 
.A(n_2198),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2210),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2213),
.Y(n_2237)
);

OR2x2_ASAP7_75t_L g2238 ( 
.A(n_2154),
.B(n_254),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2144),
.B(n_254),
.Y(n_2239)
);

NAND4xp25_ASAP7_75t_L g2240 ( 
.A(n_2219),
.B(n_257),
.C(n_255),
.D(n_256),
.Y(n_2240)
);

BUFx2_ASAP7_75t_L g2241 ( 
.A(n_2124),
.Y(n_2241)
);

OR2x2_ASAP7_75t_L g2242 ( 
.A(n_2164),
.B(n_255),
.Y(n_2242)
);

INVxp67_ASAP7_75t_L g2243 ( 
.A(n_2186),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2124),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2216),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_2179),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2157),
.B(n_256),
.Y(n_2247)
);

INVx2_ASAP7_75t_SL g2248 ( 
.A(n_2200),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2222),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2173),
.B(n_257),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_2180),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2148),
.Y(n_2252)
);

OR2x2_ASAP7_75t_L g2253 ( 
.A(n_2152),
.B(n_258),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2129),
.Y(n_2254)
);

OR2x2_ASAP7_75t_L g2255 ( 
.A(n_2163),
.B(n_258),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2160),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2203),
.B(n_259),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2145),
.B(n_260),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2174),
.B(n_261),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2127),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2190),
.B(n_262),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2193),
.B(n_262),
.Y(n_2262)
);

INVx4_ASAP7_75t_L g2263 ( 
.A(n_2171),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2208),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_2200),
.B(n_263),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2189),
.B(n_2159),
.Y(n_2266)
);

AND2x4_ASAP7_75t_L g2267 ( 
.A(n_2133),
.B(n_263),
.Y(n_2267)
);

OR2x2_ASAP7_75t_L g2268 ( 
.A(n_2141),
.B(n_264),
.Y(n_2268)
);

INVx3_ASAP7_75t_L g2269 ( 
.A(n_2218),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2155),
.B(n_2211),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2196),
.B(n_264),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2200),
.B(n_265),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2221),
.Y(n_2273)
);

NOR2xp33_ASAP7_75t_L g2274 ( 
.A(n_2201),
.B(n_265),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2169),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2204),
.B(n_266),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2140),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2206),
.B(n_266),
.Y(n_2278)
);

NAND2xp33_ASAP7_75t_R g2279 ( 
.A(n_2146),
.B(n_267),
.Y(n_2279)
);

OR2x2_ASAP7_75t_L g2280 ( 
.A(n_2125),
.B(n_268),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_2207),
.B(n_269),
.Y(n_2281)
);

AND2x6_ASAP7_75t_SL g2282 ( 
.A(n_2178),
.B(n_270),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2209),
.B(n_270),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2169),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2212),
.B(n_271),
.Y(n_2285)
);

INVxp67_ASAP7_75t_L g2286 ( 
.A(n_2131),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2149),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2220),
.B(n_271),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2165),
.B(n_272),
.Y(n_2289)
);

OR2x2_ASAP7_75t_L g2290 ( 
.A(n_2187),
.B(n_272),
.Y(n_2290)
);

OR2x2_ASAP7_75t_L g2291 ( 
.A(n_2184),
.B(n_273),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2151),
.Y(n_2292)
);

OR2x2_ASAP7_75t_L g2293 ( 
.A(n_2197),
.B(n_273),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2137),
.B(n_274),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2215),
.Y(n_2295)
);

OR2x2_ASAP7_75t_L g2296 ( 
.A(n_2167),
.B(n_274),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2176),
.B(n_275),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2215),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2166),
.Y(n_2299)
);

INVx3_ASAP7_75t_L g2300 ( 
.A(n_2170),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2181),
.B(n_2182),
.Y(n_2301)
);

HB1xp67_ASAP7_75t_L g2302 ( 
.A(n_2139),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2188),
.B(n_275),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2134),
.B(n_276),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2202),
.B(n_276),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2217),
.Y(n_2306)
);

AND2x4_ASAP7_75t_L g2307 ( 
.A(n_2153),
.B(n_277),
.Y(n_2307)
);

BUFx2_ASAP7_75t_L g2308 ( 
.A(n_2132),
.Y(n_2308)
);

OR2x2_ASAP7_75t_L g2309 ( 
.A(n_2199),
.B(n_277),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2194),
.B(n_278),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2134),
.B(n_279),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2158),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2195),
.Y(n_2313)
);

NAND2x1_ASAP7_75t_L g2314 ( 
.A(n_2175),
.B(n_279),
.Y(n_2314)
);

OR2x2_ASAP7_75t_L g2315 ( 
.A(n_2205),
.B(n_280),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2150),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2185),
.B(n_280),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2191),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2162),
.B(n_281),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2136),
.B(n_281),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_2126),
.B(n_282),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_2214),
.B(n_282),
.Y(n_2322)
);

OR2x6_ASAP7_75t_SL g2323 ( 
.A(n_2183),
.B(n_283),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_L g2324 ( 
.A(n_2171),
.B(n_284),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2135),
.Y(n_2325)
);

OR2x2_ASAP7_75t_L g2326 ( 
.A(n_2172),
.B(n_284),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2156),
.B(n_285),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2135),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2135),
.Y(n_2329)
);

OR2x2_ASAP7_75t_L g2330 ( 
.A(n_2172),
.B(n_285),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2156),
.B(n_286),
.Y(n_2331)
);

AND2x4_ASAP7_75t_SL g2332 ( 
.A(n_2144),
.B(n_286),
.Y(n_2332)
);

OR2x2_ASAP7_75t_L g2333 ( 
.A(n_2172),
.B(n_287),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2177),
.Y(n_2334)
);

OR2x6_ASAP7_75t_L g2335 ( 
.A(n_2248),
.B(n_287),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2224),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2235),
.B(n_288),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2228),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2235),
.B(n_288),
.Y(n_2339)
);

OR2x2_ASAP7_75t_L g2340 ( 
.A(n_2277),
.B(n_289),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2241),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2241),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2231),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2236),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2237),
.Y(n_2345)
);

AND2x4_ASAP7_75t_L g2346 ( 
.A(n_2269),
.B(n_289),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2233),
.B(n_290),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2245),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2302),
.B(n_290),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2249),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2226),
.B(n_291),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2325),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2328),
.Y(n_2353)
);

AND2x4_ASAP7_75t_SL g2354 ( 
.A(n_2263),
.B(n_291),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2266),
.B(n_292),
.Y(n_2355)
);

OAI21xp33_ASAP7_75t_SL g2356 ( 
.A1(n_2275),
.A2(n_292),
.B(n_293),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2329),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2256),
.Y(n_2358)
);

NOR2x1p5_ASAP7_75t_L g2359 ( 
.A(n_2314),
.B(n_293),
.Y(n_2359)
);

INVxp67_ASAP7_75t_L g2360 ( 
.A(n_2308),
.Y(n_2360)
);

OR2x2_ASAP7_75t_L g2361 ( 
.A(n_2286),
.B(n_294),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2295),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2227),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2300),
.B(n_2299),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2313),
.B(n_294),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2298),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2252),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2243),
.B(n_295),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2254),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2334),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2225),
.B(n_296),
.Y(n_2371)
);

INVxp67_ASAP7_75t_L g2372 ( 
.A(n_2308),
.Y(n_2372)
);

HB1xp67_ASAP7_75t_L g2373 ( 
.A(n_2284),
.Y(n_2373)
);

INVxp33_ASAP7_75t_SL g2374 ( 
.A(n_2311),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2301),
.B(n_2287),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2270),
.Y(n_2376)
);

OR2x2_ASAP7_75t_L g2377 ( 
.A(n_2260),
.B(n_296),
.Y(n_2377)
);

INVxp67_ASAP7_75t_L g2378 ( 
.A(n_2272),
.Y(n_2378)
);

AND2x2_ASAP7_75t_L g2379 ( 
.A(n_2292),
.B(n_297),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2264),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2312),
.B(n_297),
.Y(n_2381)
);

INVxp67_ASAP7_75t_L g2382 ( 
.A(n_2265),
.Y(n_2382)
);

NAND3xp33_ASAP7_75t_L g2383 ( 
.A(n_2318),
.B(n_2279),
.C(n_2316),
.Y(n_2383)
);

AND2x2_ASAP7_75t_L g2384 ( 
.A(n_2246),
.B(n_298),
.Y(n_2384)
);

AND2x2_ASAP7_75t_L g2385 ( 
.A(n_2251),
.B(n_298),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2244),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2273),
.Y(n_2387)
);

INVxp67_ASAP7_75t_SL g2388 ( 
.A(n_2234),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2268),
.Y(n_2389)
);

HB1xp67_ASAP7_75t_L g2390 ( 
.A(n_2223),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2306),
.Y(n_2391)
);

OR2x2_ASAP7_75t_L g2392 ( 
.A(n_2326),
.B(n_299),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2247),
.B(n_299),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2255),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2253),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2257),
.B(n_300),
.Y(n_2396)
);

HB1xp67_ASAP7_75t_L g2397 ( 
.A(n_2330),
.Y(n_2397)
);

INVx1_ASAP7_75t_SL g2398 ( 
.A(n_2327),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2238),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2333),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2230),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2242),
.Y(n_2402)
);

OR2x2_ASAP7_75t_L g2403 ( 
.A(n_2232),
.B(n_301),
.Y(n_2403)
);

OR2x2_ASAP7_75t_L g2404 ( 
.A(n_2229),
.B(n_301),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_2259),
.B(n_302),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2250),
.B(n_302),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2271),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2276),
.Y(n_2408)
);

INVx2_ASAP7_75t_SL g2409 ( 
.A(n_2267),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2261),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2331),
.B(n_2262),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2239),
.Y(n_2412)
);

AND2x4_ASAP7_75t_L g2413 ( 
.A(n_2258),
.B(n_2332),
.Y(n_2413)
);

AND2x4_ASAP7_75t_L g2414 ( 
.A(n_2280),
.B(n_303),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2278),
.B(n_303),
.Y(n_2415)
);

OR2x2_ASAP7_75t_L g2416 ( 
.A(n_2290),
.B(n_2296),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2291),
.Y(n_2417)
);

AOI22xp5_ASAP7_75t_L g2418 ( 
.A1(n_2240),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2293),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2274),
.B(n_304),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2281),
.B(n_306),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2283),
.B(n_307),
.Y(n_2422)
);

AOI322xp5_ASAP7_75t_L g2423 ( 
.A1(n_2304),
.A2(n_312),
.A3(n_311),
.B1(n_309),
.B2(n_307),
.C1(n_308),
.C2(n_310),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2285),
.B(n_308),
.Y(n_2424)
);

OR2x2_ASAP7_75t_L g2425 ( 
.A(n_2309),
.B(n_309),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2303),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2315),
.Y(n_2427)
);

AND2x4_ASAP7_75t_L g2428 ( 
.A(n_2288),
.B(n_310),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2322),
.B(n_2294),
.Y(n_2429)
);

NOR2x1_ASAP7_75t_L g2430 ( 
.A(n_2324),
.B(n_312),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2297),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2289),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2305),
.Y(n_2433)
);

AND2x2_ASAP7_75t_L g2434 ( 
.A(n_2310),
.B(n_313),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2282),
.B(n_313),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2323),
.B(n_2307),
.Y(n_2436)
);

OAI22xp5_ASAP7_75t_L g2437 ( 
.A1(n_2317),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_2321),
.B(n_314),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2320),
.B(n_315),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2319),
.B(n_316),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2224),
.Y(n_2441)
);

INVx1_ASAP7_75t_SL g2442 ( 
.A(n_2225),
.Y(n_2442)
);

AND2x2_ASAP7_75t_L g2443 ( 
.A(n_2235),
.B(n_317),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2224),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2235),
.B(n_317),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2224),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2224),
.Y(n_2447)
);

OR2x2_ASAP7_75t_L g2448 ( 
.A(n_2235),
.B(n_318),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2224),
.Y(n_2449)
);

NAND3xp33_ASAP7_75t_L g2450 ( 
.A(n_2302),
.B(n_320),
.C(n_321),
.Y(n_2450)
);

AND2x2_ASAP7_75t_L g2451 ( 
.A(n_2235),
.B(n_321),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2235),
.B(n_322),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2224),
.Y(n_2453)
);

OR2x2_ASAP7_75t_L g2454 ( 
.A(n_2235),
.B(n_322),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2224),
.Y(n_2455)
);

AND2x2_ASAP7_75t_L g2456 ( 
.A(n_2235),
.B(n_323),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2235),
.B(n_323),
.Y(n_2457)
);

OAI21xp5_ASAP7_75t_L g2458 ( 
.A1(n_2233),
.A2(n_324),
.B(n_325),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2233),
.B(n_326),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2233),
.B(n_326),
.Y(n_2460)
);

OR2x2_ASAP7_75t_L g2461 ( 
.A(n_2235),
.B(n_327),
.Y(n_2461)
);

OR2x2_ASAP7_75t_L g2462 ( 
.A(n_2235),
.B(n_327),
.Y(n_2462)
);

OR2x2_ASAP7_75t_L g2463 ( 
.A(n_2235),
.B(n_328),
.Y(n_2463)
);

HB1xp67_ASAP7_75t_SL g2464 ( 
.A(n_2308),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2224),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2235),
.B(n_329),
.Y(n_2466)
);

NOR2xp33_ASAP7_75t_L g2467 ( 
.A(n_2263),
.B(n_330),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2233),
.B(n_330),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2233),
.B(n_331),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2235),
.B(n_332),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2235),
.B(n_332),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2224),
.Y(n_2472)
);

NOR2x1_ASAP7_75t_L g2473 ( 
.A(n_2308),
.B(n_333),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2224),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2224),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2224),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2224),
.Y(n_2477)
);

NOR2xp33_ASAP7_75t_L g2478 ( 
.A(n_2263),
.B(n_333),
.Y(n_2478)
);

AND2x4_ASAP7_75t_L g2479 ( 
.A(n_2235),
.B(n_334),
.Y(n_2479)
);

OR2x2_ASAP7_75t_L g2480 ( 
.A(n_2235),
.B(n_334),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2235),
.B(n_335),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2235),
.B(n_335),
.Y(n_2482)
);

OR2x2_ASAP7_75t_L g2483 ( 
.A(n_2235),
.B(n_336),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2233),
.B(n_336),
.Y(n_2484)
);

INVx3_ASAP7_75t_L g2485 ( 
.A(n_2263),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2235),
.B(n_337),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2224),
.Y(n_2487)
);

OR2x2_ASAP7_75t_L g2488 ( 
.A(n_2235),
.B(n_338),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2224),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2235),
.B(n_338),
.Y(n_2490)
);

A2O1A1Ixp33_ASAP7_75t_L g2491 ( 
.A1(n_2308),
.A2(n_342),
.B(n_339),
.C(n_340),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2224),
.Y(n_2492)
);

HB1xp67_ASAP7_75t_L g2493 ( 
.A(n_2235),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2235),
.Y(n_2494)
);

AOI211xp5_ASAP7_75t_L g2495 ( 
.A1(n_2308),
.A2(n_342),
.B(n_339),
.C(n_340),
.Y(n_2495)
);

INVxp67_ASAP7_75t_SL g2496 ( 
.A(n_2233),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2233),
.B(n_343),
.Y(n_2497)
);

NOR2x1_ASAP7_75t_L g2498 ( 
.A(n_2308),
.B(n_343),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2224),
.Y(n_2499)
);

INVx2_ASAP7_75t_SL g2500 ( 
.A(n_2248),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2224),
.Y(n_2501)
);

OR2x2_ASAP7_75t_L g2502 ( 
.A(n_2360),
.B(n_2372),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_R g2503 ( 
.A(n_2500),
.B(n_344),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2378),
.B(n_344),
.Y(n_2504)
);

AND2x2_ASAP7_75t_L g2505 ( 
.A(n_2364),
.B(n_345),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2388),
.B(n_345),
.Y(n_2506)
);

INVx1_ASAP7_75t_SL g2507 ( 
.A(n_2464),
.Y(n_2507)
);

AOI21xp33_ASAP7_75t_SL g2508 ( 
.A1(n_2383),
.A2(n_346),
.B(n_347),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2362),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_2427),
.B(n_346),
.Y(n_2510)
);

OR2x2_ASAP7_75t_L g2511 ( 
.A(n_2416),
.B(n_347),
.Y(n_2511)
);

BUFx2_ASAP7_75t_L g2512 ( 
.A(n_2493),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2382),
.B(n_348),
.Y(n_2513)
);

INVxp67_ASAP7_75t_SL g2514 ( 
.A(n_2473),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2366),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2417),
.B(n_349),
.Y(n_2516)
);

INVx1_ASAP7_75t_SL g2517 ( 
.A(n_2442),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2419),
.B(n_349),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_SL g2519 ( 
.A(n_2485),
.B(n_350),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2402),
.B(n_350),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2494),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2375),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_SL g2523 ( 
.A(n_2374),
.B(n_351),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2389),
.B(n_351),
.Y(n_2524)
);

AND2x2_ASAP7_75t_SL g2525 ( 
.A(n_2436),
.B(n_352),
.Y(n_2525)
);

AO221x1_ASAP7_75t_L g2526 ( 
.A1(n_2341),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.C(n_355),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2391),
.B(n_356),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2373),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2390),
.B(n_356),
.Y(n_2529)
);

INVx2_ASAP7_75t_SL g2530 ( 
.A(n_2479),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2336),
.Y(n_2531)
);

INVx1_ASAP7_75t_SL g2532 ( 
.A(n_2354),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2338),
.Y(n_2533)
);

NAND2xp33_ASAP7_75t_SL g2534 ( 
.A(n_2359),
.B(n_357),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2397),
.B(n_358),
.Y(n_2535)
);

OAI31xp33_ASAP7_75t_L g2536 ( 
.A1(n_2491),
.A2(n_360),
.A3(n_358),
.B(n_359),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2343),
.Y(n_2537)
);

OR2x2_ASAP7_75t_L g2538 ( 
.A(n_2394),
.B(n_359),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2401),
.B(n_360),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2395),
.B(n_361),
.Y(n_2540)
);

INVx1_ASAP7_75t_SL g2541 ( 
.A(n_2413),
.Y(n_2541)
);

HB1xp67_ASAP7_75t_L g2542 ( 
.A(n_2342),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2399),
.B(n_361),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2344),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2400),
.B(n_362),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2349),
.B(n_362),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2345),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2412),
.Y(n_2548)
);

AOI211xp5_ASAP7_75t_SL g2549 ( 
.A1(n_2495),
.A2(n_365),
.B(n_363),
.C(n_364),
.Y(n_2549)
);

INVxp33_ASAP7_75t_L g2550 ( 
.A(n_2498),
.Y(n_2550)
);

AND2x4_ASAP7_75t_L g2551 ( 
.A(n_2496),
.B(n_2348),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2350),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2398),
.B(n_363),
.Y(n_2553)
);

AOI21xp5_ASAP7_75t_L g2554 ( 
.A1(n_2435),
.A2(n_364),
.B(n_365),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2426),
.B(n_366),
.Y(n_2555)
);

AOI22xp33_ASAP7_75t_L g2556 ( 
.A1(n_2458),
.A2(n_370),
.B1(n_367),
.B2(n_369),
.Y(n_2556)
);

OR2x2_ASAP7_75t_L g2557 ( 
.A(n_2386),
.B(n_367),
.Y(n_2557)
);

NOR3xp33_ASAP7_75t_L g2558 ( 
.A(n_2450),
.B(n_371),
.C(n_372),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2337),
.B(n_373),
.Y(n_2559)
);

AND2x2_ASAP7_75t_L g2560 ( 
.A(n_2432),
.B(n_373),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2363),
.Y(n_2561)
);

NOR3xp33_ASAP7_75t_L g2562 ( 
.A(n_2437),
.B(n_374),
.C(n_375),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2411),
.B(n_376),
.Y(n_2563)
);

OR2x2_ASAP7_75t_L g2564 ( 
.A(n_2376),
.B(n_376),
.Y(n_2564)
);

INVx1_ASAP7_75t_SL g2565 ( 
.A(n_2339),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2410),
.B(n_377),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2370),
.Y(n_2567)
);

AND2x2_ASAP7_75t_L g2568 ( 
.A(n_2431),
.B(n_377),
.Y(n_2568)
);

INVx1_ASAP7_75t_SL g2569 ( 
.A(n_2443),
.Y(n_2569)
);

NOR2xp33_ASAP7_75t_SL g2570 ( 
.A(n_2430),
.B(n_2467),
.Y(n_2570)
);

OR2x2_ASAP7_75t_L g2571 ( 
.A(n_2408),
.B(n_378),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2445),
.B(n_2451),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2352),
.Y(n_2573)
);

OR2x2_ASAP7_75t_L g2574 ( 
.A(n_2433),
.B(n_378),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2407),
.B(n_379),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2377),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2452),
.B(n_379),
.Y(n_2577)
);

OR2x2_ASAP7_75t_L g2578 ( 
.A(n_2380),
.B(n_380),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2351),
.B(n_380),
.Y(n_2579)
);

OR2x2_ASAP7_75t_L g2580 ( 
.A(n_2387),
.B(n_381),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2456),
.B(n_381),
.Y(n_2581)
);

AND2x4_ASAP7_75t_L g2582 ( 
.A(n_2353),
.B(n_2357),
.Y(n_2582)
);

BUFx2_ASAP7_75t_L g2583 ( 
.A(n_2335),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2358),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2457),
.B(n_382),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2441),
.Y(n_2586)
);

OR2x2_ASAP7_75t_L g2587 ( 
.A(n_2367),
.B(n_382),
.Y(n_2587)
);

NAND2x1_ASAP7_75t_L g2588 ( 
.A(n_2444),
.B(n_383),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2446),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2447),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2449),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2466),
.B(n_2470),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2453),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2355),
.B(n_383),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2455),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2465),
.Y(n_2596)
);

NOR2xp33_ASAP7_75t_L g2597 ( 
.A(n_2429),
.B(n_384),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2409),
.B(n_384),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2471),
.B(n_385),
.Y(n_2599)
);

NAND3xp33_ASAP7_75t_L g2600 ( 
.A(n_2423),
.B(n_385),
.C(n_386),
.Y(n_2600)
);

HB1xp67_ASAP7_75t_L g2601 ( 
.A(n_2448),
.Y(n_2601)
);

INVxp67_ASAP7_75t_L g2602 ( 
.A(n_2361),
.Y(n_2602)
);

NOR2xp33_ASAP7_75t_L g2603 ( 
.A(n_2365),
.B(n_387),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2472),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2481),
.B(n_387),
.Y(n_2605)
);

NAND3xp33_ASAP7_75t_SL g2606 ( 
.A(n_2418),
.B(n_388),
.C(n_389),
.Y(n_2606)
);

AO21x1_ASAP7_75t_L g2607 ( 
.A1(n_2347),
.A2(n_389),
.B(n_390),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2482),
.B(n_390),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2474),
.Y(n_2609)
);

NOR2xp33_ASAP7_75t_L g2610 ( 
.A(n_2381),
.B(n_391),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2475),
.Y(n_2611)
);

NAND2x1_ASAP7_75t_L g2612 ( 
.A(n_2476),
.B(n_391),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2477),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2487),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2489),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2486),
.B(n_392),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2490),
.B(n_392),
.Y(n_2617)
);

NOR4xp25_ASAP7_75t_L g2618 ( 
.A(n_2356),
.B(n_395),
.C(n_393),
.D(n_394),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2368),
.B(n_393),
.Y(n_2619)
);

AND2x2_ASAP7_75t_L g2620 ( 
.A(n_2379),
.B(n_394),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2371),
.B(n_395),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2492),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2499),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2501),
.Y(n_2624)
);

AOI31xp33_ASAP7_75t_L g2625 ( 
.A1(n_2454),
.A2(n_398),
.A3(n_396),
.B(n_397),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2514),
.B(n_2459),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2512),
.Y(n_2627)
);

AOI22xp5_ASAP7_75t_L g2628 ( 
.A1(n_2600),
.A2(n_2478),
.B1(n_2468),
.B2(n_2469),
.Y(n_2628)
);

OAI22xp5_ASAP7_75t_L g2629 ( 
.A1(n_2550),
.A2(n_2460),
.B1(n_2497),
.B2(n_2484),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2517),
.B(n_2438),
.Y(n_2630)
);

AOI22x1_ASAP7_75t_SL g2631 ( 
.A1(n_2507),
.A2(n_2369),
.B1(n_2335),
.B2(n_2428),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2583),
.B(n_2565),
.Y(n_2632)
);

AND2x4_ASAP7_75t_L g2633 ( 
.A(n_2541),
.B(n_2346),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2509),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2515),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2528),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2569),
.B(n_2414),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2609),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2613),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2614),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2576),
.B(n_2428),
.Y(n_2641)
);

OAI21xp33_ASAP7_75t_L g2642 ( 
.A1(n_2502),
.A2(n_2618),
.B(n_2570),
.Y(n_2642)
);

AOI21xp5_ASAP7_75t_L g2643 ( 
.A1(n_2534),
.A2(n_2440),
.B(n_2439),
.Y(n_2643)
);

AOI22xp33_ASAP7_75t_L g2644 ( 
.A1(n_2562),
.A2(n_2420),
.B1(n_2340),
.B2(n_2393),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2531),
.Y(n_2645)
);

OAI21xp5_ASAP7_75t_L g2646 ( 
.A1(n_2549),
.A2(n_2396),
.B(n_2461),
.Y(n_2646)
);

AOI222xp33_ASAP7_75t_L g2647 ( 
.A1(n_2606),
.A2(n_2523),
.B1(n_2597),
.B2(n_2525),
.C1(n_2526),
.C2(n_2556),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2533),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2537),
.Y(n_2649)
);

AOI222xp33_ASAP7_75t_L g2650 ( 
.A1(n_2602),
.A2(n_2424),
.B1(n_2405),
.B2(n_2415),
.C1(n_2422),
.C2(n_2421),
.Y(n_2650)
);

OAI22xp5_ASAP7_75t_L g2651 ( 
.A1(n_2572),
.A2(n_2462),
.B1(n_2480),
.B2(n_2463),
.Y(n_2651)
);

OAI22xp5_ASAP7_75t_L g2652 ( 
.A1(n_2592),
.A2(n_2483),
.B1(n_2488),
.B2(n_2404),
.Y(n_2652)
);

AND2x2_ASAP7_75t_L g2653 ( 
.A(n_2522),
.B(n_2406),
.Y(n_2653)
);

INVx1_ASAP7_75t_SL g2654 ( 
.A(n_2532),
.Y(n_2654)
);

NOR2xp33_ASAP7_75t_SL g2655 ( 
.A(n_2536),
.B(n_2425),
.Y(n_2655)
);

OAI22xp33_ASAP7_75t_L g2656 ( 
.A1(n_2625),
.A2(n_2392),
.B1(n_2403),
.B2(n_2385),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2544),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2601),
.B(n_2384),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2607),
.B(n_2434),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2530),
.B(n_397),
.Y(n_2660)
);

INVx1_ASAP7_75t_SL g2661 ( 
.A(n_2599),
.Y(n_2661)
);

INVx1_ASAP7_75t_SL g2662 ( 
.A(n_2605),
.Y(n_2662)
);

OAI221xp5_ASAP7_75t_L g2663 ( 
.A1(n_2558),
.A2(n_2508),
.B1(n_2554),
.B2(n_2521),
.C(n_2542),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2510),
.B(n_398),
.Y(n_2664)
);

INVx3_ASAP7_75t_L g2665 ( 
.A(n_2551),
.Y(n_2665)
);

NOR3xp33_ASAP7_75t_L g2666 ( 
.A(n_2516),
.B(n_399),
.C(n_400),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2547),
.Y(n_2667)
);

AND2x2_ASAP7_75t_L g2668 ( 
.A(n_2548),
.B(n_399),
.Y(n_2668)
);

NOR2xp33_ASAP7_75t_L g2669 ( 
.A(n_2511),
.B(n_400),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2552),
.Y(n_2670)
);

AOI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2551),
.A2(n_403),
.B1(n_401),
.B2(n_402),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2573),
.Y(n_2672)
);

OA22x2_ASAP7_75t_L g2673 ( 
.A1(n_2588),
.A2(n_403),
.B1(n_401),
.B2(n_402),
.Y(n_2673)
);

OAI22xp33_ASAP7_75t_SL g2674 ( 
.A1(n_2612),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.Y(n_2674)
);

NAND3xp33_ASAP7_75t_L g2675 ( 
.A(n_2561),
.B(n_405),
.C(n_406),
.Y(n_2675)
);

OAI22xp5_ASAP7_75t_L g2676 ( 
.A1(n_2506),
.A2(n_410),
.B1(n_407),
.B2(n_409),
.Y(n_2676)
);

AOI222xp33_ASAP7_75t_L g2677 ( 
.A1(n_2603),
.A2(n_409),
.B1(n_410),
.B2(n_412),
.C1(n_413),
.C2(n_414),
.Y(n_2677)
);

INVx1_ASAP7_75t_SL g2678 ( 
.A(n_2608),
.Y(n_2678)
);

OAI21xp33_ASAP7_75t_L g2679 ( 
.A1(n_2503),
.A2(n_412),
.B(n_413),
.Y(n_2679)
);

O2A1O1Ixp33_ASAP7_75t_L g2680 ( 
.A1(n_2519),
.A2(n_416),
.B(n_414),
.C(n_415),
.Y(n_2680)
);

NAND3xp33_ASAP7_75t_SL g2681 ( 
.A(n_2513),
.B(n_415),
.C(n_416),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2584),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2586),
.Y(n_2683)
);

OR2x2_ASAP7_75t_L g2684 ( 
.A(n_2567),
.B(n_418),
.Y(n_2684)
);

OAI221xp5_ASAP7_75t_L g2685 ( 
.A1(n_2610),
.A2(n_421),
.B1(n_418),
.B2(n_419),
.C(n_423),
.Y(n_2685)
);

INVx1_ASAP7_75t_SL g2686 ( 
.A(n_2621),
.Y(n_2686)
);

HB1xp67_ASAP7_75t_L g2687 ( 
.A(n_2654),
.Y(n_2687)
);

AOI21xp5_ASAP7_75t_L g2688 ( 
.A1(n_2642),
.A2(n_2535),
.B(n_2529),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2684),
.Y(n_2689)
);

INVxp67_ASAP7_75t_L g2690 ( 
.A(n_2631),
.Y(n_2690)
);

AND2x2_ASAP7_75t_L g2691 ( 
.A(n_2633),
.B(n_2505),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2632),
.Y(n_2692)
);

AOI22xp33_ASAP7_75t_L g2693 ( 
.A1(n_2647),
.A2(n_2655),
.B1(n_2666),
.B2(n_2663),
.Y(n_2693)
);

OAI221xp5_ASAP7_75t_SL g2694 ( 
.A1(n_2680),
.A2(n_2679),
.B1(n_2628),
.B2(n_2659),
.C(n_2677),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2633),
.B(n_2568),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2627),
.Y(n_2696)
);

AOI22xp5_ASAP7_75t_L g2697 ( 
.A1(n_2656),
.A2(n_2546),
.B1(n_2543),
.B2(n_2539),
.Y(n_2697)
);

OAI32xp33_ASAP7_75t_L g2698 ( 
.A1(n_2626),
.A2(n_2564),
.A3(n_2581),
.B1(n_2577),
.B2(n_2559),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2638),
.Y(n_2699)
);

OAI21xp33_ASAP7_75t_L g2700 ( 
.A1(n_2665),
.A2(n_2590),
.B(n_2589),
.Y(n_2700)
);

AOI221x1_ASAP7_75t_L g2701 ( 
.A1(n_2674),
.A2(n_2520),
.B1(n_2518),
.B2(n_2524),
.C(n_2504),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2637),
.Y(n_2702)
);

INVxp67_ASAP7_75t_L g2703 ( 
.A(n_2630),
.Y(n_2703)
);

AOI221xp5_ASAP7_75t_L g2704 ( 
.A1(n_2629),
.A2(n_2593),
.B1(n_2596),
.B2(n_2595),
.C(n_2591),
.Y(n_2704)
);

OAI221xp5_ASAP7_75t_L g2705 ( 
.A1(n_2646),
.A2(n_2611),
.B1(n_2622),
.B2(n_2615),
.C(n_2604),
.Y(n_2705)
);

AOI21xp33_ASAP7_75t_L g2706 ( 
.A1(n_2686),
.A2(n_2624),
.B(n_2623),
.Y(n_2706)
);

AND2x2_ASAP7_75t_SL g2707 ( 
.A(n_2641),
.B(n_2553),
.Y(n_2707)
);

AOI21xp5_ASAP7_75t_L g2708 ( 
.A1(n_2643),
.A2(n_2616),
.B(n_2585),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2639),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2640),
.Y(n_2710)
);

OAI32xp33_ASAP7_75t_L g2711 ( 
.A1(n_2675),
.A2(n_2617),
.A3(n_2580),
.B1(n_2587),
.B2(n_2578),
.Y(n_2711)
);

BUFx2_ASAP7_75t_L g2712 ( 
.A(n_2653),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2661),
.B(n_2662),
.Y(n_2713)
);

NOR2xp33_ASAP7_75t_L g2714 ( 
.A(n_2678),
.B(n_2538),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2650),
.B(n_2566),
.Y(n_2715)
);

AOI21xp5_ASAP7_75t_L g2716 ( 
.A1(n_2681),
.A2(n_2619),
.B(n_2557),
.Y(n_2716)
);

AOI21xp5_ASAP7_75t_L g2717 ( 
.A1(n_2652),
.A2(n_2582),
.B(n_2574),
.Y(n_2717)
);

AOI22xp5_ASAP7_75t_L g2718 ( 
.A1(n_2651),
.A2(n_2582),
.B1(n_2575),
.B2(n_2545),
.Y(n_2718)
);

INVx1_ASAP7_75t_SL g2719 ( 
.A(n_2660),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2668),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2687),
.B(n_2636),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2713),
.Y(n_2722)
);

OR2x2_ASAP7_75t_L g2723 ( 
.A(n_2719),
.B(n_2712),
.Y(n_2723)
);

XNOR2xp5_ASAP7_75t_L g2724 ( 
.A(n_2707),
.B(n_2673),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2689),
.Y(n_2725)
);

AOI21xp5_ASAP7_75t_L g2726 ( 
.A1(n_2693),
.A2(n_2658),
.B(n_2676),
.Y(n_2726)
);

OAI22xp5_ASAP7_75t_L g2727 ( 
.A1(n_2690),
.A2(n_2671),
.B1(n_2644),
.B2(n_2685),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2696),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2720),
.Y(n_2729)
);

INVxp33_ASAP7_75t_L g2730 ( 
.A(n_2714),
.Y(n_2730)
);

OAI22xp33_ASAP7_75t_SL g2731 ( 
.A1(n_2694),
.A2(n_2634),
.B1(n_2645),
.B2(n_2635),
.Y(n_2731)
);

NOR2x1_ASAP7_75t_L g2732 ( 
.A(n_2692),
.B(n_2669),
.Y(n_2732)
);

AOI21xp5_ASAP7_75t_L g2733 ( 
.A1(n_2708),
.A2(n_2664),
.B(n_2649),
.Y(n_2733)
);

OAI32xp33_ASAP7_75t_L g2734 ( 
.A1(n_2715),
.A2(n_2667),
.A3(n_2670),
.B1(n_2657),
.B2(n_2648),
.Y(n_2734)
);

NOR2x1_ASAP7_75t_L g2735 ( 
.A(n_2702),
.B(n_2571),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2695),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2691),
.Y(n_2737)
);

NOR2xp33_ASAP7_75t_L g2738 ( 
.A(n_2698),
.B(n_2563),
.Y(n_2738)
);

NOR2xp33_ASAP7_75t_L g2739 ( 
.A(n_2703),
.B(n_2672),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2723),
.Y(n_2740)
);

AOI22xp33_ASAP7_75t_L g2741 ( 
.A1(n_2731),
.A2(n_2727),
.B1(n_2738),
.B2(n_2726),
.Y(n_2741)
);

AOI221xp5_ASAP7_75t_L g2742 ( 
.A1(n_2734),
.A2(n_2705),
.B1(n_2706),
.B2(n_2688),
.C(n_2704),
.Y(n_2742)
);

AOI222xp33_ASAP7_75t_L g2743 ( 
.A1(n_2724),
.A2(n_2700),
.B1(n_2711),
.B2(n_2710),
.C1(n_2709),
.C2(n_2699),
.Y(n_2743)
);

AOI211xp5_ASAP7_75t_L g2744 ( 
.A1(n_2730),
.A2(n_2717),
.B(n_2716),
.C(n_2697),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2737),
.B(n_2718),
.Y(n_2745)
);

NOR3xp33_ASAP7_75t_L g2746 ( 
.A(n_2722),
.B(n_2721),
.C(n_2732),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2736),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2735),
.Y(n_2748)
);

AOI221xp5_ASAP7_75t_L g2749 ( 
.A1(n_2742),
.A2(n_2733),
.B1(n_2739),
.B2(n_2728),
.C(n_2725),
.Y(n_2749)
);

XNOR2xp5_ASAP7_75t_L g2750 ( 
.A(n_2744),
.B(n_2697),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2748),
.B(n_2729),
.Y(n_2751)
);

AOI221xp5_ASAP7_75t_L g2752 ( 
.A1(n_2741),
.A2(n_2683),
.B1(n_2682),
.B2(n_2540),
.C(n_2598),
.Y(n_2752)
);

AOI21xp33_ASAP7_75t_L g2753 ( 
.A1(n_2743),
.A2(n_2740),
.B(n_2745),
.Y(n_2753)
);

AOI221xp5_ASAP7_75t_L g2754 ( 
.A1(n_2746),
.A2(n_2527),
.B1(n_2560),
.B2(n_2555),
.C(n_2579),
.Y(n_2754)
);

AOI221xp5_ASAP7_75t_SL g2755 ( 
.A1(n_2747),
.A2(n_2594),
.B1(n_2620),
.B2(n_2701),
.C(n_423),
.Y(n_2755)
);

AOI21xp5_ASAP7_75t_L g2756 ( 
.A1(n_2744),
.A2(n_419),
.B(n_421),
.Y(n_2756)
);

AOI22xp5_ASAP7_75t_L g2757 ( 
.A1(n_2750),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_2757)
);

HB1xp67_ASAP7_75t_L g2758 ( 
.A(n_2751),
.Y(n_2758)
);

O2A1O1Ixp33_ASAP7_75t_L g2759 ( 
.A1(n_2753),
.A2(n_428),
.B(n_426),
.C(n_427),
.Y(n_2759)
);

OAI21xp33_ASAP7_75t_L g2760 ( 
.A1(n_2752),
.A2(n_427),
.B(n_428),
.Y(n_2760)
);

OAI22xp5_ASAP7_75t_L g2761 ( 
.A1(n_2749),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2758),
.Y(n_2762)
);

NOR2x1_ASAP7_75t_L g2763 ( 
.A(n_2759),
.B(n_2756),
.Y(n_2763)
);

NAND2x1p5_ASAP7_75t_L g2764 ( 
.A(n_2762),
.B(n_2757),
.Y(n_2764)
);

AOI22xp33_ASAP7_75t_L g2765 ( 
.A1(n_2764),
.A2(n_2761),
.B1(n_2763),
.B2(n_2760),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2765),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2766),
.Y(n_2767)
);

OA21x2_ASAP7_75t_L g2768 ( 
.A1(n_2766),
.A2(n_2755),
.B(n_2754),
.Y(n_2768)
);

AO22x2_ASAP7_75t_L g2769 ( 
.A1(n_2767),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.Y(n_2769)
);

XNOR2xp5_ASAP7_75t_L g2770 ( 
.A(n_2768),
.B(n_432),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2770),
.Y(n_2771)
);

AOI21xp5_ASAP7_75t_L g2772 ( 
.A1(n_2771),
.A2(n_2769),
.B(n_434),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2772),
.Y(n_2773)
);

OAI21xp5_ASAP7_75t_L g2774 ( 
.A1(n_2772),
.A2(n_434),
.B(n_435),
.Y(n_2774)
);

AOI22xp33_ASAP7_75t_L g2775 ( 
.A1(n_2773),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2774),
.Y(n_2776)
);

OAI221xp5_ASAP7_75t_R g2777 ( 
.A1(n_2775),
.A2(n_439),
.B1(n_436),
.B2(n_438),
.C(n_440),
.Y(n_2777)
);

AOI211xp5_ASAP7_75t_L g2778 ( 
.A1(n_2777),
.A2(n_2776),
.B(n_439),
.C(n_671),
.Y(n_2778)
);


endmodule