module fake_jpeg_23370_n_349 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_48),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_49),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_46),
.Y(n_63)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_24),
.B(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_53),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_64),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_24),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_50),
.Y(n_81)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_38),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_28),
.B1(n_34),
.B2(n_29),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_72),
.A2(n_28),
.B1(n_42),
.B2(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_76),
.Y(n_107)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_75),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_114)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_46),
.A3(n_41),
.B1(n_42),
.B2(n_29),
.Y(n_77)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_77),
.B(n_38),
.C(n_23),
.Y(n_130)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_79),
.Y(n_108)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_88),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_60),
.A2(n_50),
.B1(n_44),
.B2(n_46),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_93),
.B1(n_41),
.B2(n_39),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_28),
.B1(n_20),
.B2(n_45),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_85),
.A2(n_22),
.B1(n_36),
.B2(n_19),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_34),
.B1(n_22),
.B2(n_18),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_90),
.Y(n_135)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx6_ASAP7_75t_SL g91 ( 
.A(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_91),
.Y(n_112)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_60),
.A2(n_44),
.B1(n_51),
.B2(n_43),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_62),
.B(n_45),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_97),
.Y(n_120)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_55),
.B(n_39),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_101),
.Y(n_121)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_59),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_103),
.Y(n_132)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_67),
.A2(n_18),
.B1(n_21),
.B2(n_36),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_118),
.Y(n_141)
);

NAND2xp33_ASAP7_75t_SL g115 ( 
.A(n_77),
.B(n_58),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_130),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_43),
.B1(n_53),
.B2(n_21),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_125),
.B1(n_102),
.B2(n_95),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_49),
.B(n_19),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_129),
.B1(n_102),
.B2(n_78),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_43),
.B1(n_51),
.B2(n_49),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_127),
.Y(n_139)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_84),
.A2(n_71),
.B1(n_70),
.B2(n_64),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_133),
.Y(n_142)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_0),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_99),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_137),
.A2(n_159),
.B1(n_27),
.B2(n_23),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_132),
.B1(n_131),
.B2(n_127),
.Y(n_175)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_140),
.B(n_145),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_120),
.B(n_73),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_151),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_104),
.Y(n_144)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_148),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_110),
.A2(n_90),
.B1(n_76),
.B2(n_97),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_153),
.B1(n_157),
.B2(n_158),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_116),
.Y(n_148)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_150),
.Y(n_182)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_94),
.C(n_101),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_109),
.B1(n_130),
.B2(n_115),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_166),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_96),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_156),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_109),
.A2(n_99),
.B1(n_92),
.B2(n_86),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_130),
.A2(n_74),
.B1(n_100),
.B2(n_98),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_88),
.B1(n_79),
.B2(n_86),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_160),
.A2(n_128),
.B1(n_124),
.B2(n_113),
.Y(n_184)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_101),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_164),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_80),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_152),
.C(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_83),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_132),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_165),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_111),
.B(n_56),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_121),
.B1(n_111),
.B2(n_135),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_169),
.A2(n_175),
.B1(n_181),
.B2(n_149),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_166),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_170),
.Y(n_205)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_119),
.A3(n_121),
.B1(n_136),
.B2(n_134),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_145),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_178),
.C(n_188),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_189),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_47),
.C(n_126),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_128),
.B1(n_124),
.B2(n_113),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_184),
.A2(n_197),
.B1(n_26),
.B2(n_17),
.Y(n_226)
);

HAxp5_ASAP7_75t_SL g185 ( 
.A(n_151),
.B(n_47),
.CON(n_185),
.SN(n_185)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_185),
.A2(n_161),
.B1(n_148),
.B2(n_146),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_47),
.C(n_37),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_141),
.B(n_27),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_193),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_37),
.B(n_35),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_195),
.B(n_155),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_27),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_147),
.B(n_35),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_194),
.B(n_9),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_30),
.B(n_31),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_27),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_199),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_158),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_137),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_10),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_140),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_200),
.Y(n_220)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_167),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_213),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_203),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_204),
.A2(n_206),
.B1(n_217),
.B2(n_179),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_207),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_150),
.Y(n_208)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_172),
.B(n_23),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_188),
.C(n_199),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_159),
.Y(n_210)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_230),
.Y(n_233)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_191),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_224),
.Y(n_238)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_185),
.A2(n_183),
.B(n_170),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_222),
.B1(n_223),
.B2(n_226),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_169),
.A2(n_148),
.B1(n_32),
.B2(n_23),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_216),
.A2(n_229),
.B1(n_197),
.B2(n_186),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_10),
.Y(n_219)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_183),
.A2(n_32),
.B1(n_17),
.B2(n_26),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_180),
.A2(n_32),
.B1(n_17),
.B2(n_26),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_227),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_192),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_195),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_178),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_1),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_189),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_221),
.B(n_193),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_232),
.B(n_250),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_190),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_236),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g235 ( 
.A(n_218),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_246),
.Y(n_275)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_168),
.C(n_180),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_250),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_251),
.B1(n_216),
.B2(n_206),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_204),
.A2(n_224),
.B1(n_227),
.B2(n_207),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_248),
.A2(n_215),
.B1(n_205),
.B2(n_220),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_168),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_171),
.B1(n_174),
.B2(n_173),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_252),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_208),
.B(n_194),
.Y(n_254)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_254),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_279),
.B1(n_254),
.B2(n_242),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_257),
.Y(n_261)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_256),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_263),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_255),
.A2(n_205),
.B1(n_202),
.B2(n_215),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_265),
.A2(n_271),
.B1(n_233),
.B2(n_244),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_248),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_266),
.A2(n_4),
.B(n_5),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_237),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_268),
.B(n_273),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_243),
.A2(n_211),
.B1(n_213),
.B2(n_231),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_274),
.B1(n_246),
.B2(n_247),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_201),
.B1(n_223),
.B2(n_230),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_243),
.A2(n_229),
.B1(n_209),
.B2(n_3),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_272),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_252),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_15),
.Y(n_279)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_241),
.C(n_236),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_282),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_232),
.C(n_245),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_234),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_290),
.Y(n_299)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_240),
.C(n_238),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_293),
.Y(n_304)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_265),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_291),
.B(n_15),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_264),
.A2(n_1),
.B(n_2),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_292),
.A2(n_295),
.B(n_276),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_1),
.C(n_3),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_262),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_295),
.Y(n_303)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

AOI21xp33_ASAP7_75t_L g302 ( 
.A1(n_286),
.A2(n_276),
.B(n_275),
.Y(n_302)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_305),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_259),
.Y(n_305)
);

OAI221xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_260),
.B1(n_266),
.B2(n_267),
.C(n_12),
.Y(n_307)
);

NOR3xp33_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_293),
.C(n_306),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_287),
.A2(n_266),
.B(n_267),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_294),
.B(n_285),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_292),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_14),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_312),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_14),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_289),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_317),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_318),
.C(n_324),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_321),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_281),
.C(n_290),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_280),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_289),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_299),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_288),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_308),
.B1(n_320),
.B2(n_314),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_5),
.C(n_6),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_297),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_327),
.A2(n_328),
.B(n_329),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_304),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_321),
.A2(n_309),
.B(n_312),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_13),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_323),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_11),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_334),
.B(n_335),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_331),
.A2(n_11),
.B(n_5),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_336),
.A2(n_338),
.B(n_340),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_4),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_334),
.C(n_339),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_325),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_342),
.B(n_7),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_341),
.B(n_331),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_344),
.B(n_345),
.Y(n_346)
);

NOR2x1p5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_343),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_7),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_8),
.Y(n_349)
);


endmodule