module fake_jpeg_26451_n_295 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_32),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_38),
.Y(n_45)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_30),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_8),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_29),
.Y(n_48)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_19),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_56),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_17),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_25),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_40),
.B(n_39),
.C(n_36),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_24),
.B1(n_19),
.B2(n_25),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_41),
.B1(n_18),
.B2(n_20),
.Y(n_84)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_32),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_75),
.C(n_77),
.Y(n_102)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_63),
.B(n_69),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_34),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_30),
.B1(n_33),
.B2(n_24),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_70),
.A2(n_72),
.B1(n_23),
.B2(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_40),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_30),
.B1(n_33),
.B2(n_25),
.Y(n_72)
);

FAx1_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_39),
.CI(n_36),
.CON(n_73),
.SN(n_73)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_74),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_26),
.Y(n_74)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_39),
.C(n_36),
.Y(n_75)
);

OR2x2_ASAP7_75t_SL g76 ( 
.A(n_48),
.B(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_81),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_36),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_51),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_41),
.B1(n_21),
.B2(n_23),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_84),
.B1(n_90),
.B2(n_21),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_17),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_29),
.Y(n_115)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_55),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_18),
.B(n_22),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_46),
.B1(n_43),
.B2(n_54),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_41),
.B1(n_20),
.B2(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_93),
.B(n_105),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_108),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_50),
.B1(n_54),
.B2(n_46),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_90),
.B1(n_87),
.B2(n_61),
.Y(n_120)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_114),
.B1(n_60),
.B2(n_85),
.Y(n_130)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_110),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_55),
.C(n_44),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_111),
.C(n_112),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_67),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_55),
.C(n_17),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_55),
.C(n_31),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_117),
.Y(n_119)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_120),
.A2(n_135),
.B1(n_140),
.B2(n_146),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_133),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_117),
.A2(n_66),
.B1(n_88),
.B2(n_72),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_123),
.A2(n_125),
.B1(n_129),
.B2(n_130),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_132),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_114),
.A2(n_88),
.B1(n_70),
.B2(n_71),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_77),
.B1(n_63),
.B2(n_69),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_126),
.A2(n_135),
.B1(n_138),
.B2(n_140),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_77),
.B(n_86),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_62),
.B1(n_86),
.B2(n_61),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_68),
.B1(n_65),
.B2(n_64),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_62),
.Y(n_132)
);

INVxp67_ASAP7_75t_SL g133 ( 
.A(n_100),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_96),
.A2(n_74),
.B1(n_68),
.B2(n_64),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_65),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_141),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_76),
.B1(n_42),
.B2(n_31),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_27),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_144),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_91),
.A2(n_42),
.B1(n_31),
.B2(n_27),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_31),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_42),
.B1(n_27),
.B2(n_28),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_27),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_99),
.A2(n_98),
.B1(n_110),
.B2(n_97),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_28),
.C(n_42),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_116),
.C(n_113),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_92),
.B(n_0),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_124),
.Y(n_172)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_159),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_92),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_152),
.B(n_155),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_97),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_153),
.A2(n_142),
.B(n_136),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_154),
.B(n_162),
.C(n_9),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_118),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_118),
.B1(n_101),
.B2(n_95),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_173),
.B1(n_176),
.B2(n_1),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_28),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_144),
.Y(n_185)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_101),
.C(n_95),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_177),
.B1(n_125),
.B2(n_141),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_121),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_166),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_137),
.Y(n_166)
);

OAI32xp33_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_28),
.A3(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_168)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_107),
.Y(n_170)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_172),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_128),
.A2(n_107),
.B1(n_28),
.B2(n_2),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_143),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_179),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_126),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_1),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_177),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_143),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_180),
.A2(n_182),
.B(n_190),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_129),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_204),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_189),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_174),
.A2(n_136),
.B(n_123),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_191),
.A2(n_169),
.B1(n_161),
.B2(n_178),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_193),
.B(n_195),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_174),
.A2(n_158),
.B(n_151),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_197),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_153),
.A2(n_139),
.B(n_4),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_154),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_12),
.C(n_11),
.Y(n_226)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_201),
.Y(n_210)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_202),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_15),
.Y(n_203)
);

NOR3xp33_ASAP7_75t_SL g220 ( 
.A(n_203),
.B(n_7),
.C(n_12),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_158),
.A2(n_153),
.B1(n_160),
.B2(n_171),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_150),
.C(n_10),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_206),
.A2(n_207),
.B1(n_211),
.B2(n_183),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_204),
.A2(n_169),
.B1(n_159),
.B2(n_160),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_196),
.A2(n_168),
.B1(n_157),
.B2(n_150),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_213),
.B(n_11),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_10),
.C(n_14),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_217),
.C(n_219),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_15),
.C(n_8),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_14),
.C(n_7),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_203),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_199),
.B1(n_188),
.B2(n_187),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_13),
.C(n_7),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_226),
.C(n_195),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_228),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_214),
.B(n_186),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_184),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_194),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_233),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_190),
.Y(n_233)
);

AO22x1_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_196),
.B1(n_202),
.B2(n_182),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_236),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_222),
.A2(n_182),
.B(n_180),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_237),
.B(n_241),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_242),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_216),
.A2(n_189),
.B1(n_184),
.B2(n_200),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_192),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_226),
.B(n_192),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_243),
.A2(n_212),
.B1(n_210),
.B2(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_238),
.A2(n_224),
.B1(n_207),
.B2(n_221),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_250),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_206),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_249),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_232),
.B(n_211),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_240),
.A2(n_209),
.B1(n_213),
.B2(n_223),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_219),
.C(n_217),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_237),
.C(n_234),
.Y(n_258)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_230),
.B(n_236),
.CI(n_235),
.CON(n_253),
.SN(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_253),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_249),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_234),
.C(n_227),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_263),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_255),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_253),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_235),
.Y(n_262)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_256),
.Y(n_263)
);

AO21x1_ASAP7_75t_L g265 ( 
.A1(n_255),
.A2(n_220),
.B(n_12),
.Y(n_265)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_6),
.C(n_251),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_268),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_6),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_270),
.B(n_275),
.Y(n_282)
);

AOI221xp5_ASAP7_75t_L g272 ( 
.A1(n_267),
.A2(n_250),
.B1(n_254),
.B2(n_246),
.C(n_247),
.Y(n_272)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_272),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_248),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_244),
.C(n_253),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_276),
.B(n_278),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_281),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_276),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_262),
.B(n_263),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_283),
.A2(n_273),
.B(n_259),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_284),
.B(n_274),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_286),
.Y(n_289)
);

AND2x2_ASAP7_75t_SL g288 ( 
.A(n_279),
.B(n_270),
.Y(n_288)
);

NOR3xp33_ASAP7_75t_SL g290 ( 
.A(n_288),
.B(n_282),
.C(n_269),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_265),
.B(n_287),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_291),
.A2(n_269),
.B(n_289),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_292),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_275),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_244),
.Y(n_295)
);


endmodule