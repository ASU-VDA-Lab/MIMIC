module fake_netlist_5_379_n_1892 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1892);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1892;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1865;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g189 ( 
.A(n_42),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_96),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_133),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_12),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_153),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_63),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_102),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_73),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_121),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_92),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_115),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_98),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_155),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_13),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_72),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_75),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_119),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_130),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_150),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_125),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_25),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_62),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_25),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_74),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_27),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_160),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_2),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_136),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_114),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_18),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_186),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_39),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_169),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_173),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_27),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_10),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_62),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_176),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_156),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_59),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_87),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_57),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_158),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_34),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_124),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_109),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_1),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_117),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_59),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_97),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_49),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_131),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_143),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_45),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_13),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_69),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_100),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_57),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_187),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_129),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_144),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_10),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_81),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_104),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_157),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_36),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_167),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_20),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_31),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_90),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_185),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_17),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_79),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_64),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_24),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_99),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_180),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_33),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_18),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_171),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_137),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_54),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_61),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_37),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_120),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_149),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_105),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_110),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_175),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_139),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_70),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_78),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_30),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_15),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_56),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_123),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_31),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_45),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_108),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_4),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_85),
.Y(n_295)
);

BUFx8_ASAP7_75t_SL g296 ( 
.A(n_111),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_88),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_2),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_159),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_14),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_21),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_145),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_4),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_127),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_16),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_181),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_17),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_141),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_140),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_147),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_3),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_36),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_54),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_26),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_68),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_5),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_15),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_28),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_83),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_8),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_6),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_38),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_61),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_29),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_39),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_8),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_165),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_49),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_82),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_11),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_43),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_174),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_16),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_146),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_19),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_46),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_46),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_154),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_1),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_11),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_101),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_178),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_80),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_134),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_135),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_41),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_188),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_12),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_116),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_0),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_132),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_152),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_41),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_93),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_161),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_103),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_89),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_3),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_30),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_142),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_122),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_56),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_29),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_64),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_95),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_94),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_112),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_126),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_71),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_9),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_26),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_32),
.Y(n_372)
);

INVxp33_ASAP7_75t_R g373 ( 
.A(n_164),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_168),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_67),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_48),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_42),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_53),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_218),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_200),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_206),
.Y(n_381)
);

INVxp33_ASAP7_75t_SL g382 ( 
.A(n_207),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_296),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_254),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_231),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_235),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_211),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_218),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_192),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_257),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_218),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_290),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_315),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_240),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_242),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_218),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_218),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_243),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_246),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_341),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_247),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_267),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_233),
.B(n_0),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_250),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_243),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_253),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_283),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_243),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_334),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_243),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_259),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_342),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_374),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_243),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_264),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_295),
.B(n_5),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_265),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_R g418 ( 
.A(n_190),
.B(n_128),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_256),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_270),
.Y(n_420)
);

INVxp33_ASAP7_75t_L g421 ( 
.A(n_189),
.Y(n_421)
);

BUFx6f_ASAP7_75t_SL g422 ( 
.A(n_267),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_256),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_256),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_205),
.B(n_6),
.Y(n_425)
);

INVxp33_ASAP7_75t_SL g426 ( 
.A(n_207),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_256),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_256),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_321),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_321),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_199),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_321),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_271),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_205),
.B(n_7),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_321),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_280),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_281),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_366),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_321),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_282),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_286),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_330),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_194),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_192),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_293),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_297),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_302),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_225),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_366),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_304),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_228),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_230),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_214),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_306),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_308),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_285),
.B(n_329),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_285),
.B(n_7),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_241),
.Y(n_458)
);

CKINVDCx14_ASAP7_75t_R g459 ( 
.A(n_192),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_252),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_309),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_269),
.B(n_9),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_278),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_276),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_277),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_310),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_278),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_319),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_327),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_287),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_214),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_288),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_329),
.B(n_14),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_379),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_408),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_379),
.Y(n_476)
);

OA21x2_ASAP7_75t_L g477 ( 
.A1(n_456),
.A2(n_391),
.B(n_388),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_449),
.B(n_191),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_388),
.B(n_391),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_402),
.B(n_216),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_396),
.B(n_191),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_396),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_397),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_403),
.B(n_221),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_SL g485 ( 
.A(n_462),
.B(n_216),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_397),
.B(n_195),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_398),
.B(n_201),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_402),
.B(n_203),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_398),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_380),
.A2(n_223),
.B1(n_234),
.B2(n_238),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_442),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_405),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_405),
.B(n_232),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g494 ( 
.A(n_457),
.B(n_229),
.C(n_236),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_R g495 ( 
.A(n_382),
.B(n_215),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_410),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_410),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_414),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_414),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_419),
.B(n_193),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_419),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_423),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_423),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_424),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_424),
.B(n_251),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_438),
.B(n_255),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_427),
.Y(n_507)
);

CKINVDCx8_ASAP7_75t_R g508 ( 
.A(n_383),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_427),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_389),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_428),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_428),
.B(n_193),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_429),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_418),
.B(n_278),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_429),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_463),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_430),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_430),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_438),
.B(n_261),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_432),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_432),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_435),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_435),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_439),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_439),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_443),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_425),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_443),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_434),
.Y(n_529)
);

NAND2xp33_ASAP7_75t_L g530 ( 
.A(n_462),
.B(n_258),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_448),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_448),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_381),
.B(n_387),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_451),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_451),
.Y(n_535)
);

INVx6_ASAP7_75t_L g536 ( 
.A(n_422),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_452),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_452),
.Y(n_538)
);

BUFx12f_ASAP7_75t_L g539 ( 
.A(n_385),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_458),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_458),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_460),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_426),
.B(n_384),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_460),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_L g545 ( 
.A(n_464),
.B(n_258),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_464),
.Y(n_546)
);

OAI21x1_ASAP7_75t_L g547 ( 
.A1(n_473),
.A2(n_279),
.B(n_275),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_465),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_465),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_470),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_453),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_470),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_484),
.A2(n_441),
.B1(n_454),
.B2(n_446),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_539),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_531),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_477),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_531),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_476),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_491),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_488),
.B(n_407),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_529),
.B(n_386),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_531),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_529),
.A2(n_409),
.B1(n_416),
.B2(n_291),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_527),
.B(n_258),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_531),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_476),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_475),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_475),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_475),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_475),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_474),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_L g572 ( 
.A(n_527),
.B(n_258),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_528),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_529),
.B(n_394),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_528),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_480),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_486),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_527),
.B(n_258),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_534),
.Y(n_579)
);

BUFx4f_ASAP7_75t_L g580 ( 
.A(n_527),
.Y(n_580)
);

AO22x2_ASAP7_75t_L g581 ( 
.A1(n_494),
.A2(n_314),
.B1(n_377),
.B2(n_300),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_484),
.B(n_395),
.Y(n_582)
);

BUFx4f_ASAP7_75t_L g583 ( 
.A(n_527),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_491),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_534),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_529),
.B(n_399),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_543),
.B(n_401),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_537),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_551),
.Y(n_589)
);

OAI21xp33_ASAP7_75t_SL g590 ( 
.A1(n_547),
.A2(n_303),
.B(n_301),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_486),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_482),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_480),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_482),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_527),
.B(n_404),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_533),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_L g597 ( 
.A(n_527),
.B(n_274),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_476),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_499),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_527),
.B(n_478),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_535),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_537),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_480),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_499),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_478),
.Y(n_605)
);

BUFx10_ASAP7_75t_L g606 ( 
.A(n_543),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_541),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_541),
.Y(n_608)
);

INVx5_ASAP7_75t_L g609 ( 
.A(n_474),
.Y(n_609)
);

OR2x6_ASAP7_75t_L g610 ( 
.A(n_539),
.B(n_536),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_499),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_535),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_501),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_514),
.B(n_406),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_535),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_544),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_530),
.B(n_411),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_510),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_544),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_501),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_501),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_486),
.B(n_274),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_514),
.B(n_415),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_502),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_546),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_510),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_546),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_550),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_536),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_530),
.B(n_417),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_486),
.B(n_487),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_486),
.B(n_274),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_488),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_550),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_535),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_488),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_474),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_502),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_552),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_502),
.Y(n_640)
);

OA22x2_ASAP7_75t_L g641 ( 
.A1(n_506),
.A2(n_471),
.B1(n_359),
.B2(n_311),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_506),
.B(n_274),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_485),
.A2(n_353),
.B1(n_371),
.B2(n_370),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_495),
.A2(n_440),
.B1(n_455),
.B2(n_466),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_518),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_L g646 ( 
.A(n_494),
.B(n_274),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_539),
.B(n_373),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_552),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_551),
.B(n_444),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_510),
.B(n_420),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_485),
.A2(n_333),
.B1(n_364),
.B2(n_316),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_533),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_518),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_487),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_487),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_474),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_487),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_506),
.B(n_472),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_518),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_487),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_493),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_520),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_481),
.B(n_433),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_SL g664 ( 
.A(n_508),
.B(n_431),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_481),
.B(n_436),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_493),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_500),
.B(n_437),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_493),
.Y(n_668)
);

BUFx8_ASAP7_75t_SL g669 ( 
.A(n_516),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_493),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_493),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_477),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_520),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_505),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_505),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_489),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_533),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_474),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_520),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_535),
.Y(n_680)
);

NAND3xp33_ASAP7_75t_L g681 ( 
.A(n_500),
.B(n_447),
.C(n_445),
.Y(n_681)
);

CKINVDCx11_ASAP7_75t_R g682 ( 
.A(n_508),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_489),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_519),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_505),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_505),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_505),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_496),
.Y(n_688)
);

AND2x6_ASAP7_75t_L g689 ( 
.A(n_519),
.B(n_299),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_519),
.B(n_472),
.Y(n_690)
);

NOR3xp33_ASAP7_75t_L g691 ( 
.A(n_490),
.B(n_467),
.C(n_331),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_496),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_512),
.B(n_450),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_498),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_535),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_L g696 ( 
.A1(n_495),
.A2(n_292),
.B1(n_340),
.B2(n_378),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_526),
.B(n_459),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_516),
.A2(n_469),
.B1(n_468),
.B2(n_461),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_512),
.B(n_237),
.Y(n_699)
);

AND2x6_ASAP7_75t_L g700 ( 
.A(n_549),
.B(n_299),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_516),
.B(n_422),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_535),
.B(n_299),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_498),
.Y(n_703)
);

NAND3xp33_ASAP7_75t_SL g704 ( 
.A(n_508),
.B(n_305),
.C(n_268),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_504),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_605),
.B(n_477),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_605),
.B(n_477),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_654),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_580),
.B(n_583),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_576),
.B(n_421),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_580),
.B(n_583),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_655),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_600),
.B(n_477),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_705),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_657),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_660),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_661),
.Y(n_717)
);

NOR2xp67_ASAP7_75t_L g718 ( 
.A(n_553),
.B(n_549),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_576),
.B(n_390),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_633),
.B(n_526),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_582),
.B(n_477),
.Y(n_721)
);

NOR2xp67_ASAP7_75t_L g722 ( 
.A(n_644),
.B(n_549),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_666),
.Y(n_723)
);

AND2x4_ASAP7_75t_SL g724 ( 
.A(n_610),
.B(n_647),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_633),
.B(n_526),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_683),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_636),
.B(n_532),
.Y(n_727)
);

AND2x6_ASAP7_75t_SL g728 ( 
.A(n_647),
.B(n_317),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_683),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_577),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_593),
.B(n_549),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_593),
.B(n_549),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_577),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_603),
.B(n_492),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_614),
.A2(n_623),
.B1(n_603),
.B2(n_561),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_580),
.B(n_547),
.Y(n_736)
);

NAND2xp33_ASAP7_75t_L g737 ( 
.A(n_595),
.B(n_332),
.Y(n_737)
);

AND2x4_ASAP7_75t_SL g738 ( 
.A(n_610),
.B(n_392),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_699),
.B(n_492),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_682),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_574),
.B(n_239),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_556),
.A2(n_547),
.B1(n_336),
.B2(n_318),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_SL g743 ( 
.A(n_554),
.B(n_393),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_591),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_668),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_688),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_636),
.B(n_492),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_705),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_670),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_684),
.B(n_663),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_684),
.B(n_492),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_650),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_690),
.B(n_532),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_618),
.B(n_490),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_556),
.A2(n_325),
.B1(n_339),
.B2(n_320),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_688),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_583),
.B(n_299),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_558),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_658),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_556),
.B(n_299),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_665),
.B(n_492),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_667),
.B(n_535),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_693),
.B(n_504),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_586),
.B(n_509),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_682),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_555),
.B(n_509),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_618),
.B(n_215),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_557),
.B(n_511),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_626),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_658),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_685),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_587),
.A2(n_400),
.B1(n_412),
.B2(n_413),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_672),
.B(n_244),
.Y(n_773)
);

AND2x6_ASAP7_75t_SL g774 ( 
.A(n_647),
.B(n_343),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_681),
.B(n_338),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_692),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_686),
.Y(n_777)
);

OAI221xp5_ASAP7_75t_L g778 ( 
.A1(n_563),
.A2(n_352),
.B1(n_355),
.B2(n_347),
.C(n_365),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_687),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_562),
.B(n_511),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_573),
.Y(n_781)
);

NOR2xp67_ASAP7_75t_L g782 ( 
.A(n_698),
.B(n_532),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_565),
.B(n_517),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_672),
.B(n_354),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_692),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_575),
.B(n_517),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_672),
.A2(n_346),
.B1(n_357),
.B2(n_220),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_579),
.B(n_523),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_560),
.B(n_538),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_626),
.B(n_220),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_585),
.B(n_523),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_694),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_696),
.B(n_196),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_588),
.Y(n_794)
);

NAND2xp33_ASAP7_75t_SL g795 ( 
.A(n_649),
.B(n_422),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_694),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_592),
.Y(n_797)
);

NOR3xp33_ASAP7_75t_L g798 ( 
.A(n_704),
.B(n_677),
.C(n_596),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_617),
.B(n_630),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_560),
.B(n_538),
.Y(n_800)
);

NAND3xp33_ASAP7_75t_L g801 ( 
.A(n_646),
.B(n_307),
.C(n_245),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_592),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_606),
.B(n_602),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_559),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_594),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_607),
.B(n_524),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_608),
.B(n_524),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_L g808 ( 
.A(n_642),
.B(n_196),
.Y(n_808)
);

NAND2x1p5_ASAP7_75t_L g809 ( 
.A(n_591),
.B(n_538),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_697),
.B(n_606),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_616),
.B(n_525),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_619),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_589),
.B(n_337),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_625),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_671),
.B(n_674),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_581),
.A2(n_350),
.B1(n_337),
.B2(n_376),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_584),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_671),
.B(n_197),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_697),
.B(n_540),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_627),
.B(n_525),
.Y(n_820)
);

OAI221xp5_ASAP7_75t_L g821 ( 
.A1(n_643),
.A2(n_548),
.B1(n_542),
.B2(n_540),
.C(n_323),
.Y(n_821)
);

NOR2xp67_ASAP7_75t_L g822 ( 
.A(n_554),
.B(n_701),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_628),
.B(n_483),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_674),
.B(n_197),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_675),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_581),
.A2(n_358),
.B1(n_348),
.B2(n_376),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_558),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_606),
.B(n_690),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_634),
.B(n_198),
.Y(n_829)
);

NOR2xp67_ASAP7_75t_SL g830 ( 
.A(n_675),
.B(n_536),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_646),
.A2(n_536),
.B1(n_219),
.B2(n_375),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_581),
.A2(n_350),
.B1(n_348),
.B2(n_363),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_639),
.B(n_483),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_648),
.B(n_483),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_703),
.B(n_483),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_594),
.B(n_676),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_641),
.B(n_198),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_590),
.B(n_202),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_567),
.Y(n_839)
);

BUFx8_ASAP7_75t_L g840 ( 
.A(n_649),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_568),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_690),
.B(n_540),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_651),
.B(n_647),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_676),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_664),
.B(n_641),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_566),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_566),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_569),
.B(n_483),
.Y(n_848)
);

AND2x6_ASAP7_75t_L g849 ( 
.A(n_570),
.B(n_503),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_631),
.B(n_503),
.Y(n_850)
);

OR2x6_ASAP7_75t_L g851 ( 
.A(n_610),
.B(n_536),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_641),
.B(n_202),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_631),
.B(n_204),
.Y(n_853)
);

NOR2xp67_ASAP7_75t_L g854 ( 
.A(n_622),
.B(n_542),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_564),
.B(n_204),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_564),
.B(n_601),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_691),
.B(n_610),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_598),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_572),
.A2(n_358),
.B1(n_362),
.B2(n_363),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_572),
.A2(n_545),
.B(n_548),
.C(n_542),
.Y(n_860)
);

BUFx6f_ASAP7_75t_SL g861 ( 
.A(n_669),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_598),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_599),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_578),
.B(n_503),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_622),
.A2(n_632),
.B1(n_536),
.B2(n_208),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_599),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_632),
.B(n_208),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_571),
.B(n_209),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_571),
.B(n_209),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_571),
.B(n_210),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_604),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_669),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_578),
.B(n_503),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_597),
.B(n_503),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_702),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_597),
.B(n_515),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_741),
.B(n_789),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_753),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_778),
.A2(n_702),
.B(n_545),
.C(n_679),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_733),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_709),
.A2(n_601),
.B(n_695),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_741),
.B(n_642),
.Y(n_882)
);

NOR2x1_ASAP7_75t_L g883 ( 
.A(n_822),
.B(n_750),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_735),
.B(n_601),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_721),
.A2(n_640),
.B(n_611),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_719),
.Y(n_886)
);

INVx11_ASAP7_75t_L g887 ( 
.A(n_840),
.Y(n_887)
);

NOR2x1p5_ASAP7_75t_L g888 ( 
.A(n_754),
.B(n_362),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_800),
.B(n_642),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_769),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_763),
.B(n_642),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_752),
.B(n_629),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_733),
.B(n_601),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_710),
.B(n_548),
.Y(n_894)
);

BUFx8_ASAP7_75t_L g895 ( 
.A(n_861),
.Y(n_895)
);

AOI21x1_ASAP7_75t_L g896 ( 
.A1(n_760),
.A2(n_624),
.B(n_604),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_760),
.A2(n_640),
.B(n_613),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_706),
.A2(n_638),
.B(n_613),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_787),
.A2(n_368),
.B1(n_361),
.B2(n_284),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_810),
.B(n_248),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_709),
.A2(n_635),
.B(n_695),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_815),
.A2(n_642),
.B1(n_689),
.B2(n_637),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_803),
.B(n_793),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_797),
.Y(n_904)
);

NOR3xp33_ASAP7_75t_L g905 ( 
.A(n_798),
.B(n_349),
.C(n_227),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_711),
.A2(n_635),
.B(n_695),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_819),
.B(n_764),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_753),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_720),
.B(n_642),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_759),
.B(n_637),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_770),
.B(n_652),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_711),
.A2(n_713),
.B(n_762),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_720),
.B(n_689),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_828),
.B(n_767),
.Y(n_914)
);

OAI21xp33_ASAP7_75t_L g915 ( 
.A1(n_793),
.A2(n_787),
.B(n_816),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_725),
.B(n_689),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_799),
.A2(n_601),
.B(n_695),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_725),
.B(n_689),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_797),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_736),
.A2(n_635),
.B(n_695),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_727),
.B(n_689),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_727),
.B(n_689),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_845),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_853),
.B(n_708),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_842),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_853),
.B(n_637),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_736),
.A2(n_612),
.B(n_680),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_SL g928 ( 
.A(n_743),
.B(n_652),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_712),
.B(n_656),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_744),
.B(n_612),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_850),
.A2(n_612),
.B(n_680),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_775),
.A2(n_656),
.B(n_678),
.C(n_620),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_707),
.A2(n_360),
.B1(n_345),
.B2(n_349),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_784),
.A2(n_612),
.B(n_680),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_802),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_784),
.A2(n_612),
.B(n_680),
.Y(n_936)
);

NOR2x1_ASAP7_75t_L g937 ( 
.A(n_803),
.B(n_656),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_804),
.B(n_249),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_817),
.B(n_260),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_761),
.A2(n_615),
.B(n_680),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_715),
.B(n_678),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_755),
.A2(n_224),
.B1(n_227),
.B2(n_226),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_716),
.B(n_678),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_802),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_731),
.A2(n_615),
.B(n_635),
.Y(n_945)
);

NOR3xp33_ASAP7_75t_L g946 ( 
.A(n_775),
.B(n_843),
.C(n_857),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_773),
.A2(n_624),
.B(n_673),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_867),
.A2(n_611),
.B(n_673),
.C(n_662),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_790),
.B(n_262),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_867),
.A2(n_620),
.B(n_662),
.C(n_659),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_732),
.A2(n_615),
.B(n_635),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_773),
.A2(n_615),
.B(n_609),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_739),
.A2(n_615),
.B(n_609),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_815),
.A2(n_609),
.B(n_659),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_734),
.A2(n_609),
.B(n_653),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_747),
.A2(n_609),
.B(n_645),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_842),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_717),
.B(n_621),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_744),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_723),
.B(n_638),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_744),
.B(n_210),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_745),
.B(n_645),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_751),
.A2(n_856),
.B(n_836),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_742),
.A2(n_700),
.B(n_515),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_856),
.A2(n_479),
.B(n_515),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_749),
.B(n_515),
.Y(n_966)
);

NOR3xp33_ASAP7_75t_L g967 ( 
.A(n_837),
.B(n_369),
.C(n_284),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_840),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_744),
.Y(n_969)
);

INVxp67_ASAP7_75t_L g970 ( 
.A(n_813),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_781),
.B(n_263),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_755),
.A2(n_730),
.B1(n_742),
.B2(n_875),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_838),
.A2(n_479),
.B(n_700),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_771),
.A2(n_212),
.B(n_213),
.C(n_217),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_730),
.B(n_212),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_777),
.A2(n_213),
.B(n_217),
.C(n_219),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_722),
.A2(n_345),
.B1(n_224),
.B2(n_226),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_779),
.A2(n_351),
.B(n_344),
.C(n_222),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_805),
.B(n_515),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_772),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_740),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_757),
.A2(n_474),
.B(n_522),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_805),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_SL g984 ( 
.A(n_765),
.B(n_222),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_844),
.B(n_794),
.Y(n_985)
);

AO21x1_ASAP7_75t_L g986 ( 
.A1(n_838),
.A2(n_700),
.B(n_20),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_757),
.A2(n_474),
.B(n_522),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_714),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_855),
.A2(n_351),
.B(n_344),
.C(n_356),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_812),
.B(n_356),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_814),
.B(n_360),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_839),
.B(n_361),
.Y(n_992)
);

AOI21x1_ASAP7_75t_L g993 ( 
.A1(n_766),
.A2(n_700),
.B(n_522),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_714),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_818),
.A2(n_824),
.B(n_852),
.C(n_837),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_848),
.A2(n_700),
.B(n_367),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_852),
.B(n_372),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_841),
.B(n_726),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_718),
.A2(n_368),
.B1(n_369),
.B2(n_367),
.Y(n_999)
);

BUFx8_ASAP7_75t_L g1000 ( 
.A(n_861),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_726),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_825),
.A2(n_375),
.B1(n_266),
.B2(n_324),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_825),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_729),
.B(n_700),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_737),
.A2(n_522),
.B(n_521),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_782),
.B(n_522),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_729),
.B(n_522),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_823),
.A2(n_326),
.B(n_273),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_SL g1009 ( 
.A1(n_864),
.A2(n_19),
.B(n_21),
.C(n_22),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_746),
.B(n_522),
.Y(n_1010)
);

AOI21x1_ASAP7_75t_L g1011 ( 
.A1(n_768),
.A2(n_522),
.B(n_521),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_809),
.A2(n_521),
.B(n_513),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_809),
.A2(n_328),
.B1(n_289),
.B2(n_294),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_746),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_818),
.B(n_272),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_833),
.A2(n_298),
.B(n_312),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_834),
.A2(n_521),
.B(n_513),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_748),
.B(n_521),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_728),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_748),
.B(n_521),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_756),
.B(n_521),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_824),
.B(n_313),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_756),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_738),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_835),
.A2(n_521),
.B(n_513),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_873),
.A2(n_513),
.B(n_507),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_874),
.A2(n_513),
.B(n_507),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_851),
.A2(n_335),
.B1(n_322),
.B2(n_372),
.Y(n_1028)
);

BUFx4f_ASAP7_75t_L g1029 ( 
.A(n_738),
.Y(n_1029)
);

BUFx12f_ASAP7_75t_L g1030 ( 
.A(n_774),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_829),
.B(n_513),
.Y(n_1031)
);

OR2x2_ASAP7_75t_L g1032 ( 
.A(n_816),
.B(n_22),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_776),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_776),
.B(n_513),
.Y(n_1034)
);

OR2x6_ASAP7_75t_L g1035 ( 
.A(n_872),
.B(n_513),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_829),
.B(n_786),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_855),
.A2(n_507),
.B(n_497),
.C(n_474),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_724),
.B(n_183),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_785),
.B(n_507),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_724),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_851),
.B(n_182),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_868),
.A2(n_507),
.B(n_497),
.C(n_28),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_785),
.B(n_507),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_792),
.B(n_507),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_792),
.B(n_507),
.Y(n_1045)
);

OAI321xp33_ASAP7_75t_L g1046 ( 
.A1(n_826),
.A2(n_23),
.A3(n_24),
.B1(n_32),
.B2(n_33),
.C(n_34),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_796),
.A2(n_497),
.B(n_66),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_796),
.B(n_788),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_791),
.B(n_497),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_868),
.A2(n_497),
.B(n_35),
.C(n_37),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_846),
.A2(n_497),
.B(n_76),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_876),
.A2(n_497),
.B(n_177),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_801),
.B(n_497),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_806),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_831),
.B(n_166),
.Y(n_1055)
);

NOR2xp67_ASAP7_75t_L g1056 ( 
.A(n_821),
.B(n_163),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_871),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_807),
.B(n_23),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_811),
.B(n_35),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_820),
.B(n_870),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_826),
.B(n_151),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_780),
.B(n_38),
.Y(n_1062)
);

NAND2x1p5_ASAP7_75t_L g1063 ( 
.A(n_830),
.B(n_148),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_851),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_L g1065 ( 
.A(n_832),
.B(n_40),
.C(n_43),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_969),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1036),
.B(n_832),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_903),
.B(n_795),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_912),
.A2(n_808),
.B(n_783),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_890),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_915),
.A2(n_870),
.B(n_869),
.C(n_854),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1036),
.B(n_877),
.Y(n_1072)
);

INVx4_ASAP7_75t_L g1073 ( 
.A(n_969),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_903),
.B(n_869),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_907),
.A2(n_860),
.B(n_847),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_895),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_R g1077 ( 
.A(n_981),
.B(n_871),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1032),
.A2(n_924),
.B1(n_972),
.B2(n_1065),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_887),
.Y(n_1079)
);

BUFx4f_ASAP7_75t_L g1080 ( 
.A(n_1064),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_995),
.A2(n_859),
.B(n_865),
.C(n_866),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_926),
.A2(n_863),
.B(n_862),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1054),
.B(n_859),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_1015),
.A2(n_858),
.B(n_862),
.C(n_863),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_1015),
.A2(n_847),
.B(n_827),
.C(n_758),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_904),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1054),
.B(n_849),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_919),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1060),
.A2(n_1061),
.B1(n_1041),
.B2(n_923),
.Y(n_1089)
);

NOR3xp33_ASAP7_75t_SL g1090 ( 
.A(n_1046),
.B(n_40),
.C(n_44),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1041),
.A2(n_849),
.B1(n_47),
.B2(n_48),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_946),
.B(n_849),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_894),
.B(n_849),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_886),
.B(n_849),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_923),
.B(n_44),
.Y(n_1095)
);

OA22x2_ASAP7_75t_L g1096 ( 
.A1(n_970),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_963),
.A2(n_138),
.B(n_118),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_900),
.B(n_50),
.Y(n_1098)
);

INVx2_ASAP7_75t_SL g1099 ( 
.A(n_890),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_914),
.B(n_51),
.Y(n_1100)
);

INVx4_ASAP7_75t_L g1101 ( 
.A(n_969),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_946),
.B(n_113),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_980),
.B(n_52),
.Y(n_1103)
);

INVxp67_ASAP7_75t_L g1104 ( 
.A(n_911),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_940),
.A2(n_889),
.B(n_1048),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_970),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_895),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_1022),
.A2(n_52),
.B(n_53),
.C(n_55),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_900),
.B(n_1033),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1033),
.Y(n_1110)
);

NOR2xp67_ASAP7_75t_SL g1111 ( 
.A(n_1064),
.B(n_55),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_1064),
.B(n_77),
.Y(n_1112)
);

INVxp67_ASAP7_75t_L g1113 ( 
.A(n_938),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_997),
.B(n_58),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1064),
.B(n_84),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1022),
.B(n_58),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_883),
.B(n_86),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_949),
.B(n_60),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_1000),
.Y(n_1119)
);

AND2x6_ASAP7_75t_L g1120 ( 
.A(n_1038),
.B(n_91),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_985),
.B(n_106),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_989),
.A2(n_60),
.B(n_63),
.C(n_65),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_967),
.A2(n_65),
.B1(n_908),
.B2(n_878),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_967),
.A2(n_925),
.B1(n_957),
.B2(n_1062),
.Y(n_1124)
);

AND2x2_ASAP7_75t_SL g1125 ( 
.A(n_1029),
.B(n_928),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_SL g1126 ( 
.A1(n_1019),
.A2(n_1030),
.B1(n_1024),
.B2(n_949),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_SL g1127 ( 
.A1(n_1062),
.A2(n_1047),
.B(n_1051),
.C(n_971),
.Y(n_1127)
);

O2A1O1Ixp5_ASAP7_75t_L g1128 ( 
.A1(n_882),
.A2(n_973),
.B(n_1006),
.C(n_884),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_983),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_920),
.A2(n_927),
.B(n_896),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_1000),
.Y(n_1131)
);

INVx5_ASAP7_75t_L g1132 ( 
.A(n_969),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1055),
.A2(n_1056),
.B1(n_975),
.B2(n_905),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1006),
.A2(n_885),
.B(n_917),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_931),
.A2(n_898),
.B(n_953),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_938),
.B(n_939),
.Y(n_1136)
);

AOI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_930),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_893),
.A2(n_930),
.B(n_945),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1038),
.B(n_1003),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_971),
.A2(n_1059),
.B(n_1058),
.C(n_891),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1008),
.A2(n_1016),
.B(n_939),
.C(n_976),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_888),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_974),
.A2(n_978),
.B(n_999),
.C(n_879),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1050),
.A2(n_944),
.B1(n_935),
.B2(n_1042),
.Y(n_1144)
);

AND2x4_ASAP7_75t_SL g1145 ( 
.A(n_880),
.B(n_959),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1023),
.B(n_988),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_1040),
.B(n_880),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_893),
.A2(n_951),
.B(n_921),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_998),
.Y(n_1149)
);

XOR2x2_ASAP7_75t_L g1150 ( 
.A(n_905),
.B(n_899),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_959),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_910),
.B(n_1003),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_990),
.B(n_991),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_909),
.A2(n_916),
.B(n_918),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_994),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_977),
.A2(n_1029),
.B1(n_964),
.B2(n_922),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_910),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1028),
.B(n_984),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_932),
.A2(n_948),
.B(n_950),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_992),
.B(n_937),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1001),
.B(n_1014),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_SL g1162 ( 
.A(n_968),
.B(n_1063),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_958),
.Y(n_1163)
);

CKINVDCx16_ASAP7_75t_R g1164 ( 
.A(n_1035),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_913),
.A2(n_1049),
.B(n_936),
.Y(n_1165)
);

OAI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1035),
.A2(n_942),
.B1(n_1013),
.B2(n_1002),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_961),
.A2(n_965),
.B(n_996),
.C(n_962),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1057),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_933),
.A2(n_1009),
.B(n_960),
.C(n_1037),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1057),
.B(n_943),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_966),
.A2(n_929),
.B(n_941),
.C(n_892),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_L g1172 ( 
.A(n_1035),
.B(n_902),
.C(n_1052),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_979),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1034),
.B(n_1044),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1063),
.Y(n_1175)
);

OAI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1004),
.A2(n_1007),
.B1(n_1018),
.B2(n_1045),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_897),
.A2(n_881),
.B1(n_901),
.B2(n_906),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1010),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_947),
.A2(n_934),
.B(n_1027),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1020),
.A2(n_1043),
.B1(n_1039),
.B2(n_1021),
.Y(n_1180)
);

CKINVDCx8_ASAP7_75t_R g1181 ( 
.A(n_986),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_952),
.A2(n_955),
.B(n_956),
.Y(n_1182)
);

NAND3xp33_ASAP7_75t_SL g1183 ( 
.A(n_1053),
.B(n_954),
.C(n_982),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_1044),
.B(n_1034),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1026),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_993),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1012),
.A2(n_987),
.B1(n_1017),
.B2(n_1025),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1005),
.A2(n_583),
.B(n_580),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_915),
.A2(n_903),
.B(n_995),
.C(n_1036),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_903),
.A2(n_915),
.B(n_752),
.C(n_778),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_903),
.B(n_752),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1064),
.Y(n_1192)
);

OR2x6_ASAP7_75t_L g1193 ( 
.A(n_1064),
.B(n_1041),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_904),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_904),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_903),
.A2(n_915),
.B1(n_787),
.B2(n_755),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_903),
.B(n_752),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1036),
.B(n_877),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_903),
.A2(n_915),
.B(n_752),
.C(n_778),
.Y(n_1199)
);

O2A1O1Ixp5_ASAP7_75t_L g1200 ( 
.A1(n_903),
.A2(n_709),
.B(n_711),
.C(n_1036),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_SL g1201 ( 
.A1(n_903),
.A2(n_582),
.B(n_623),
.C(n_614),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1064),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_SL g1203 ( 
.A(n_915),
.B(n_903),
.Y(n_1203)
);

O2A1O1Ixp5_ASAP7_75t_SL g1204 ( 
.A1(n_884),
.A2(n_838),
.B(n_1061),
.C(n_975),
.Y(n_1204)
);

BUFx8_ASAP7_75t_SL g1205 ( 
.A(n_981),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_895),
.Y(n_1206)
);

BUFx12f_ASAP7_75t_L g1207 ( 
.A(n_895),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_911),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_SL g1209 ( 
.A1(n_1061),
.A2(n_711),
.B(n_709),
.C(n_1050),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_911),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1036),
.B(n_877),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_912),
.A2(n_583),
.B(n_580),
.Y(n_1212)
);

INVx4_ASAP7_75t_L g1213 ( 
.A(n_969),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_904),
.Y(n_1214)
);

AOI21x1_ASAP7_75t_L g1215 ( 
.A1(n_884),
.A2(n_736),
.B(n_711),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1036),
.B(n_877),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1036),
.B(n_877),
.Y(n_1217)
);

NOR3xp33_ASAP7_75t_SL g1218 ( 
.A(n_915),
.B(n_704),
.C(n_490),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_903),
.A2(n_915),
.B1(n_787),
.B2(n_755),
.Y(n_1219)
);

NAND2xp33_ASAP7_75t_L g1220 ( 
.A(n_1064),
.B(n_915),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_903),
.B(n_735),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_912),
.A2(n_583),
.B(n_580),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_904),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1212),
.A2(n_1222),
.B(n_1188),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1134),
.A2(n_1069),
.B(n_1135),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1118),
.A2(n_1199),
.B(n_1190),
.C(n_1141),
.Y(n_1226)
);

OAI22x1_ASAP7_75t_L g1227 ( 
.A1(n_1191),
.A2(n_1197),
.B1(n_1103),
.B2(n_1221),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1130),
.A2(n_1148),
.B(n_1138),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1200),
.A2(n_1128),
.B(n_1196),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1105),
.A2(n_1071),
.B(n_1167),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1136),
.A2(n_1203),
.B1(n_1150),
.B2(n_1158),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1127),
.A2(n_1140),
.B(n_1075),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1070),
.Y(n_1233)
);

AO32x2_ASAP7_75t_L g1234 ( 
.A1(n_1196),
.A2(n_1219),
.A3(n_1078),
.B1(n_1144),
.B2(n_1089),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1129),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1072),
.B(n_1198),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1146),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1113),
.B(n_1125),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1074),
.A2(n_1179),
.B(n_1165),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1082),
.A2(n_1182),
.B(n_1154),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1201),
.A2(n_1116),
.B(n_1219),
.C(n_1203),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1179),
.A2(n_1177),
.B(n_1211),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1216),
.B(n_1217),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1153),
.A2(n_1067),
.B(n_1098),
.C(n_1143),
.Y(n_1244)
);

OA21x2_ASAP7_75t_L g1245 ( 
.A1(n_1159),
.A2(n_1084),
.B(n_1172),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1193),
.B(n_1147),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1104),
.A2(n_1068),
.B1(n_1210),
.B2(n_1208),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_1159),
.A2(n_1185),
.B(n_1085),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1086),
.Y(n_1249)
);

BUFx10_ASAP7_75t_L g1250 ( 
.A(n_1100),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1187),
.A2(n_1137),
.B(n_1180),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1204),
.A2(n_1078),
.B(n_1169),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1144),
.A2(n_1180),
.A3(n_1156),
.B(n_1089),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1218),
.B(n_1109),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1156),
.A2(n_1184),
.A3(n_1186),
.B(n_1121),
.Y(n_1255)
);

NAND3xp33_ASAP7_75t_L g1256 ( 
.A(n_1133),
.B(n_1123),
.C(n_1124),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1097),
.A2(n_1170),
.B(n_1183),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1149),
.B(n_1083),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_1121),
.A2(n_1108),
.A3(n_1091),
.B(n_1178),
.Y(n_1259)
);

NOR4xp25_ASAP7_75t_L g1260 ( 
.A(n_1122),
.B(n_1166),
.C(n_1081),
.D(n_1091),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_SL g1261 ( 
.A1(n_1093),
.A2(n_1175),
.B(n_1102),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1193),
.B(n_1147),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1092),
.A2(n_1209),
.B(n_1220),
.Y(n_1263)
);

OAI21xp33_ASAP7_75t_L g1264 ( 
.A1(n_1090),
.A2(n_1114),
.B(n_1095),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1193),
.B(n_1202),
.Y(n_1265)
);

BUFx8_ASAP7_75t_L g1266 ( 
.A(n_1207),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1181),
.A2(n_1163),
.B1(n_1096),
.B2(n_1164),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1171),
.A2(n_1146),
.B(n_1161),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1173),
.B(n_1094),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1176),
.A2(n_1139),
.B(n_1160),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1087),
.A2(n_1152),
.B(n_1132),
.Y(n_1271)
);

AO31x2_ASAP7_75t_L g1272 ( 
.A1(n_1155),
.A2(n_1223),
.A3(n_1214),
.B(n_1195),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1088),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1157),
.B(n_1099),
.Y(n_1274)
);

AO31x2_ASAP7_75t_L g1275 ( 
.A1(n_1194),
.A2(n_1168),
.A3(n_1073),
.B(n_1066),
.Y(n_1275)
);

BUFx12f_ASAP7_75t_L g1276 ( 
.A(n_1107),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1106),
.B(n_1157),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1066),
.A2(n_1073),
.A3(n_1213),
.B(n_1101),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1157),
.B(n_1120),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1174),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1077),
.Y(n_1281)
);

INVx5_ASAP7_75t_L g1282 ( 
.A(n_1205),
.Y(n_1282)
);

NAND3xp33_ASAP7_75t_L g1283 ( 
.A(n_1111),
.B(n_1162),
.C(n_1115),
.Y(n_1283)
);

BUFx2_ASAP7_75t_SL g1284 ( 
.A(n_1192),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1151),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1151),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1192),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1132),
.A2(n_1162),
.B(n_1117),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1096),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1132),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1132),
.A2(n_1175),
.B(n_1080),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1175),
.A2(n_1112),
.B(n_1213),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_SL g1293 ( 
.A1(n_1101),
.A2(n_1202),
.B(n_1192),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1202),
.A2(n_1126),
.B1(n_1142),
.B2(n_1145),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_SL g1295 ( 
.A1(n_1120),
.A2(n_1076),
.B(n_1119),
.C(n_1131),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1120),
.A2(n_1079),
.B(n_1206),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1120),
.B(n_1072),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1212),
.A2(n_583),
.B(n_580),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1072),
.B(n_1198),
.Y(n_1299)
);

CKINVDCx11_ASAP7_75t_R g1300 ( 
.A(n_1207),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1110),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1130),
.A2(n_1148),
.B(n_1138),
.Y(n_1302)
);

AOI221xp5_ASAP7_75t_L g1303 ( 
.A1(n_1196),
.A2(n_915),
.B1(n_1219),
.B2(n_903),
.C(n_1118),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1189),
.A2(n_1200),
.B(n_1128),
.Y(n_1304)
);

NAND3xp33_ASAP7_75t_L g1305 ( 
.A(n_1201),
.B(n_1118),
.C(n_903),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1212),
.A2(n_583),
.B(n_580),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1151),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1212),
.A2(n_583),
.B(n_580),
.Y(n_1308)
);

OAI211xp5_ASAP7_75t_SL g1309 ( 
.A1(n_1218),
.A2(n_752),
.B(n_1113),
.C(n_915),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1212),
.A2(n_583),
.B(n_580),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1118),
.A2(n_903),
.B(n_1199),
.C(n_1190),
.Y(n_1311)
);

NOR2xp67_ASAP7_75t_L g1312 ( 
.A(n_1104),
.B(n_804),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1136),
.B(n_710),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1110),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1070),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1136),
.B(n_710),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1212),
.A2(n_583),
.B(n_580),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1212),
.A2(n_583),
.B(n_580),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1136),
.B(n_710),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1072),
.B(n_1198),
.Y(n_1320)
);

INVx5_ASAP7_75t_L g1321 ( 
.A(n_1205),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1130),
.A2(n_1148),
.B(n_1138),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1212),
.A2(n_583),
.B(n_580),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1151),
.Y(n_1324)
);

OAI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1067),
.A2(n_928),
.B1(n_752),
.B2(n_743),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_1106),
.Y(n_1326)
);

AO32x2_ASAP7_75t_L g1327 ( 
.A1(n_1196),
.A2(n_1219),
.A3(n_1078),
.B1(n_1144),
.B2(n_1089),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1118),
.A2(n_915),
.B1(n_903),
.B2(n_1150),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1128),
.A2(n_1159),
.B(n_1134),
.Y(n_1329)
);

O2A1O1Ixp5_ASAP7_75t_L g1330 ( 
.A1(n_1201),
.A2(n_1118),
.B(n_903),
.C(n_1068),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1110),
.Y(n_1331)
);

AOI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1212),
.A2(n_1222),
.B(n_1215),
.Y(n_1332)
);

O2A1O1Ixp33_ASAP7_75t_SL g1333 ( 
.A1(n_1201),
.A2(n_1141),
.B(n_1189),
.C(n_1127),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1130),
.A2(n_1148),
.B(n_1138),
.Y(n_1334)
);

AOI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1212),
.A2(n_1222),
.B(n_1215),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1212),
.A2(n_583),
.B(n_580),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1130),
.A2(n_1148),
.B(n_1138),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1072),
.B(n_1198),
.Y(n_1338)
);

OAI22x1_ASAP7_75t_L g1339 ( 
.A1(n_1118),
.A2(n_903),
.B1(n_1197),
.B2(n_1191),
.Y(n_1339)
);

AOI221x1_ASAP7_75t_L g1340 ( 
.A1(n_1196),
.A2(n_1219),
.B1(n_1189),
.B2(n_915),
.C(n_1118),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1118),
.A2(n_903),
.B(n_1199),
.C(n_1190),
.Y(n_1341)
);

NAND2xp33_ASAP7_75t_L g1342 ( 
.A(n_1189),
.B(n_1064),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1136),
.B(n_710),
.Y(n_1343)
);

INVx2_ASAP7_75t_SL g1344 ( 
.A(n_1070),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1118),
.A2(n_903),
.B(n_1199),
.C(n_1190),
.Y(n_1345)
);

AO21x2_ASAP7_75t_L g1346 ( 
.A1(n_1159),
.A2(n_1135),
.B(n_1179),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1208),
.B(n_980),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1072),
.B(n_1198),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1208),
.Y(n_1349)
);

O2A1O1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1201),
.A2(n_1118),
.B(n_903),
.C(n_1221),
.Y(n_1350)
);

NOR2xp67_ASAP7_75t_L g1351 ( 
.A(n_1104),
.B(n_804),
.Y(n_1351)
);

O2A1O1Ixp33_ASAP7_75t_SL g1352 ( 
.A1(n_1201),
.A2(n_1141),
.B(n_1189),
.C(n_1127),
.Y(n_1352)
);

AOI211x1_ASAP7_75t_L g1353 ( 
.A1(n_1067),
.A2(n_915),
.B(n_1219),
.C(n_1196),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1208),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_SL g1355 ( 
.A1(n_1136),
.A2(n_915),
.B(n_1118),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1189),
.A2(n_1200),
.B(n_1128),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1130),
.A2(n_1148),
.B(n_1138),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1189),
.A2(n_1200),
.B(n_1128),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1212),
.A2(n_583),
.B(n_580),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1110),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1136),
.B(n_710),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1189),
.A2(n_1200),
.B(n_1128),
.Y(n_1362)
);

AOI221x1_ASAP7_75t_L g1363 ( 
.A1(n_1196),
.A2(n_1219),
.B1(n_1189),
.B2(n_915),
.C(n_1118),
.Y(n_1363)
);

CKINVDCx6p67_ASAP7_75t_R g1364 ( 
.A(n_1207),
.Y(n_1364)
);

O2A1O1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1201),
.A2(n_1118),
.B(n_903),
.C(n_1221),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1128),
.A2(n_1159),
.B(n_1134),
.Y(n_1366)
);

INVx4_ASAP7_75t_L g1367 ( 
.A(n_1132),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1072),
.B(n_1198),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1212),
.A2(n_583),
.B(n_580),
.Y(n_1369)
);

AOI221x1_ASAP7_75t_L g1370 ( 
.A1(n_1196),
.A2(n_1219),
.B1(n_1189),
.B2(n_915),
.C(n_1118),
.Y(n_1370)
);

AOI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1212),
.A2(n_1222),
.B(n_1215),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1118),
.A2(n_903),
.B1(n_772),
.B2(n_582),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1212),
.A2(n_583),
.B(n_580),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1212),
.A2(n_583),
.B(n_580),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1072),
.B(n_1198),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1070),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1212),
.A2(n_583),
.B(n_580),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1072),
.B(n_1198),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1212),
.A2(n_583),
.B(n_580),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1282),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_SL g1381 ( 
.A1(n_1256),
.A2(n_1267),
.B1(n_1342),
.B2(n_1305),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1328),
.A2(n_1372),
.B1(n_1256),
.B2(n_1303),
.Y(n_1382)
);

INVx6_ASAP7_75t_L g1383 ( 
.A(n_1246),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1243),
.B(n_1236),
.Y(n_1384)
);

INVx4_ASAP7_75t_L g1385 ( 
.A(n_1367),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1367),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1231),
.A2(n_1305),
.B1(n_1339),
.B2(n_1227),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_SL g1388 ( 
.A1(n_1281),
.A2(n_1282),
.B1(n_1321),
.B2(n_1283),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1249),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1325),
.A2(n_1254),
.B1(n_1309),
.B2(n_1264),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1354),
.Y(n_1391)
);

INVx6_ASAP7_75t_L g1392 ( 
.A(n_1262),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1264),
.A2(n_1267),
.B1(n_1320),
.B2(n_1338),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_1300),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1348),
.A2(n_1368),
.B1(n_1375),
.B2(n_1299),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_1349),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1349),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1225),
.A2(n_1230),
.B(n_1239),
.Y(n_1398)
);

OAI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1355),
.A2(n_1236),
.B1(n_1378),
.B2(n_1299),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1238),
.A2(n_1316),
.B1(n_1343),
.B2(n_1361),
.Y(n_1400)
);

INVx4_ASAP7_75t_L g1401 ( 
.A(n_1321),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1355),
.A2(n_1319),
.B1(n_1313),
.B2(n_1283),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1321),
.Y(n_1403)
);

BUFx2_ASAP7_75t_SL g1404 ( 
.A(n_1312),
.Y(n_1404)
);

CKINVDCx11_ASAP7_75t_R g1405 ( 
.A(n_1364),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1331),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1297),
.A2(n_1347),
.B1(n_1250),
.B2(n_1346),
.Y(n_1407)
);

BUFx8_ASAP7_75t_L g1408 ( 
.A(n_1277),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1360),
.Y(n_1409)
);

INVx6_ASAP7_75t_L g1410 ( 
.A(n_1262),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1378),
.B(n_1311),
.Y(n_1411)
);

CKINVDCx11_ASAP7_75t_R g1412 ( 
.A(n_1281),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1250),
.A2(n_1346),
.B1(n_1289),
.B2(n_1263),
.Y(n_1413)
);

INVx8_ASAP7_75t_L g1414 ( 
.A(n_1265),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_1266),
.Y(n_1415)
);

BUFx12f_ASAP7_75t_L g1416 ( 
.A(n_1266),
.Y(n_1416)
);

OAI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1340),
.A2(n_1370),
.B1(n_1363),
.B2(n_1258),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1233),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1296),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1301),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1341),
.A2(n_1345),
.B1(n_1226),
.B2(n_1244),
.Y(n_1421)
);

INVx6_ASAP7_75t_L g1422 ( 
.A(n_1284),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1263),
.A2(n_1269),
.B1(n_1280),
.B2(n_1247),
.Y(n_1423)
);

CKINVDCx11_ASAP7_75t_R g1424 ( 
.A(n_1314),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1273),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1350),
.A2(n_1365),
.B(n_1241),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1248),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1272),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1344),
.Y(n_1429)
);

OAI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1237),
.A2(n_1252),
.B1(n_1304),
.B2(n_1362),
.Y(n_1430)
);

CKINVDCx11_ASAP7_75t_R g1431 ( 
.A(n_1287),
.Y(n_1431)
);

AOI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1351),
.A2(n_1294),
.B1(n_1279),
.B2(n_1295),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1252),
.A2(n_1356),
.B1(n_1358),
.B2(n_1362),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1304),
.A2(n_1356),
.B1(n_1358),
.B2(n_1229),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1229),
.A2(n_1242),
.B1(n_1245),
.B2(n_1232),
.Y(n_1435)
);

BUFx4f_ASAP7_75t_SL g1436 ( 
.A(n_1287),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1275),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1315),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1270),
.A2(n_1245),
.B1(n_1376),
.B2(n_1326),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1329),
.A2(n_1366),
.B1(n_1248),
.B2(n_1260),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1329),
.A2(n_1366),
.B1(n_1260),
.B2(n_1294),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1353),
.A2(n_1327),
.B1(n_1234),
.B2(n_1274),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_SL g1443 ( 
.A1(n_1234),
.A2(n_1327),
.B1(n_1288),
.B2(n_1253),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_1285),
.Y(n_1444)
);

OAI21xp33_ASAP7_75t_L g1445 ( 
.A1(n_1261),
.A2(n_1292),
.B(n_1268),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1286),
.Y(n_1446)
);

BUFx12f_ASAP7_75t_L g1447 ( 
.A(n_1293),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1307),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1290),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1324),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1234),
.A2(n_1327),
.B1(n_1291),
.B2(n_1271),
.Y(n_1451)
);

BUFx4_ASAP7_75t_SL g1452 ( 
.A(n_1330),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_1251),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1224),
.A2(n_1257),
.B1(n_1377),
.B2(n_1374),
.Y(n_1454)
);

OAI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1333),
.A2(n_1352),
.B1(n_1373),
.B2(n_1369),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1259),
.B(n_1253),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1298),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1278),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1259),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1306),
.A2(n_1379),
.B1(n_1359),
.B2(n_1336),
.Y(n_1460)
);

BUFx12f_ASAP7_75t_L g1461 ( 
.A(n_1259),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1308),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1310),
.A2(n_1323),
.B1(n_1318),
.B2(n_1317),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1228),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1240),
.A2(n_1334),
.B1(n_1357),
.B2(n_1302),
.Y(n_1465)
);

NAND2xp33_ASAP7_75t_SL g1466 ( 
.A(n_1253),
.B(n_1255),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_SL g1467 ( 
.A1(n_1322),
.A2(n_1337),
.B1(n_1255),
.B2(n_1335),
.Y(n_1467)
);

OAI21xp33_ASAP7_75t_L g1468 ( 
.A1(n_1332),
.A2(n_1371),
.B(n_1255),
.Y(n_1468)
);

CKINVDCx11_ASAP7_75t_R g1469 ( 
.A(n_1300),
.Y(n_1469)
);

CKINVDCx11_ASAP7_75t_R g1470 ( 
.A(n_1300),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_1233),
.Y(n_1471)
);

BUFx8_ASAP7_75t_L g1472 ( 
.A(n_1276),
.Y(n_1472)
);

OAI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1372),
.A2(n_1231),
.B1(n_1067),
.B2(n_1203),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1249),
.Y(n_1474)
);

BUFx8_ASAP7_75t_L g1475 ( 
.A(n_1276),
.Y(n_1475)
);

INVx6_ASAP7_75t_L g1476 ( 
.A(n_1246),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1349),
.Y(n_1477)
);

BUFx10_ASAP7_75t_L g1478 ( 
.A(n_1344),
.Y(n_1478)
);

CKINVDCx20_ASAP7_75t_R g1479 ( 
.A(n_1300),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1235),
.Y(n_1480)
);

BUFx4_ASAP7_75t_SL g1481 ( 
.A(n_1347),
.Y(n_1481)
);

CKINVDCx6p67_ASAP7_75t_R g1482 ( 
.A(n_1282),
.Y(n_1482)
);

BUFx10_ASAP7_75t_L g1483 ( 
.A(n_1344),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1354),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1313),
.B(n_1316),
.Y(n_1485)
);

BUFx2_ASAP7_75t_SL g1486 ( 
.A(n_1282),
.Y(n_1486)
);

CKINVDCx20_ASAP7_75t_R g1487 ( 
.A(n_1300),
.Y(n_1487)
);

CKINVDCx11_ASAP7_75t_R g1488 ( 
.A(n_1300),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1235),
.Y(n_1489)
);

INVx3_ASAP7_75t_SL g1490 ( 
.A(n_1282),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1347),
.B(n_1349),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1347),
.B(n_1349),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1328),
.A2(n_1150),
.B1(n_915),
.B2(n_1372),
.Y(n_1493)
);

INVx6_ASAP7_75t_L g1494 ( 
.A(n_1246),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1235),
.Y(n_1495)
);

INVx4_ASAP7_75t_L g1496 ( 
.A(n_1367),
.Y(n_1496)
);

CKINVDCx11_ASAP7_75t_R g1497 ( 
.A(n_1300),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1328),
.A2(n_1150),
.B1(n_915),
.B2(n_1372),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1265),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1354),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1328),
.A2(n_1150),
.B1(n_915),
.B2(n_1372),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1243),
.B(n_1236),
.Y(n_1502)
);

INVx6_ASAP7_75t_L g1503 ( 
.A(n_1246),
.Y(n_1503)
);

AO21x2_ASAP7_75t_L g1504 ( 
.A1(n_1398),
.A2(n_1434),
.B(n_1455),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1469),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1384),
.B(n_1502),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1493),
.A2(n_1501),
.B(n_1498),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1428),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1419),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1456),
.B(n_1433),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1408),
.Y(n_1511)
);

CKINVDCx20_ASAP7_75t_R g1512 ( 
.A(n_1470),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1437),
.Y(n_1513)
);

OR2x6_ASAP7_75t_L g1514 ( 
.A(n_1426),
.B(n_1461),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1488),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1459),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1433),
.B(n_1443),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1427),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1454),
.A2(n_1463),
.B(n_1460),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1465),
.A2(n_1453),
.B(n_1468),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1458),
.Y(n_1521)
);

OAI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1382),
.A2(n_1421),
.B(n_1473),
.Y(n_1522)
);

AND2x6_ASAP7_75t_L g1523 ( 
.A(n_1419),
.B(n_1432),
.Y(n_1523)
);

AOI222xp33_ASAP7_75t_L g1524 ( 
.A1(n_1473),
.A2(n_1390),
.B1(n_1393),
.B2(n_1387),
.C1(n_1411),
.C2(n_1434),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1381),
.A2(n_1445),
.B(n_1393),
.C(n_1411),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1430),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1430),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1442),
.Y(n_1528)
);

CKINVDCx11_ASAP7_75t_R g1529 ( 
.A(n_1497),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1442),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1381),
.A2(n_1388),
.B1(n_1407),
.B2(n_1402),
.Y(n_1531)
);

NAND2x1p5_ASAP7_75t_L g1532 ( 
.A(n_1419),
.B(n_1464),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1451),
.Y(n_1533)
);

INVx3_ASAP7_75t_L g1534 ( 
.A(n_1462),
.Y(n_1534)
);

AOI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1449),
.A2(n_1495),
.B(n_1480),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1395),
.A2(n_1502),
.B(n_1384),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1466),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1447),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1489),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1443),
.B(n_1441),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1395),
.B(n_1423),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1408),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1491),
.B(n_1492),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1453),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1435),
.A2(n_1440),
.B(n_1441),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1412),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1406),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1409),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1399),
.B(n_1485),
.Y(n_1549)
);

INVx4_ASAP7_75t_SL g1550 ( 
.A(n_1490),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1425),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1420),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_1396),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_1422),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_SL g1555 ( 
.A1(n_1413),
.A2(n_1439),
.B(n_1435),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1422),
.Y(n_1556)
);

OR2x6_ASAP7_75t_L g1557 ( 
.A(n_1486),
.B(n_1401),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1440),
.A2(n_1386),
.B(n_1467),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1457),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1389),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1399),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1474),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1417),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1417),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1455),
.A2(n_1467),
.B(n_1450),
.Y(n_1565)
);

AOI221x1_ASAP7_75t_SL g1566 ( 
.A1(n_1452),
.A2(n_1481),
.B1(n_1400),
.B2(n_1404),
.C(n_1424),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1452),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1405),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1471),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1436),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1471),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1448),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1391),
.A2(n_1484),
.B1(n_1500),
.B2(n_1401),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_SL g1574 ( 
.A1(n_1385),
.A2(n_1496),
.B(n_1418),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1397),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1477),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1436),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1444),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1438),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1429),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1383),
.Y(n_1581)
);

OA21x2_ASAP7_75t_L g1582 ( 
.A1(n_1380),
.A2(n_1403),
.B(n_1481),
.Y(n_1582)
);

AOI21x1_ASAP7_75t_L g1583 ( 
.A1(n_1383),
.A2(n_1503),
.B(n_1392),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1431),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1392),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1499),
.B(n_1503),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1410),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_SL g1588 ( 
.A(n_1416),
.B(n_1394),
.Y(n_1588)
);

OAI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1414),
.A2(n_1494),
.B(n_1476),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1482),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1494),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1446),
.B(n_1414),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1478),
.B(n_1483),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1510),
.B(n_1478),
.Y(n_1594)
);

OAI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1522),
.A2(n_1415),
.B(n_1487),
.Y(n_1595)
);

A2O1A1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1525),
.A2(n_1479),
.B(n_1472),
.C(n_1475),
.Y(n_1596)
);

OAI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1507),
.A2(n_1475),
.B(n_1524),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1541),
.A2(n_1534),
.B1(n_1531),
.B2(n_1559),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1534),
.B(n_1543),
.Y(n_1599)
);

NOR2x1_ASAP7_75t_R g1600 ( 
.A(n_1529),
.B(n_1505),
.Y(n_1600)
);

OR2x6_ASAP7_75t_L g1601 ( 
.A(n_1514),
.B(n_1555),
.Y(n_1601)
);

OA21x2_ASAP7_75t_L g1602 ( 
.A1(n_1520),
.A2(n_1545),
.B(n_1558),
.Y(n_1602)
);

OAI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1519),
.A2(n_1536),
.B(n_1527),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1539),
.Y(n_1604)
);

OAI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1526),
.A2(n_1527),
.B(n_1561),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1518),
.Y(n_1606)
);

CKINVDCx20_ASAP7_75t_R g1607 ( 
.A(n_1512),
.Y(n_1607)
);

O2A1O1Ixp33_ASAP7_75t_L g1608 ( 
.A1(n_1555),
.A2(n_1526),
.B(n_1567),
.C(n_1563),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1506),
.B(n_1549),
.Y(n_1609)
);

OAI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1561),
.A2(n_1567),
.B(n_1563),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_SL g1611 ( 
.A1(n_1517),
.A2(n_1540),
.B1(n_1504),
.B2(n_1523),
.Y(n_1611)
);

NAND3xp33_ASAP7_75t_SL g1612 ( 
.A(n_1588),
.B(n_1546),
.C(n_1515),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1546),
.Y(n_1613)
);

NAND3xp33_ASAP7_75t_L g1614 ( 
.A(n_1564),
.B(n_1573),
.C(n_1572),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1577),
.A2(n_1570),
.B1(n_1580),
.B2(n_1582),
.Y(n_1615)
);

NOR2x1_ASAP7_75t_SL g1616 ( 
.A(n_1583),
.B(n_1504),
.Y(n_1616)
);

NAND2xp33_ASAP7_75t_L g1617 ( 
.A(n_1538),
.B(n_1523),
.Y(n_1617)
);

A2O1A1Ixp33_ASAP7_75t_L g1618 ( 
.A1(n_1517),
.A2(n_1566),
.B(n_1545),
.C(n_1540),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_SL g1619 ( 
.A1(n_1574),
.A2(n_1535),
.B(n_1582),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1557),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1535),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1579),
.B(n_1575),
.Y(n_1622)
);

NAND4xp25_ASAP7_75t_L g1623 ( 
.A(n_1576),
.B(n_1571),
.C(n_1569),
.D(n_1579),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1547),
.B(n_1586),
.Y(n_1624)
);

AO32x2_ASAP7_75t_L g1625 ( 
.A1(n_1554),
.A2(n_1556),
.A3(n_1528),
.B1(n_1530),
.B2(n_1533),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1582),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1553),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1518),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1509),
.B(n_1589),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1548),
.B(n_1551),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1523),
.A2(n_1538),
.B1(n_1578),
.B2(n_1582),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1552),
.B(n_1528),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1565),
.A2(n_1544),
.B(n_1532),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1587),
.B(n_1578),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1560),
.B(n_1562),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1589),
.B(n_1550),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1602),
.B(n_1565),
.Y(n_1637)
);

NAND3xp33_ASAP7_75t_L g1638 ( 
.A(n_1597),
.B(n_1538),
.C(n_1581),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1626),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1625),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1625),
.B(n_1537),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1606),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1633),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1625),
.B(n_1508),
.Y(n_1644)
);

INVx2_ASAP7_75t_SL g1645 ( 
.A(n_1629),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1621),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1611),
.B(n_1516),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1614),
.B(n_1585),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1604),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1616),
.B(n_1513),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1603),
.B(n_1624),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_SL g1652 ( 
.A1(n_1595),
.A2(n_1523),
.B1(n_1617),
.B2(n_1610),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1606),
.B(n_1628),
.Y(n_1653)
);

BUFx2_ASAP7_75t_L g1654 ( 
.A(n_1629),
.Y(n_1654)
);

CKINVDCx20_ASAP7_75t_R g1655 ( 
.A(n_1607),
.Y(n_1655)
);

OR2x2_ASAP7_75t_SL g1656 ( 
.A(n_1612),
.B(n_1591),
.Y(n_1656)
);

NOR2xp67_ASAP7_75t_L g1657 ( 
.A(n_1636),
.B(n_1521),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_L g1658 ( 
.A(n_1636),
.B(n_1521),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_1622),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1632),
.Y(n_1660)
);

NAND4xp25_ASAP7_75t_L g1661 ( 
.A(n_1638),
.B(n_1596),
.C(n_1598),
.D(n_1608),
.Y(n_1661)
);

BUFx3_ASAP7_75t_L g1662 ( 
.A(n_1639),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1640),
.B(n_1623),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1646),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1657),
.B(n_1620),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1654),
.B(n_1645),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1645),
.B(n_1601),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1649),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1640),
.B(n_1601),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1640),
.B(n_1630),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1642),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1644),
.B(n_1599),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1642),
.Y(n_1673)
);

OAI21xp33_ASAP7_75t_L g1674 ( 
.A1(n_1652),
.A2(n_1596),
.B(n_1618),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1650),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1648),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1650),
.Y(n_1677)
);

AO21x2_ASAP7_75t_L g1678 ( 
.A1(n_1637),
.A2(n_1619),
.B(n_1618),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1639),
.Y(n_1679)
);

AOI211xp5_ASAP7_75t_L g1680 ( 
.A1(n_1638),
.A2(n_1615),
.B(n_1622),
.C(n_1600),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1660),
.B(n_1605),
.Y(n_1681)
);

NOR3xp33_ASAP7_75t_SL g1682 ( 
.A(n_1638),
.B(n_1505),
.C(n_1515),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1648),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1652),
.A2(n_1609),
.B1(n_1523),
.B2(n_1634),
.Y(n_1684)
);

OR2x2_ASAP7_75t_SL g1685 ( 
.A(n_1656),
.B(n_1635),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1644),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1659),
.B(n_1594),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1686),
.B(n_1643),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1673),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1664),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1673),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1668),
.Y(n_1692)
);

INVx2_ASAP7_75t_SL g1693 ( 
.A(n_1662),
.Y(n_1693)
);

NOR2x1_ASAP7_75t_L g1694 ( 
.A(n_1662),
.B(n_1657),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1663),
.B(n_1653),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1676),
.B(n_1659),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1668),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1663),
.B(n_1653),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1666),
.B(n_1641),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1676),
.B(n_1651),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1663),
.B(n_1660),
.Y(n_1701)
);

BUFx2_ASAP7_75t_L g1702 ( 
.A(n_1662),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_1662),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1665),
.B(n_1658),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1675),
.B(n_1647),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1677),
.B(n_1647),
.Y(n_1706)
);

AND2x6_ASAP7_75t_SL g1707 ( 
.A(n_1687),
.B(n_1593),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1683),
.B(n_1681),
.Y(n_1708)
);

NAND2x1p5_ASAP7_75t_L g1709 ( 
.A(n_1679),
.B(n_1658),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1683),
.B(n_1656),
.Y(n_1710)
);

NOR2x1p5_ASAP7_75t_L g1711 ( 
.A(n_1703),
.B(n_1661),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1689),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1710),
.A2(n_1674),
.B1(n_1661),
.B2(n_1680),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1708),
.B(n_1670),
.Y(n_1714)
);

INVx3_ASAP7_75t_L g1715 ( 
.A(n_1709),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1689),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1694),
.B(n_1658),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1708),
.B(n_1670),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1699),
.B(n_1669),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1705),
.B(n_1706),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1691),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1691),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1690),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1710),
.B(n_1670),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1699),
.B(n_1669),
.Y(n_1725)
);

INVx3_ASAP7_75t_L g1726 ( 
.A(n_1709),
.Y(n_1726)
);

OAI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1696),
.A2(n_1674),
.B(n_1680),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1696),
.B(n_1613),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1701),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1700),
.B(n_1671),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1690),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1694),
.B(n_1665),
.Y(n_1732)
);

INVx2_ASAP7_75t_SL g1733 ( 
.A(n_1709),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1700),
.B(n_1682),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1702),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1701),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1695),
.B(n_1685),
.Y(n_1737)
);

INVxp67_ASAP7_75t_SL g1738 ( 
.A(n_1688),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1695),
.B(n_1671),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1695),
.B(n_1672),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1701),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1704),
.B(n_1665),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1703),
.B(n_1705),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1703),
.B(n_1667),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1692),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1697),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1703),
.B(n_1667),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1705),
.B(n_1667),
.Y(n_1748)
);

INVxp67_ASAP7_75t_SL g1749 ( 
.A(n_1688),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1728),
.B(n_1568),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1744),
.B(n_1702),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1744),
.B(n_1702),
.Y(n_1752)
);

INVxp67_ASAP7_75t_L g1753 ( 
.A(n_1711),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1717),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1720),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1713),
.B(n_1687),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1724),
.B(n_1698),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1735),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1720),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1724),
.B(n_1698),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1747),
.B(n_1743),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1747),
.B(n_1693),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1712),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1720),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1712),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1713),
.B(n_1707),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_SL g1767 ( 
.A(n_1727),
.B(n_1735),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_SL g1768 ( 
.A(n_1727),
.B(n_1655),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1714),
.B(n_1698),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1716),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1723),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1716),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1743),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1721),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1721),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1722),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1714),
.B(n_1688),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_SL g1778 ( 
.A(n_1734),
.B(n_1682),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1722),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1745),
.Y(n_1780)
);

CKINVDCx16_ASAP7_75t_R g1781 ( 
.A(n_1737),
.Y(n_1781)
);

BUFx2_ASAP7_75t_L g1782 ( 
.A(n_1717),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1711),
.B(n_1707),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1737),
.B(n_1693),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1723),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1742),
.A2(n_1684),
.B1(n_1678),
.B2(n_1617),
.Y(n_1786)
);

OAI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1768),
.A2(n_1749),
.B(n_1738),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1782),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1758),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1753),
.B(n_1613),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1780),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1780),
.Y(n_1792)
);

A2O1A1Ixp33_ASAP7_75t_L g1793 ( 
.A1(n_1768),
.A2(n_1584),
.B(n_1749),
.C(n_1738),
.Y(n_1793)
);

OAI222xp33_ASAP7_75t_L g1794 ( 
.A1(n_1766),
.A2(n_1718),
.B1(n_1740),
.B2(n_1684),
.C1(n_1730),
.C2(n_1733),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1761),
.B(n_1751),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1781),
.B(n_1748),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1781),
.B(n_1748),
.Y(n_1797)
);

OAI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1767),
.A2(n_1631),
.B1(n_1685),
.B2(n_1718),
.Y(n_1798)
);

OAI21xp33_ASAP7_75t_L g1799 ( 
.A1(n_1767),
.A2(n_1730),
.B(n_1739),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1773),
.Y(n_1800)
);

NOR2x1_ASAP7_75t_L g1801 ( 
.A(n_1778),
.B(n_1783),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1756),
.B(n_1719),
.Y(n_1802)
);

INVxp67_ASAP7_75t_L g1803 ( 
.A(n_1751),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1763),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1763),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1761),
.B(n_1719),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1752),
.B(n_1725),
.Y(n_1807)
);

INVx1_ASAP7_75t_SL g1808 ( 
.A(n_1773),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1765),
.Y(n_1809)
);

OAI21xp5_ASAP7_75t_SL g1810 ( 
.A1(n_1786),
.A2(n_1732),
.B(n_1726),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1757),
.B(n_1740),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1752),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1795),
.B(n_1762),
.Y(n_1813)
);

OAI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1787),
.A2(n_1784),
.B1(n_1760),
.B2(n_1757),
.C(n_1782),
.Y(n_1814)
);

OAI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1793),
.A2(n_1762),
.B(n_1760),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1795),
.B(n_1755),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1788),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1790),
.B(n_1750),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1788),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1791),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1793),
.A2(n_1685),
.B1(n_1656),
.B2(n_1755),
.Y(n_1821)
);

INVx1_ASAP7_75t_SL g1822 ( 
.A(n_1795),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1803),
.B(n_1755),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1792),
.Y(n_1824)
);

INVxp67_ASAP7_75t_L g1825 ( 
.A(n_1789),
.Y(n_1825)
);

AND2x4_ASAP7_75t_SL g1826 ( 
.A(n_1790),
.B(n_1655),
.Y(n_1826)
);

INVx2_ASAP7_75t_SL g1827 ( 
.A(n_1807),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1804),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1805),
.Y(n_1829)
);

OAI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1799),
.A2(n_1769),
.B1(n_1759),
.B2(n_1764),
.C(n_1715),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1800),
.B(n_1759),
.Y(n_1831)
);

OAI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1798),
.A2(n_1764),
.B1(n_1759),
.B2(n_1769),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1822),
.B(n_1808),
.Y(n_1833)
);

OAI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1832),
.A2(n_1801),
.B(n_1798),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1819),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1819),
.Y(n_1836)
);

INVxp67_ASAP7_75t_L g1837 ( 
.A(n_1818),
.Y(n_1837)
);

INVx5_ASAP7_75t_L g1838 ( 
.A(n_1816),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1821),
.A2(n_1810),
.B1(n_1812),
.B2(n_1796),
.Y(n_1839)
);

INVxp67_ASAP7_75t_L g1840 ( 
.A(n_1818),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1826),
.Y(n_1841)
);

AOI211xp5_ASAP7_75t_L g1842 ( 
.A1(n_1814),
.A2(n_1794),
.B(n_1797),
.C(n_1802),
.Y(n_1842)
);

NAND2x1p5_ASAP7_75t_L g1843 ( 
.A(n_1817),
.B(n_1584),
.Y(n_1843)
);

AND2x4_ASAP7_75t_SL g1844 ( 
.A(n_1827),
.B(n_1607),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1833),
.B(n_1831),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1835),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1838),
.B(n_1825),
.Y(n_1847)
);

NAND3xp33_ASAP7_75t_L g1848 ( 
.A(n_1834),
.B(n_1825),
.C(n_1815),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1837),
.B(n_1823),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1838),
.B(n_1813),
.Y(n_1850)
);

AOI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1841),
.A2(n_1830),
.B1(n_1806),
.B2(n_1764),
.Y(n_1851)
);

NOR3xp33_ASAP7_75t_SL g1852 ( 
.A(n_1836),
.B(n_1824),
.C(n_1820),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1844),
.Y(n_1853)
);

AOI321xp33_ASAP7_75t_L g1854 ( 
.A1(n_1842),
.A2(n_1829),
.A3(n_1828),
.B1(n_1809),
.B2(n_1811),
.C(n_1754),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1843),
.B(n_1725),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1853),
.B(n_1838),
.Y(n_1856)
);

AOI321xp33_ASAP7_75t_L g1857 ( 
.A1(n_1851),
.A2(n_1839),
.A3(n_1840),
.B1(n_1754),
.B2(n_1774),
.C(n_1779),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_R g1858 ( 
.A(n_1850),
.B(n_1568),
.Y(n_1858)
);

AOI221xp5_ASAP7_75t_L g1859 ( 
.A1(n_1848),
.A2(n_1754),
.B1(n_1770),
.B2(n_1779),
.C(n_1765),
.Y(n_1859)
);

OAI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1852),
.A2(n_1847),
.B(n_1845),
.Y(n_1860)
);

AOI222xp33_ASAP7_75t_L g1861 ( 
.A1(n_1846),
.A2(n_1772),
.B1(n_1770),
.B2(n_1776),
.C1(n_1775),
.C2(n_1774),
.Y(n_1861)
);

OAI211xp5_ASAP7_75t_L g1862 ( 
.A1(n_1854),
.A2(n_1754),
.B(n_1590),
.C(n_1715),
.Y(n_1862)
);

NOR3xp33_ASAP7_75t_L g1863 ( 
.A(n_1849),
.B(n_1590),
.C(n_1542),
.Y(n_1863)
);

AOI221xp5_ASAP7_75t_L g1864 ( 
.A1(n_1860),
.A2(n_1855),
.B1(n_1772),
.B2(n_1776),
.C(n_1775),
.Y(n_1864)
);

INVxp67_ASAP7_75t_SL g1865 ( 
.A(n_1856),
.Y(n_1865)
);

OAI21xp5_ASAP7_75t_L g1866 ( 
.A1(n_1862),
.A2(n_1777),
.B(n_1733),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1863),
.A2(n_1715),
.B1(n_1726),
.B2(n_1742),
.Y(n_1867)
);

AOI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1859),
.A2(n_1715),
.B1(n_1726),
.B2(n_1732),
.Y(n_1868)
);

AOI322xp5_ASAP7_75t_L g1869 ( 
.A1(n_1857),
.A2(n_1733),
.A3(n_1739),
.B1(n_1729),
.B2(n_1741),
.C1(n_1736),
.C2(n_1726),
.Y(n_1869)
);

NAND3xp33_ASAP7_75t_SL g1870 ( 
.A(n_1858),
.B(n_1861),
.C(n_1577),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1865),
.B(n_1777),
.Y(n_1871)
);

NAND4xp75_ASAP7_75t_L g1872 ( 
.A(n_1864),
.B(n_1785),
.C(n_1771),
.D(n_1693),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1870),
.B(n_1511),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1866),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1867),
.B(n_1742),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1868),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1874),
.B(n_1869),
.Y(n_1877)
);

XOR2x2_ASAP7_75t_L g1878 ( 
.A(n_1871),
.B(n_1511),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1876),
.B(n_1729),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1878),
.B(n_1873),
.Y(n_1880)
);

OAI22x1_ASAP7_75t_L g1881 ( 
.A1(n_1880),
.A2(n_1873),
.B1(n_1877),
.B2(n_1879),
.Y(n_1881)
);

OAI21xp33_ASAP7_75t_L g1882 ( 
.A1(n_1881),
.A2(n_1875),
.B(n_1872),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1881),
.A2(n_1785),
.B1(n_1771),
.B2(n_1736),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1882),
.B(n_1771),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1883),
.Y(n_1885)
);

OAI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1884),
.A2(n_1785),
.B(n_1741),
.Y(n_1886)
);

OAI21xp33_ASAP7_75t_L g1887 ( 
.A1(n_1885),
.A2(n_1542),
.B(n_1580),
.Y(n_1887)
);

OA22x2_ASAP7_75t_L g1888 ( 
.A1(n_1886),
.A2(n_1593),
.B1(n_1732),
.B2(n_1731),
.Y(n_1888)
);

OAI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1888),
.A2(n_1887),
.B(n_1627),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1889),
.Y(n_1890)
);

AOI221xp5_ASAP7_75t_L g1891 ( 
.A1(n_1890),
.A2(n_1723),
.B1(n_1731),
.B2(n_1745),
.C(n_1746),
.Y(n_1891)
);

AOI211xp5_ASAP7_75t_L g1892 ( 
.A1(n_1891),
.A2(n_1570),
.B(n_1592),
.C(n_1731),
.Y(n_1892)
);


endmodule