module real_jpeg_8860_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_1),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g94 ( 
.A1(n_1),
.A2(n_3),
.B(n_61),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_1),
.A2(n_71),
.B1(n_76),
.B2(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_1),
.B(n_110),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_1),
.A2(n_39),
.B(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_1),
.B(n_39),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_1),
.A2(n_27),
.B1(n_34),
.B2(n_160),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_1),
.A2(n_60),
.B(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_1),
.B(n_60),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_2),
.A2(n_71),
.B1(n_76),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_2),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_2),
.A2(n_60),
.B1(n_61),
.B2(n_89),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_89),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_89),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_3),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_3),
.A2(n_60),
.B1(n_61),
.B2(n_72),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_7),
.A2(n_60),
.B(n_62),
.C(n_63),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_7),
.B(n_60),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_7),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_10),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_56),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_11),
.A2(n_60),
.B1(n_61),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_11),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_11),
.A2(n_39),
.B1(n_40),
.B2(n_66),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_66),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_12),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_12),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_12),
.A2(n_60),
.B1(n_61),
.B2(n_77),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_77),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_12),
.A2(n_39),
.B1(n_40),
.B2(n_77),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_15),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_15),
.A2(n_30),
.B1(n_31),
.B2(n_41),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_16),
.A2(n_39),
.B1(n_40),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_16),
.A2(n_30),
.B1(n_31),
.B2(n_48),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_17),
.A2(n_71),
.B1(n_76),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_17),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_17),
.A2(n_60),
.B1(n_61),
.B2(n_79),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_17),
.A2(n_30),
.B1(n_31),
.B2(n_79),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_17),
.A2(n_39),
.B1(n_40),
.B2(n_79),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_117),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_116),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_99),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_22),
.B(n_99),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_81),
.B2(n_98),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_49),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_37),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_27),
.A2(n_32),
.B1(n_34),
.B2(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_27),
.A2(n_34),
.B1(n_52),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_27),
.A2(n_34),
.B1(n_143),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_27),
.A2(n_34),
.B1(n_145),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_27),
.A2(n_34),
.B1(n_176),
.B2(n_192),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_28),
.A2(n_29),
.B1(n_97),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_28),
.A2(n_29),
.B1(n_142),
.B2(n_144),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_30),
.A2(n_31),
.B1(n_43),
.B2(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_30),
.B(n_46),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_30),
.B(n_165),
.Y(n_164)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_31),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_34),
.B(n_93),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_42),
.B1(n_45),
.B2(n_54),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_43),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_39),
.B(n_64),
.Y(n_189)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_40),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_187)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_42),
.A2(n_45),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_42),
.A2(n_45),
.B1(n_151),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_42),
.A2(n_45),
.B1(n_174),
.B2(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_42),
.A2(n_45),
.B1(n_113),
.B2(n_182),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_44),
.Y(n_155)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_45),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_45),
.B(n_93),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_57),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_53),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_55),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_68),
.B1(n_69),
.B2(n_80),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_59),
.A2(n_63),
.B1(n_84),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_59),
.A2(n_63),
.B1(n_106),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_59),
.A2(n_63),
.B1(n_129),
.B2(n_184),
.Y(n_183)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_62),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_63),
.B(n_93),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_74),
.B1(n_75),
.B2(n_78),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_74),
.B1(n_75),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B(n_73),
.C(n_74),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_72),
.Y(n_73)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_72),
.B(n_93),
.C(n_94),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_74),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_81),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_85),
.C(n_90),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.C(n_103),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_103),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.C(n_111),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_105),
.B1(n_111),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_111),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_135),
.B(n_214),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_133),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_119),
.B(n_133),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.C(n_125),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_120),
.B(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_123),
.A2(n_125),
.B1(n_126),
.B2(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_123),
.Y(n_212)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.C(n_131),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_127),
.A2(n_128),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_130),
.B(n_131),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_132),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_208),
.B(n_213),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_194),
.B(n_207),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_178),
.B(n_193),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_168),
.B(n_177),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_157),
.B(n_167),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_146),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_141),
.B(n_146),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_152),
.B2(n_156),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_147),
.B(n_156),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_150),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_152),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_162),
.B(n_166),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_161),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_169),
.B(n_170),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_173),
.C(n_175),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_180),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_180),
.Y(n_195)
);

FAx1_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_183),
.CI(n_186),
.CON(n_180),
.SN(n_180)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_185),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_191),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_195),
.B(n_196),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_204),
.C(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_203),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_204),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_209),
.B(n_210),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);


endmodule