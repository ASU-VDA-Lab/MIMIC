module fake_jpeg_27325_n_164 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx4f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_14),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_28),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_11),
.B1(n_13),
.B2(n_17),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_19),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_24),
.A2(n_11),
.B1(n_15),
.B2(n_19),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_11),
.B1(n_20),
.B2(n_18),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_46),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_31),
.B(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_39),
.B1(n_33),
.B2(n_30),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_54),
.B1(n_42),
.B2(n_49),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_48),
.A2(n_39),
.B1(n_30),
.B2(n_32),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_39),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_64),
.B1(n_65),
.B2(n_57),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_43),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_71),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_50),
.B1(n_51),
.B2(n_44),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_70),
.B1(n_66),
.B2(n_60),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_50),
.B1(n_51),
.B2(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_75),
.Y(n_87)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_64),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_37),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_59),
.C(n_37),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_40),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_69),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_77),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_86),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_63),
.B1(n_59),
.B2(n_57),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_84),
.B1(n_79),
.B2(n_78),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_76),
.C(n_79),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_91),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_0),
.B(n_1),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NOR3xp33_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_61),
.C(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_94),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_76),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_103),
.C(n_91),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_90),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_105),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_99),
.A2(n_104),
.B1(n_84),
.B2(n_82),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_71),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_102),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_83),
.B1(n_88),
.B2(n_86),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_87),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_68),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_70),
.B1(n_61),
.B2(n_31),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_74),
.Y(n_105)
);

BUFx24_ASAP7_75t_SL g106 ( 
.A(n_102),
.Y(n_106)
);

BUFx24_ASAP7_75t_SL g123 ( 
.A(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_103),
.B(n_80),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_115),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_117),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_25),
.B1(n_24),
.B2(n_13),
.Y(n_126)
);

INVxp33_ASAP7_75t_SL g112 ( 
.A(n_93),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_112),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_94),
.C(n_28),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_20),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_28),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

AO21x1_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_16),
.B(n_21),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_17),
.B(n_21),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_122),
.B1(n_110),
.B2(n_7),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_98),
.B1(n_96),
.B2(n_100),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_28),
.C(n_27),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g133 ( 
.A(n_125),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_129),
.B1(n_0),
.B2(n_1),
.Y(n_136)
);

AOI31xp67_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_13),
.A3(n_20),
.B(n_18),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_107),
.B(n_13),
.C(n_18),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_18),
.B1(n_20),
.B2(n_8),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_110),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_131),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_128),
.B(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_136),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_138),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_28),
.Y(n_138)
);

OAI21x1_ASAP7_75t_SL g140 ( 
.A1(n_138),
.A2(n_127),
.B(n_119),
.Y(n_140)
);

OAI321xp33_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_144),
.A3(n_132),
.B1(n_7),
.B2(n_9),
.C(n_4),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_27),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_146),
.Y(n_151)
);

AOI31xp67_ASAP7_75t_SL g144 ( 
.A1(n_133),
.A2(n_123),
.A3(n_8),
.B(n_9),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_147),
.A2(n_151),
.B1(n_2),
.B2(n_3),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_145),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_149),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_141),
.A2(n_7),
.B1(n_10),
.B2(n_9),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_6),
.B(n_10),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_150),
.A2(n_0),
.B(n_2),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_27),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_27),
.C(n_28),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_27),
.Y(n_160)
);

FAx1_ASAP7_75t_SL g154 ( 
.A(n_152),
.B(n_4),
.CI(n_10),
.CON(n_154),
.SN(n_154)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_156),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_157),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_160),
.C(n_153),
.Y(n_161)
);

OAI21x1_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_162),
.B(n_154),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_154),
.C(n_3),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_3),
.Y(n_164)
);


endmodule