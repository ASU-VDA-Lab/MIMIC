module fake_aes_2151_n_16 (n_1, n_2, n_0, n_16);
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
NOR2x1_ASAP7_75t_L g4 ( .A(n_0), .B(n_1), .Y(n_4) );
NAND2x1p5_ASAP7_75t_L g5 ( .A(n_3), .B(n_0), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g6 ( .A(n_3), .B(n_4), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
INVx2_ASAP7_75t_R g8 ( .A(n_6), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
NOR2xp33_ASAP7_75t_SL g10 ( .A(n_7), .B(n_0), .Y(n_10) );
NOR3xp33_ASAP7_75t_SL g11 ( .A(n_10), .B(n_8), .C(n_1), .Y(n_11) );
O2A1O1Ixp33_ASAP7_75t_L g12 ( .A1(n_9), .A2(n_8), .B(n_2), .C(n_0), .Y(n_12) );
NAND2x1p5_ASAP7_75t_L g13 ( .A(n_11), .B(n_9), .Y(n_13) );
NAND2xp33_ASAP7_75t_SL g14 ( .A(n_12), .B(n_8), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_13), .B(n_2), .Y(n_15) );
OAI21xp5_ASAP7_75t_L g16 ( .A1(n_15), .A2(n_14), .B(n_2), .Y(n_16) );
endmodule