module fake_netlist_5_1864_n_458 (n_91, n_82, n_122, n_10, n_24, n_124, n_86, n_83, n_61, n_90, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_105, n_80, n_4, n_35, n_73, n_17, n_92, n_19, n_120, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_458);

input n_91;
input n_82;
input n_122;
input n_10;
input n_24;
input n_124;
input n_86;
input n_83;
input n_61;
input n_90;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_105;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_458;

wire n_137;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_444;
wire n_194;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_136;
wire n_146;
wire n_315;
wire n_268;
wire n_451;
wire n_408;
wire n_376;
wire n_127;
wire n_235;
wire n_226;
wire n_353;
wire n_351;
wire n_367;
wire n_452;
wire n_397;
wire n_155;
wire n_423;
wire n_284;
wire n_245;
wire n_139;
wire n_280;
wire n_378;
wire n_382;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_321;
wire n_292;
wire n_455;
wire n_417;
wire n_212;
wire n_385;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_330;
wire n_373;
wire n_147;
wire n_307;
wire n_439;
wire n_150;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_186;
wire n_134;
wire n_191;
wire n_171;
wire n_153;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_325;
wire n_449;
wire n_132;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_152;
wire n_317;
wire n_323;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_335;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_457;
wire n_297;
wire n_156;
wire n_225;
wire n_377;
wire n_219;
wire n_442;
wire n_157;
wire n_131;
wire n_192;
wire n_223;
wire n_392;
wire n_158;
wire n_138;
wire n_264;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_287;
wire n_344;
wire n_422;
wire n_415;
wire n_141;
wire n_355;
wire n_336;
wire n_145;
wire n_337;
wire n_430;
wire n_313;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_165;
wire n_213;
wire n_129;
wire n_342;
wire n_361;
wire n_363;
wire n_402;
wire n_413;
wire n_197;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_277;
wire n_338;
wire n_149;
wire n_333;
wire n_309;
wire n_130;
wire n_322;
wire n_258;
wire n_151;
wire n_306;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_239;
wire n_420;
wire n_310;
wire n_358;
wire n_362;
wire n_332;
wire n_170;
wire n_273;
wire n_161;
wire n_349;
wire n_270;
wire n_230;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_441;
wire n_450;
wire n_312;
wire n_429;
wire n_345;
wire n_210;
wire n_365;
wire n_176;
wire n_182;
wire n_143;
wire n_354;
wire n_237;
wire n_425;
wire n_407;
wire n_180;
wire n_340;
wire n_207;
wire n_346;
wire n_393;
wire n_229;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_405;
wire n_359;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_246;
wire n_179;
wire n_125;
wire n_410;
wire n_269;
wire n_128;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_426;
wire n_409;
wire n_154;
wire n_148;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_391;
wire n_434;
wire n_175;
wire n_262;
wire n_238;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_242;
wire n_360;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_278;

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

INVxp67_ASAP7_75t_SL g127 ( 
.A(n_114),
.Y(n_127)
);

NOR2xp67_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_8),
.Y(n_128)
);

INVxp33_ASAP7_75t_SL g129 ( 
.A(n_17),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

INVxp67_ASAP7_75t_SL g133 ( 
.A(n_56),
.Y(n_133)
);

INVxp67_ASAP7_75t_SL g134 ( 
.A(n_48),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_86),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_52),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_3),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_51),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_0),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_7),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_107),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_23),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_3),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_27),
.Y(n_150)
);

INVxp33_ASAP7_75t_SL g151 ( 
.A(n_92),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_96),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_40),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_2),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_42),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_73),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_41),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_5),
.Y(n_158)
);

INVxp67_ASAP7_75t_SL g159 ( 
.A(n_66),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_75),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_84),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_102),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_32),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_16),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_74),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_5),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_34),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_79),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_55),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_10),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_90),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_64),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_54),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_95),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_30),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_46),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_10),
.Y(n_183)
);

INVxp67_ASAP7_75t_SL g184 ( 
.A(n_99),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_72),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_62),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_2),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_31),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_19),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_29),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_57),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_58),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_77),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_18),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_9),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_83),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_37),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_12),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_139),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_0),
.B(n_1),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_145),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_144),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_1),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_169),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_154),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_157),
.B(n_125),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_155),
.B(n_4),
.Y(n_214)
);

AND2x4_ASAP7_75t_L g215 ( 
.A(n_125),
.B(n_13),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_153),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_165),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_180),
.B(n_4),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_164),
.B(n_194),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_172),
.B(n_6),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_130),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_135),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_126),
.B(n_6),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_136),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_131),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_132),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_178),
.B(n_7),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_178),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_212),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_129),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_8),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_127),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_208),
.A2(n_151),
.B1(n_128),
.B2(n_146),
.Y(n_247)
);

AND2x4_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_127),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_167),
.B1(n_181),
.B2(n_159),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

AND2x6_ASAP7_75t_L g252 ( 
.A(n_201),
.B(n_140),
.Y(n_252)
);

BUFx4f_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_199),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_207),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_220),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_220),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_200),
.B(n_215),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_225),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_214),
.A2(n_133),
.B1(n_134),
.B2(n_159),
.Y(n_263)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_215),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_222),
.B(n_214),
.Y(n_266)
);

NAND3xp33_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_147),
.C(n_137),
.Y(n_267)
);

BUFx4f_ASAP7_75t_L g268 ( 
.A(n_201),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_221),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_230),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_228),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_227),
.A2(n_224),
.B1(n_231),
.B2(n_200),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_200),
.B(n_141),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_229),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_232),
.Y(n_275)
);

AND2x6_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_142),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_240),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

BUFx8_ASAP7_75t_L g280 ( 
.A(n_244),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_235),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_223),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_266),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_210),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_251),
.Y(n_286)
);

AND2x4_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_202),
.Y(n_287)
);

AND2x4_ASAP7_75t_L g288 ( 
.A(n_248),
.B(n_246),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_255),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_259),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_259),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_247),
.B(n_150),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_223),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_245),
.B(n_210),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_133),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_251),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_258),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_269),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_269),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_258),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_237),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_249),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_264),
.B(n_134),
.Y(n_309)
);

OR2x6_ASAP7_75t_L g310 ( 
.A(n_239),
.B(n_205),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_238),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_242),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_258),
.Y(n_313)
);

NOR3xp33_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_147),
.C(n_184),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_262),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_253),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_243),
.A2(n_184),
.B1(n_197),
.B2(n_161),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_246),
.B(n_233),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_265),
.B(n_206),
.Y(n_319)
);

O2A1O1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_270),
.A2(n_216),
.B(n_209),
.C(n_218),
.Y(n_320)
);

A2O1A1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_284),
.A2(n_268),
.B(n_288),
.C(n_281),
.Y(n_321)
);

INVx5_ASAP7_75t_L g322 ( 
.A(n_316),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_315),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_204),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_287),
.B(n_291),
.Y(n_326)
);

NAND2x1p5_ASAP7_75t_L g327 ( 
.A(n_287),
.B(n_316),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_279),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_314),
.A2(n_283),
.B1(n_252),
.B2(n_296),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_299),
.A2(n_250),
.B(n_241),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_301),
.A2(n_309),
.B1(n_317),
.B2(n_308),
.Y(n_332)
);

AND2x4_ASAP7_75t_L g333 ( 
.A(n_290),
.B(n_218),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_252),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_285),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_310),
.A2(n_219),
.B(n_226),
.C(n_204),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_294),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_292),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_278),
.Y(n_340)
);

AOI21xp33_ASAP7_75t_L g341 ( 
.A1(n_310),
.A2(n_203),
.B(n_143),
.Y(n_341)
);

CKINVDCx6p67_ASAP7_75t_R g342 ( 
.A(n_293),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_289),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_297),
.B(n_148),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_278),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_316),
.B(n_152),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_304),
.B(n_300),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_282),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_307),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_311),
.B(n_160),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_312),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_306),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_295),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_298),
.B(n_162),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_282),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_313),
.Y(n_357)
);

INVx8_ASAP7_75t_L g358 ( 
.A(n_277),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_326),
.B(n_347),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_324),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_338),
.Y(n_361)
);

OA21x2_ASAP7_75t_L g362 ( 
.A1(n_341),
.A2(n_193),
.B(n_166),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_343),
.Y(n_363)
);

AOI221xp5_ASAP7_75t_SL g364 ( 
.A1(n_337),
.A2(n_321),
.B1(n_329),
.B2(n_338),
.C(n_332),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_328),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_348),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_333),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_325),
.A2(n_280),
.B1(n_203),
.B2(n_170),
.Y(n_368)
);

OAI22xp33_ASAP7_75t_L g369 ( 
.A1(n_325),
.A2(n_188),
.B1(n_168),
.B2(n_171),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_335),
.A2(n_320),
.B(n_286),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_345),
.A2(n_190),
.B1(n_179),
.B2(n_182),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_340),
.A2(n_191),
.B1(n_185),
.B2(n_186),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_336),
.B(n_280),
.Y(n_373)
);

O2A1O1Ixp33_ASAP7_75t_SL g374 ( 
.A1(n_346),
.A2(n_192),
.B(n_173),
.C(n_177),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_339),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_331),
.A2(n_303),
.B(n_302),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_330),
.A2(n_198),
.B1(n_176),
.B2(n_175),
.Y(n_377)
);

O2A1O1Ixp33_ASAP7_75t_L g378 ( 
.A1(n_334),
.A2(n_233),
.B(n_303),
.C(n_302),
.Y(n_378)
);

AOI221xp5_ASAP7_75t_L g379 ( 
.A1(n_350),
.A2(n_219),
.B1(n_226),
.B2(n_233),
.C(n_156),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_L g380 ( 
.A1(n_322),
.A2(n_163),
.B1(n_286),
.B2(n_313),
.Y(n_380)
);

OAI222xp33_ASAP7_75t_L g381 ( 
.A1(n_327),
.A2(n_9),
.B1(n_11),
.B2(n_14),
.C1(n_15),
.C2(n_20),
.Y(n_381)
);

OAI221xp5_ASAP7_75t_L g382 ( 
.A1(n_351),
.A2(n_11),
.B1(n_276),
.B2(n_22),
.C(n_24),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_347),
.B(n_276),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_350),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_361),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_377),
.A2(n_382),
.B1(n_368),
.B2(n_365),
.Y(n_386)
);

AOI222xp33_ASAP7_75t_L g387 ( 
.A1(n_381),
.A2(n_326),
.B1(n_358),
.B2(n_354),
.C1(n_344),
.C2(n_323),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_354),
.Y(n_388)
);

OAI21x1_ASAP7_75t_L g389 ( 
.A1(n_376),
.A2(n_356),
.B(n_339),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_359),
.A2(n_358),
.B1(n_322),
.B2(n_344),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_375),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_360),
.A2(n_349),
.B1(n_353),
.B2(n_352),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_379),
.A2(n_342),
.B1(n_322),
.B2(n_348),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_367),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_384),
.B(n_355),
.Y(n_395)
);

OAI22xp33_ASAP7_75t_L g396 ( 
.A1(n_363),
.A2(n_357),
.B1(n_355),
.B2(n_26),
.Y(n_396)
);

OAI22xp33_ASAP7_75t_L g397 ( 
.A1(n_383),
.A2(n_373),
.B1(n_369),
.B2(n_379),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_L g398 ( 
.A1(n_362),
.A2(n_357),
.B1(n_25),
.B2(n_28),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_366),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_362),
.A2(n_21),
.B1(n_33),
.B2(n_35),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_378),
.A2(n_36),
.B(n_38),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_364),
.Y(n_402)
);

AOI221xp5_ASAP7_75t_L g403 ( 
.A1(n_397),
.A2(n_372),
.B1(n_371),
.B2(n_374),
.C(n_380),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_385),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_394),
.B(n_370),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_391),
.Y(n_406)
);

OAI31xp33_ASAP7_75t_L g407 ( 
.A1(n_396),
.A2(n_39),
.A3(n_43),
.B(n_44),
.Y(n_407)
);

OAI221xp5_ASAP7_75t_L g408 ( 
.A1(n_393),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.C(n_50),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_391),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_389),
.Y(n_410)
);

AOI221xp5_ASAP7_75t_L g411 ( 
.A1(n_393),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.C(n_63),
.Y(n_411)
);

NAND3xp33_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_65),
.C(n_67),
.Y(n_412)
);

AOI21xp33_ASAP7_75t_L g413 ( 
.A1(n_402),
.A2(n_68),
.B(n_69),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_388),
.B(n_70),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_412),
.A2(n_390),
.B1(n_386),
.B2(n_408),
.Y(n_415)
);

AO21x2_ASAP7_75t_L g416 ( 
.A1(n_410),
.A2(n_400),
.B(n_401),
.Y(n_416)
);

OAI31xp33_ASAP7_75t_L g417 ( 
.A1(n_408),
.A2(n_386),
.A3(n_398),
.B(n_395),
.Y(n_417)
);

AND2x2_ASAP7_75t_SL g418 ( 
.A(n_411),
.B(n_395),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_414),
.B(n_392),
.Y(n_419)
);

NAND3xp33_ASAP7_75t_SL g420 ( 
.A(n_403),
.B(n_392),
.C(n_399),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_404),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_406),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_409),
.Y(n_423)
);

OAI31xp33_ASAP7_75t_L g424 ( 
.A1(n_407),
.A2(n_80),
.A3(n_81),
.B(n_82),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_405),
.B(n_85),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_413),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_413),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_421),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_419),
.B(n_88),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_422),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_423),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_425),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_427),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_91),
.Y(n_434)
);

OR2x6_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_94),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_426),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_420),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_429),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_433),
.B(n_416),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_433),
.B(n_417),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_424),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_435),
.A2(n_97),
.B(n_101),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_442),
.A2(n_435),
.B(n_437),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_438),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_439),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_443),
.A2(n_435),
.B1(n_441),
.B2(n_440),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_445),
.B(n_436),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_446),
.A2(n_444),
.B1(n_436),
.B2(n_434),
.Y(n_448)
);

O2A1O1Ixp33_ASAP7_75t_L g449 ( 
.A1(n_447),
.A2(n_428),
.B(n_430),
.C(n_431),
.Y(n_449)
);

OAI21xp33_ASAP7_75t_SL g450 ( 
.A1(n_448),
.A2(n_449),
.B(n_108),
.Y(n_450)
);

XOR2x1_ASAP7_75t_L g451 ( 
.A(n_450),
.B(n_110),
.Y(n_451)
);

NOR3x2_ASAP7_75t_L g452 ( 
.A(n_451),
.B(n_111),
.C(n_112),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_452),
.A2(n_113),
.B1(n_115),
.B2(n_118),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_452),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_454),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_455),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_456),
.Y(n_457)
);

AOI221xp5_ASAP7_75t_L g458 ( 
.A1(n_457),
.A2(n_453),
.B1(n_120),
.B2(n_121),
.C(n_122),
.Y(n_458)
);


endmodule