module real_jpeg_359_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_1),
.A2(n_59),
.B1(n_60),
.B2(n_72),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_1),
.A2(n_39),
.B1(n_41),
.B2(n_72),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_72),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_2),
.A2(n_27),
.B1(n_39),
.B2(n_41),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_2),
.A2(n_27),
.B1(n_59),
.B2(n_60),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_2),
.A2(n_27),
.B1(n_71),
.B2(n_73),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_4),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_4),
.A2(n_34),
.B1(n_71),
.B2(n_73),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_4),
.A2(n_34),
.B1(n_59),
.B2(n_60),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_9),
.A2(n_38),
.B1(n_59),
.B2(n_60),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_38),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_9),
.A2(n_38),
.B1(n_71),
.B2(n_73),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_9),
.B(n_60),
.C(n_68),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_9),
.B(n_66),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_9),
.B(n_39),
.C(n_54),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_9),
.B(n_23),
.C(n_45),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_9),
.B(n_52),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_9),
.B(n_30),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_9),
.B(n_50),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_309),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_271),
.B(n_306),
.Y(n_14)
);

A2O1A1O1Ixp25_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_133),
.B(n_251),
.C(n_252),
.D(n_270),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_111),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_17),
.B(n_111),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_78),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_18),
.B(n_79),
.C(n_105),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_51),
.C(n_63),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_19),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_20),
.B(n_35),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_28),
.B(n_31),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_21),
.A2(n_29),
.B(n_86),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_22),
.A2(n_23),
.B1(n_44),
.B2(n_45),
.Y(n_47)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_23),
.B(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_28),
.B(n_33),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_28),
.A2(n_29),
.B(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_28),
.B(n_85),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_28),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_29),
.B(n_215),
.Y(n_229)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_30),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_31),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_32),
.B(n_214),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_48),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_36),
.B(n_200),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_42),
.Y(n_36)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_37),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_37),
.B(n_50),
.Y(n_186)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_41),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_39),
.B(n_209),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_42),
.B(n_49),
.Y(n_90)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_42),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

OAI21x1_ASAP7_75t_R g108 ( 
.A1(n_48),
.A2(n_89),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_48),
.B(n_187),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_50),
.B(n_188),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_51),
.A2(n_63),
.B1(n_64),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_51),
.A2(n_115),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_56),
.B(n_62),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_52),
.B(n_62),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_52),
.B(n_126),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_52),
.A2(n_152),
.B(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_54),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_56),
.B(n_62),
.Y(n_103)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_57),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_57),
.B(n_101),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_57),
.A2(n_285),
.B(n_286),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_60),
.B(n_183),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_74),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_66),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_66),
.B(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_66),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_73),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_75),
.Y(n_97)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_71),
.B(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_74),
.A2(n_263),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_104),
.B2(n_105),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_91),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_81),
.B(n_92),
.C(n_99),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_87),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_82),
.B(n_87),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_83),
.B(n_213),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_86),
.B(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B(n_90),
.Y(n_87)
);

AOI21x1_ASAP7_75t_SL g149 ( 
.A1(n_88),
.A2(n_109),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_90),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_90),
.B(n_186),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_98),
.B2(n_99),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_96),
.B(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_96),
.A2(n_147),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_100),
.B(n_124),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_100),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_103),
.B(n_154),
.Y(n_201)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_106),
.A2(n_107),
.B1(n_181),
.B2(n_182),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_106),
.A2(n_107),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_107),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_107),
.B(n_108),
.Y(n_259)
);

AOI21xp33_ASAP7_75t_L g275 ( 
.A1(n_107),
.A2(n_259),
.B(n_261),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_108),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_132),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_113),
.B1(n_132),
.B2(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.C(n_127),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_119),
.B(n_281),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_119),
.A2(n_147),
.B(n_299),
.Y(n_313)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_122),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_128),
.A2(n_129),
.B1(n_131),
.B2(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

OAI21x1_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_155),
.B(n_248),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_135),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_136),
.B(n_139),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_143),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_143),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.C(n_151),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_146),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_148),
.A2(n_149),
.B1(n_151),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_148),
.A2(n_149),
.B1(n_284),
.B2(n_287),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_148),
.A2(n_149),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_149),
.B(n_279),
.C(n_284),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_149),
.B(n_303),
.C(n_305),
.Y(n_315)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_152),
.B(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_173),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_157),
.B(n_159),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.C(n_166),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_160),
.A2(n_161),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_166),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.C(n_169),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_172),
.B(n_229),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_192),
.B(n_247),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_189),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_175),
.B(n_189),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_180),
.C(n_184),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_177),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_180),
.A2(n_184),
.B1(n_185),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI21x1_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_203),
.B(n_246),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_194),
.B(n_198),
.Y(n_246)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.C(n_202),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_201),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_241),
.B(n_245),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_223),
.B(n_240),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_211),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_216),
.B1(n_217),
.B2(n_222),
.Y(n_211)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_220),
.C(n_222),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_230),
.B(n_239),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_227),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_235),
.B(n_238),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_237),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_243),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_254),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_257),
.C(n_265),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_264),
.B2(n_265),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B(n_269),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_267),
.Y(n_269)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_269),
.A2(n_277),
.B1(n_278),
.B2(n_288),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_269),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_275),
.C(n_277),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_289),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_273),
.B(n_274),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_279),
.A2(n_280),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_280),
.B(n_292),
.C(n_296),
.Y(n_316)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_284),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_289),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_291),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_300),
.B1(n_301),
.B2(n_305),
.Y(n_297)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_317),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_316),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_311),
.B(n_316),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_315),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_313),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);


endmodule