module fake_jpeg_12860_n_491 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_491);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_491;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_61),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_57),
.Y(n_134)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_19),
.B(n_11),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_65),
.B(n_69),
.Y(n_125)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_19),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_71),
.B(n_72),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_77),
.B(n_80),
.Y(n_133)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_27),
.B(n_17),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_37),
.B(n_16),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_84),
.B(n_85),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_27),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_34),
.B(n_17),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_93),
.B(n_97),
.Y(n_146)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_34),
.B(n_17),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

BUFx8_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

BUFx16f_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_70),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_100),
.B(n_101),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_60),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_28),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_110),
.B(n_151),
.C(n_18),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_40),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_111),
.B(n_124),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_66),
.A2(n_39),
.B1(n_28),
.B2(n_40),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_120),
.A2(n_94),
.B1(n_53),
.B2(n_52),
.Y(n_160)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_68),
.A2(n_35),
.B(n_48),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_122),
.A2(n_26),
.B(n_35),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_41),
.Y(n_124)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_98),
.B(n_48),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_153),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_71),
.A2(n_46),
.B(n_58),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_98),
.B(n_26),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_157),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_99),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_159),
.B(n_162),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_160),
.A2(n_51),
.B1(n_134),
.B2(n_102),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_106),
.B(n_49),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_57),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_49),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_169),
.B(n_178),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

HAxp5_ASAP7_75t_SL g172 ( 
.A(n_149),
.B(n_68),
.CON(n_172),
.SN(n_172)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_172),
.A2(n_206),
.B(n_159),
.Y(n_213)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_173),
.Y(n_242)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_177),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_99),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_113),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_181),
.Y(n_228)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_116),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_182),
.Y(n_225)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_185),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_106),
.B(n_49),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_186),
.B(n_192),
.Y(n_229)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_104),
.Y(n_188)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_140),
.Y(n_191)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_43),
.B1(n_114),
.B2(n_55),
.Y(n_220)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_195),
.Y(n_231)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_129),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_115),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_197),
.Y(n_239)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_198),
.B(n_200),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_110),
.B(n_67),
.C(n_60),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_199),
.B(n_204),
.C(n_18),
.Y(n_250)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_129),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_205),
.Y(n_249)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_130),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_133),
.B(n_64),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_109),
.Y(n_205)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_127),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_207),
.A2(n_209),
.B1(n_192),
.B2(n_165),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_133),
.B(n_41),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_36),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_114),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_213),
.A2(n_29),
.B(n_165),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_183),
.A2(n_123),
.B1(n_131),
.B2(n_89),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_218),
.A2(n_219),
.B1(n_223),
.B2(n_238),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_167),
.A2(n_123),
.B1(n_131),
.B2(n_142),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_220),
.B(n_248),
.C(n_31),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_160),
.A2(n_87),
.B1(n_155),
.B2(n_130),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_233),
.B(n_15),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_236),
.A2(n_244),
.B1(n_172),
.B2(n_192),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_142),
.B1(n_109),
.B2(n_136),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_177),
.A2(n_155),
.B1(n_136),
.B2(n_62),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_243),
.A2(n_252),
.B1(n_254),
.B2(n_219),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_169),
.A2(n_138),
.B1(n_91),
.B2(n_86),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_158),
.B(n_145),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_138),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_168),
.A2(n_63),
.B1(n_96),
.B2(n_92),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_161),
.A2(n_79),
.B1(n_74),
.B2(n_75),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_228),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_255),
.B(n_266),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_215),
.B(n_158),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_256),
.B(n_262),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_257),
.A2(n_267),
.B1(n_271),
.B2(n_281),
.Y(n_323)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_217),
.Y(n_259)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_178),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_260),
.B(n_264),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_213),
.A2(n_31),
.B(n_18),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_261),
.A2(n_287),
.B(n_291),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_170),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_212),
.Y(n_263)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_263),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_173),
.Y(n_264)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_212),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_265),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_215),
.B(n_36),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_235),
.A2(n_203),
.B1(n_157),
.B2(n_82),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_226),
.Y(n_268)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_217),
.Y(n_269)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_270),
.A2(n_253),
.B1(n_221),
.B2(n_227),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_235),
.A2(n_152),
.B1(n_105),
.B2(n_59),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_272),
.B(n_276),
.C(n_288),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_218),
.A2(n_144),
.B1(n_171),
.B2(n_188),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_273),
.A2(n_242),
.B1(n_232),
.B2(n_234),
.Y(n_301)
);

O2A1O1Ixp33_ASAP7_75t_L g274 ( 
.A1(n_239),
.A2(n_145),
.B(n_31),
.C(n_113),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_274),
.B(n_279),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_216),
.B(n_181),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_278),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_67),
.C(n_39),
.Y(n_276)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_277),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_231),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_210),
.B(n_29),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_237),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_222),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_284),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_230),
.Y(n_283)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_283),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_226),
.Y(n_285)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_285),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_216),
.B(n_30),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_289),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_222),
.B(n_128),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_220),
.B(n_39),
.C(n_47),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_224),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_230),
.Y(n_290)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_290),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_238),
.B(n_29),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_240),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_295),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_229),
.B(n_47),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_293),
.Y(n_305)
);

CKINVDCx12_ASAP7_75t_R g294 ( 
.A(n_221),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_294),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_249),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_233),
.B(n_47),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_296),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_L g346 ( 
.A1(n_301),
.A2(n_312),
.B1(n_287),
.B2(n_267),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_258),
.A2(n_232),
.B1(n_242),
.B2(n_254),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_308),
.A2(n_320),
.B1(n_330),
.B2(n_291),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_241),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_309),
.B(n_321),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_234),
.B1(n_253),
.B2(n_241),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_313),
.B(n_316),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_257),
.A2(n_211),
.B1(n_240),
.B2(n_237),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_314),
.A2(n_328),
.B1(n_273),
.B2(n_274),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_258),
.A2(n_211),
.B1(n_224),
.B2(n_245),
.Y(n_320)
);

OAI32xp33_ASAP7_75t_L g321 ( 
.A1(n_260),
.A2(n_245),
.A3(n_214),
.B1(n_225),
.B2(n_227),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_323),
.B(n_285),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_281),
.A2(n_225),
.B(n_214),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_326),
.A2(n_329),
.B(n_287),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_291),
.A2(n_39),
.B1(n_32),
.B2(n_30),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_279),
.A2(n_47),
.B(n_1),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_277),
.A2(n_32),
.B1(n_30),
.B2(n_42),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_264),
.Y(n_333)
);

INVx13_ASAP7_75t_L g365 ( 
.A(n_333),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_334),
.A2(n_353),
.B1(n_314),
.B2(n_346),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_318),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_335),
.B(n_356),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_278),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_336),
.B(n_347),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_337),
.A2(n_317),
.B(n_362),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_272),
.C(n_276),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_339),
.B(n_342),
.Y(n_371)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_340),
.Y(n_366)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_297),
.Y(n_341)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_341),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_311),
.B(n_272),
.C(n_270),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_298),
.B(n_280),
.C(n_255),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_352),
.Y(n_372)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_344),
.Y(n_370)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_319),
.Y(n_345)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_345),
.Y(n_375)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_346),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_306),
.B(n_284),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_348),
.A2(n_322),
.B1(n_308),
.B2(n_320),
.Y(n_374)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_332),
.Y(n_349)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_349),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_282),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_350),
.B(n_351),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_305),
.B(n_263),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_298),
.B(n_261),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_322),
.A2(n_288),
.B1(n_259),
.B2(n_269),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_332),
.Y(n_354)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_354),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_305),
.B(n_290),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_302),
.Y(n_357)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_357),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_307),
.B(n_304),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_358),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_307),
.B(n_300),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_359),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_313),
.B(n_292),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_321),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_333),
.B(n_289),
.Y(n_361)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_361),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_317),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_317),
.Y(n_368)
);

FAx1_ASAP7_75t_SL g363 ( 
.A(n_310),
.B(n_265),
.CI(n_14),
.CON(n_363),
.SN(n_363)
);

NOR2x1_ASAP7_75t_L g382 ( 
.A(n_363),
.B(n_303),
.Y(n_382)
);

O2A1O1Ixp33_ASAP7_75t_L g377 ( 
.A1(n_364),
.A2(n_303),
.B(n_326),
.C(n_329),
.Y(n_377)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_368),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_369),
.Y(n_415)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_340),
.Y(n_373)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_373),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_374),
.A2(n_377),
.B1(n_334),
.B2(n_364),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_302),
.Y(n_378)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_379),
.B(n_355),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_380),
.A2(n_337),
.B1(n_365),
.B2(n_310),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_382),
.B(n_328),
.Y(n_413)
);

NOR4xp25_ASAP7_75t_L g385 ( 
.A(n_342),
.B(n_343),
.C(n_339),
.D(n_361),
.Y(n_385)
);

NAND3xp33_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_363),
.C(n_349),
.Y(n_405)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_365),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_391),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_338),
.B(n_309),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_393),
.B(n_352),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_390),
.A2(n_338),
.B1(n_348),
.B2(n_330),
.Y(n_394)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_394),
.Y(n_423)
);

MAJx2_ASAP7_75t_L g395 ( 
.A(n_371),
.B(n_355),
.C(n_360),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_398),
.Y(n_419)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_397),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_353),
.C(n_316),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_400),
.C(n_406),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_372),
.B(n_379),
.C(n_368),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_367),
.B(n_299),
.Y(n_401)
);

NAND3xp33_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_405),
.C(n_411),
.Y(n_432)
);

XNOR2x1_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_364),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_380),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_404),
.A2(n_381),
.B1(n_389),
.B2(n_393),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_388),
.B(n_325),
.C(n_344),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_381),
.A2(n_301),
.B1(n_341),
.B2(n_363),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_408),
.B(n_413),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_410),
.A2(n_391),
.B1(n_370),
.B2(n_384),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_376),
.B(n_325),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_324),
.C(n_327),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_414),
.C(n_370),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_389),
.B(n_324),
.C(n_327),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_378),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_416),
.B(n_383),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_404),
.A2(n_369),
.B(n_377),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_417),
.B(n_425),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_397),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_421),
.A2(n_428),
.B1(n_433),
.B2(n_409),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_422),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_399),
.A2(n_382),
.B(n_392),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_424),
.A2(n_431),
.B(n_12),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_426),
.A2(n_409),
.B1(n_268),
.B2(n_32),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_396),
.A2(n_384),
.B1(n_366),
.B2(n_387),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_373),
.C(n_375),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_429),
.B(n_434),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_386),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_430),
.B(n_407),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_396),
.A2(n_410),
.B(n_415),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_SL g433 ( 
.A1(n_402),
.A2(n_386),
.B1(n_375),
.B2(n_315),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_414),
.A2(n_315),
.B(n_285),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_429),
.B(n_395),
.C(n_398),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_438),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_439),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_418),
.B(n_406),
.C(n_412),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_407),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_444),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_441),
.Y(n_457)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_443),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_419),
.B(n_268),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_445),
.B(n_446),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_418),
.B(n_83),
.C(n_73),
.Y(n_446)
);

BUFx12f_ASAP7_75t_SL g447 ( 
.A(n_432),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g462 ( 
.A(n_447),
.Y(n_462)
);

XOR2x1_ASAP7_75t_SL g448 ( 
.A(n_431),
.B(n_16),
.Y(n_448)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_448),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_438),
.B(n_425),
.C(n_420),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_452),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_449),
.A2(n_423),
.B1(n_422),
.B2(n_435),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_437),
.A2(n_426),
.B1(n_427),
.B2(n_417),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_460),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_430),
.C(n_428),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_447),
.A2(n_42),
.B1(n_14),
.B2(n_13),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_463),
.B(n_448),
.C(n_450),
.Y(n_465)
);

AND2x4_ASAP7_75t_SL g464 ( 
.A(n_462),
.B(n_442),
.Y(n_464)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_464),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_468),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_436),
.C(n_439),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_466),
.B(n_469),
.C(n_456),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_451),
.A2(n_446),
.B(n_444),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_467),
.B(n_453),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_460),
.A2(n_14),
.B(n_13),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_459),
.B(n_13),
.C(n_12),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_47),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_473),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_461),
.B(n_0),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_474),
.B(n_477),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_472),
.B(n_456),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_479),
.A2(n_470),
.B1(n_452),
.B2(n_464),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_480),
.A2(n_483),
.B(n_475),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_476),
.A2(n_454),
.B(n_458),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_482),
.A2(n_478),
.B(n_42),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_478),
.A2(n_473),
.B(n_457),
.Y(n_483)
);

AOI322xp5_ASAP7_75t_L g486 ( 
.A1(n_484),
.A2(n_485),
.A3(n_481),
.B1(n_1),
.B2(n_2),
.C1(n_4),
.C2(n_0),
.Y(n_486)
);

OAI21x1_ASAP7_75t_SL g487 ( 
.A1(n_486),
.A2(n_1),
.B(n_2),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_487),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_488),
.B(n_9),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_489),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_490)
);

MAJx2_ASAP7_75t_L g491 ( 
.A(n_490),
.B(n_7),
.C(n_9),
.Y(n_491)
);


endmodule