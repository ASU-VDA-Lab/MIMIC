module fake_jpeg_4305_n_345 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_32),
.B1(n_21),
.B2(n_26),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_30),
.B1(n_32),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_48),
.A2(n_50),
.B1(n_53),
.B2(n_66),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_49),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_32),
.B1(n_24),
.B2(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_27),
.B1(n_20),
.B2(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_62),
.Y(n_82)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_17),
.B1(n_20),
.B2(n_39),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_71),
.B1(n_25),
.B2(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g87 ( 
.A(n_65),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_17),
.B1(n_25),
.B2(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_37),
.A2(n_22),
.B1(n_25),
.B2(n_29),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_42),
.C(n_35),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_46),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_75),
.A2(n_88),
.B1(n_91),
.B2(n_55),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_97),
.B(n_95),
.Y(n_119)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_86),
.Y(n_103)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_89),
.Y(n_109)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_54),
.A2(n_25),
.B1(n_13),
.B2(n_11),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_54),
.A2(n_14),
.B1(n_15),
.B2(n_12),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_94),
.Y(n_114)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_98),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_33),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_101),
.Y(n_140)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_105),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_71),
.B1(n_64),
.B2(n_51),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_94),
.B1(n_78),
.B2(n_96),
.Y(n_135)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_113),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_57),
.B(n_47),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_111),
.A2(n_118),
.B(n_119),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_62),
.Y(n_113)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_72),
.B1(n_86),
.B2(n_73),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_58),
.C(n_55),
.Y(n_118)
);

NAND2x1_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_90),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_46),
.B(n_33),
.Y(n_153)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_124),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_19),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_19),
.Y(n_125)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_99),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_138),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_133),
.B(n_141),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_90),
.B1(n_96),
.B2(n_79),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_135),
.B1(n_139),
.B2(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_64),
.B1(n_92),
.B2(n_72),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_110),
.B(n_83),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_59),
.B1(n_73),
.B2(n_58),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_152),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_83),
.B(n_19),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_145),
.A2(n_153),
.B(n_33),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_104),
.A2(n_93),
.B1(n_81),
.B2(n_98),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_148),
.A2(n_101),
.B1(n_100),
.B2(n_105),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_120),
.A2(n_70),
.B1(n_65),
.B2(n_56),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_155),
.B1(n_102),
.B2(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_109),
.A2(n_23),
.B1(n_29),
.B2(n_31),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_156),
.Y(n_160)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_158),
.B(n_168),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_113),
.C(n_118),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_159),
.B(n_163),
.C(n_132),
.Y(n_213)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_140),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_161),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_125),
.C(n_126),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_139),
.B1(n_135),
.B2(n_141),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_108),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_140),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_170),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_147),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_171),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_123),
.B1(n_107),
.B2(n_116),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_172),
.A2(n_176),
.B1(n_138),
.B2(n_148),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_19),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_150),
.A2(n_106),
.B1(n_112),
.B2(n_23),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_186),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_46),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_155),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_129),
.A2(n_112),
.B1(n_106),
.B2(n_19),
.Y(n_176)
);

AOI32xp33_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_67),
.A3(n_99),
.B1(n_115),
.B2(n_42),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_177),
.A2(n_179),
.B(n_185),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_18),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_182),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_131),
.A2(n_42),
.B(n_35),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_181),
.B(n_115),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_99),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_0),
.Y(n_184)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_142),
.A2(n_23),
.B1(n_29),
.B2(n_31),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_187),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_177),
.A2(n_131),
.B1(n_153),
.B2(n_151),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_190),
.A2(n_205),
.B(n_206),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_195),
.B1(n_169),
.B2(n_174),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_159),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_137),
.B1(n_136),
.B2(n_132),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_204),
.A2(n_172),
.B1(n_164),
.B2(n_170),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_146),
.Y(n_205)
);

AO22x1_ASAP7_75t_SL g206 ( 
.A1(n_184),
.A2(n_146),
.B1(n_31),
.B2(n_23),
.Y(n_206)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

AOI21x1_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_35),
.B(n_132),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_183),
.B(n_166),
.Y(n_235)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_160),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_215),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_163),
.C(n_182),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_165),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_214),
.Y(n_219)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_224),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_220),
.A2(n_190),
.B1(n_197),
.B2(n_211),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_232),
.C(n_237),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_222),
.B(n_225),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_173),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_227),
.B(n_228),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_236),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_202),
.A2(n_161),
.B1(n_167),
.B2(n_178),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_231),
.A2(n_234),
.B1(n_212),
.B2(n_196),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_181),
.C(n_168),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_158),
.B1(n_162),
.B2(n_180),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_235),
.A2(n_189),
.B(n_201),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_169),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_180),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_208),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_206),
.Y(n_240)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_187),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_242),
.C(n_192),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_115),
.C(n_31),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_244),
.A2(n_255),
.B1(n_257),
.B2(n_1),
.Y(n_283)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_249),
.A2(n_251),
.B(n_260),
.Y(n_276)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_254),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_266),
.Y(n_277)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_223),
.A2(n_191),
.B1(n_189),
.B2(n_211),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_218),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_223),
.A2(n_206),
.B1(n_208),
.B2(n_188),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_258),
.B(n_264),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_217),
.A2(n_214),
.B(n_215),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_209),
.C(n_198),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_263),
.C(n_265),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_0),
.C(n_1),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_1),
.C(n_2),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_220),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_271),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_246),
.A2(n_219),
.B1(n_226),
.B2(n_216),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_238),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_244),
.B(n_232),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_241),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_274),
.Y(n_292)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_282),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_217),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_280),
.C(n_281),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_243),
.B(n_240),
.C(n_228),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_233),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_8),
.Y(n_282)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_8),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_263),
.C(n_261),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_262),
.B(n_248),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_287),
.A2(n_300),
.B(n_15),
.Y(n_310)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_293),
.C(n_298),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_279),
.B(n_247),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_277),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_15),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_255),
.C(n_245),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_2),
.C(n_3),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_2),
.C(n_3),
.Y(n_312)
);

XOR2x2_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_9),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_284),
.Y(n_302)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_286),
.B(n_285),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_303),
.A2(n_312),
.B(n_315),
.Y(n_319)
);

OAI321xp33_ASAP7_75t_L g304 ( 
.A1(n_300),
.A2(n_269),
.A3(n_275),
.B1(n_271),
.B2(n_10),
.C(n_14),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_304),
.A2(n_308),
.B(n_310),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_294),
.A2(n_275),
.B1(n_9),
.B2(n_10),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_307),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_292),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

INVx11_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_313),
.A2(n_296),
.B1(n_4),
.B2(n_5),
.Y(n_325)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_298),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_314),
.A2(n_293),
.B1(n_299),
.B2(n_289),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_3),
.C(n_4),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_289),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_318),
.B(n_3),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_294),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_315),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_291),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_323),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_324),
.A2(n_311),
.B(n_306),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_327),
.A2(n_331),
.B(n_332),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_330),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_312),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_10),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_316),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_333),
.B(n_317),
.Y(n_336)
);

NOR2x1_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_325),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_335),
.A2(n_336),
.B(n_338),
.Y(n_340)
);

OAI321xp33_ASAP7_75t_L g338 ( 
.A1(n_332),
.A2(n_316),
.A3(n_319),
.B1(n_323),
.B2(n_12),
.C(n_4),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_334),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_339),
.A2(n_328),
.B(n_337),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_341),
.A2(n_340),
.B(n_5),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_342),
.Y(n_343)
);

NOR4xp25_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_344),
.B(n_6),
.Y(n_345)
);


endmodule