module fake_jpeg_13931_n_190 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_190);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_25),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_10),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_6),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_32),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_7),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_83),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_1),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_72),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

BUFx16f_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_70),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_98),
.C(n_104),
.Y(n_124)
);

OR2x2_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_70),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_57),
.B1(n_67),
.B2(n_74),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_76),
.B1(n_74),
.B2(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_75),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_55),
.C(n_77),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_59),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_SL g102 ( 
.A(n_90),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_102),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_60),
.C(n_62),
.Y(n_104)
);

INVxp67_ASAP7_75t_R g107 ( 
.A(n_106),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_109),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_68),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_112),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_120),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_64),
.B(n_61),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_123),
.B(n_69),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_63),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_92),
.B(n_65),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_117),
.B(n_20),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_96),
.B(n_73),
.Y(n_120)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_30),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_76),
.B1(n_56),
.B2(n_67),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_2),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_5),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_128),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_111),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_137),
.B1(n_147),
.B2(n_27),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_3),
.B(n_4),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_136),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_12),
.B1(n_14),
.B2(n_17),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_142),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_18),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_144),
.B(n_146),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_145),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_150),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_138),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_152),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_156),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_133),
.Y(n_156)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_135),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_160),
.B(n_135),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_163),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_37),
.A3(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_162),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_134),
.C(n_136),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_154),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_175),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_155),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_167),
.B(n_158),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_179),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_181),
.B(n_148),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_177),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_176),
.B(n_182),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_180),
.B(n_172),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_170),
.B(n_164),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_187),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_188),
.A2(n_170),
.B1(n_162),
.B2(n_165),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_168),
.Y(n_190)
);


endmodule