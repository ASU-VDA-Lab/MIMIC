module fake_jpeg_6646_n_176 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_26),
.B1(n_13),
.B2(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_26),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_50),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_46),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_31),
.B(n_22),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_28),
.A2(n_27),
.B1(n_15),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_23),
.B1(n_16),
.B2(n_21),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_24),
.Y(n_50)
);

CKINVDCx6p67_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_52),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_23),
.B1(n_16),
.B2(n_15),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_49),
.B1(n_61),
.B2(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_38),
.B(n_21),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_25),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_25),
.Y(n_83)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_68),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_51),
.C(n_42),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_75),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_52),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_70),
.A2(n_45),
.B(n_40),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_67),
.B(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_78),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_76),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_67),
.B(n_61),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_41),
.B1(n_51),
.B2(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_39),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NOR3xp33_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_40),
.C(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_14),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_69),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_41),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_92),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_70),
.A2(n_41),
.B(n_48),
.Y(n_92)
);

OAI211xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_96),
.B(n_81),
.C(n_77),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_74),
.A2(n_49),
.B1(n_66),
.B2(n_53),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_97),
.B(n_100),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_25),
.B(n_21),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_99),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_75),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_93),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_94),
.B(n_72),
.Y(n_104)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_76),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_64),
.B(n_17),
.Y(n_128)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_74),
.B1(n_83),
.B2(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

OAI321xp33_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_82),
.A3(n_21),
.B1(n_10),
.B2(n_12),
.C(n_11),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_98),
.Y(n_125)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_114),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_99),
.B(n_82),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_87),
.B(n_53),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_91),
.C(n_89),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_124),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_108),
.C(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_126),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_64),
.C(n_17),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_140)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_117),
.Y(n_135)
);

XNOR2x1_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_17),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_115),
.B(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_132),
.Y(n_149)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_1),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_122),
.A2(n_111),
.B1(n_107),
.B2(n_115),
.Y(n_134)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_105),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_141),
.B(n_1),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_140),
.A2(n_126),
.B(n_127),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_12),
.B1(n_2),
.B2(n_5),
.Y(n_142)
);

OA21x2_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_125),
.B(n_5),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_6),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_119),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_148),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_128),
.C(n_121),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_133),
.C(n_136),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_140),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_153),
.B(n_160),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_154),
.A2(n_151),
.B(n_148),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_150),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_143),
.A2(n_141),
.B1(n_142),
.B2(n_8),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_159),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_6),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_164),
.B(n_166),
.Y(n_170)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_163),
.B(n_157),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_144),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_170),
.B(n_165),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_153),
.B1(n_147),
.B2(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_169),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_157),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_173),
.C(n_7),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_169),
.A2(n_163),
.B(n_145),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_6),
.C(n_7),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);


endmodule