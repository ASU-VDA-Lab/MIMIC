module fake_jpeg_13190_n_525 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_525);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_361;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_51),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_21),
.B(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_21),
.B(n_7),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_54),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_7),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_60),
.Y(n_118)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_22),
.B(n_7),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_65),
.B(n_66),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_6),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_67),
.B(n_70),
.Y(n_126)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_32),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_22),
.B(n_14),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_71),
.B(n_73),
.Y(n_142)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_23),
.B(n_6),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

BUFx12f_ASAP7_75t_SL g75 ( 
.A(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_92),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_82),
.Y(n_111)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_24),
.B(n_44),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_66),
.A2(n_43),
.B1(n_34),
.B2(n_37),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_99),
.A2(n_139),
.B1(n_141),
.B2(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_54),
.B(n_42),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_134),
.B(n_148),
.Y(n_161)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_75),
.A2(n_40),
.B1(n_43),
.B2(n_34),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_45),
.A2(n_43),
.B1(n_37),
.B2(n_40),
.Y(n_141)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_57),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_48),
.A2(n_46),
.B1(n_50),
.B2(n_60),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_50),
.B(n_44),
.Y(n_148)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_68),
.A2(n_37),
.B1(n_28),
.B2(n_39),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_28),
.B1(n_38),
.B2(n_42),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_47),
.A2(n_37),
.B1(n_27),
.B2(n_15),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_15),
.B1(n_27),
.B2(n_24),
.Y(n_173)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_94),
.B1(n_90),
.B2(n_93),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_162),
.B1(n_183),
.B2(n_186),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_156),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_126),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_170),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_52),
.B1(n_55),
.B2(n_69),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_146),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_163),
.B(n_192),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_165),
.Y(n_236)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_166),
.Y(n_225)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_101),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_119),
.A2(n_85),
.B1(n_25),
.B2(n_20),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_199),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_187),
.Y(n_216)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_113),
.Y(n_174)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_174),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_103),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_193),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_25),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_184),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_99),
.A2(n_139),
.B1(n_128),
.B2(n_109),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_SL g213 ( 
.A1(n_181),
.A2(n_157),
.B(n_162),
.C(n_185),
.Y(n_213)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_124),
.B(n_20),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_104),
.A2(n_78),
.B(n_39),
.C(n_38),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_185),
.B(n_114),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_106),
.A2(n_87),
.B1(n_82),
.B2(n_89),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_123),
.A2(n_80),
.B1(n_41),
.B2(n_59),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_200),
.B1(n_111),
.B2(n_114),
.Y(n_205)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_97),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_63),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_121),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_125),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_195),
.Y(n_227)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_95),
.Y(n_196)
);

INVx13_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_201),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_132),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_153),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_119),
.A2(n_59),
.B1(n_63),
.B2(n_41),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_138),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_133),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_205),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_209),
.B(n_219),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_165),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_218),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_213),
.A2(n_193),
.B(n_175),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_111),
.C(n_147),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_201),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_161),
.B(n_122),
.Y(n_219)
);

CKINVDCx12_ASAP7_75t_R g221 ( 
.A(n_160),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_221),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_167),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_232),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_184),
.B(n_121),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_191),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_181),
.B(n_116),
.Y(n_232)
);

OR2x2_ASAP7_75t_SL g234 ( 
.A(n_181),
.B(n_169),
.Y(n_234)
);

NAND2xp67_ASAP7_75t_SL g238 ( 
.A(n_234),
.B(n_181),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_SL g270 ( 
.A1(n_238),
.A2(n_244),
.B(n_249),
.C(n_260),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_209),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_239),
.A2(n_250),
.B(n_254),
.Y(n_292)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_241),
.B(n_237),
.Y(n_301)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_242),
.Y(n_274)
);

AO22x2_ASAP7_75t_SL g244 ( 
.A1(n_213),
.A2(n_183),
.B1(n_168),
.B2(n_187),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_213),
.B1(n_204),
.B2(n_234),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_245),
.A2(n_236),
.B1(n_229),
.B2(n_98),
.Y(n_294)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_197),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_248),
.B(n_255),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_212),
.A2(n_191),
.B1(n_182),
.B2(n_175),
.Y(n_249)
);

NAND2xp33_ASAP7_75t_SL g250 ( 
.A(n_212),
.B(n_201),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_252),
.Y(n_286)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_253),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_189),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_223),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_210),
.Y(n_279)
);

OAI32xp33_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_180),
.A3(n_174),
.B1(n_194),
.B2(n_195),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_259),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_172),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_172),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_266),
.Y(n_296)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_227),
.Y(n_262)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_227),
.Y(n_263)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_263),
.Y(n_298)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_267),
.Y(n_293)
);

OA21x2_ASAP7_75t_L g266 ( 
.A1(n_216),
.A2(n_154),
.B(n_196),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_215),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_231),
.B(n_158),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_269),
.B(n_226),
.Y(n_281)
);

AO22x1_ASAP7_75t_SL g272 ( 
.A1(n_244),
.A2(n_245),
.B1(n_260),
.B2(n_238),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_272),
.B(n_281),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_248),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_280),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_243),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_277),
.B(n_285),
.Y(n_307)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_243),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_244),
.A2(n_268),
.B1(n_266),
.B2(n_259),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_282),
.A2(n_284),
.B1(n_294),
.B2(n_299),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_250),
.A2(n_212),
.B(n_211),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_283),
.A2(n_288),
.B(n_262),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_244),
.A2(n_204),
.B1(n_216),
.B2(n_205),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_269),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g288 ( 
.A(n_244),
.B(n_229),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_249),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_291),
.Y(n_319)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_241),
.B(n_230),
.C(n_214),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_295),
.B(n_297),
.C(n_242),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_215),
.C(n_236),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_266),
.A2(n_221),
.B1(n_203),
.B2(n_158),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_261),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_257),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_240),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_284),
.A2(n_239),
.B1(n_254),
.B2(n_247),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_302),
.A2(n_306),
.B1(n_308),
.B2(n_329),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g304 ( 
.A(n_297),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_304),
.B(n_322),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_282),
.A2(n_239),
.B1(n_247),
.B2(n_265),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_275),
.A2(n_265),
.B1(n_255),
.B2(n_256),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_309),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_288),
.A2(n_266),
.B1(n_252),
.B2(n_246),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_310),
.A2(n_314),
.B1(n_321),
.B2(n_294),
.Y(n_337)
);

AO21x1_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_264),
.B(n_263),
.Y(n_311)
);

AO21x1_ASAP7_75t_L g352 ( 
.A1(n_311),
.A2(n_312),
.B(n_333),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_313),
.B(n_316),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_288),
.A2(n_275),
.B1(n_296),
.B2(n_291),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_315),
.Y(n_358)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_317),
.Y(n_344)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_274),
.Y(n_318)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_318),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_320),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_288),
.A2(n_267),
.B1(n_258),
.B2(n_251),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_293),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_293),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_323),
.B(n_324),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_293),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_271),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_325),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_251),
.C(n_203),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_326),
.B(n_270),
.C(n_278),
.Y(n_346)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_327),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_296),
.A2(n_235),
.B1(n_208),
.B2(n_190),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_280),
.B(n_225),
.Y(n_331)
);

BUFx24_ASAP7_75t_SL g350 ( 
.A(n_331),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_276),
.B(n_225),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_332),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_290),
.B(n_298),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_298),
.Y(n_334)
);

INVxp33_ASAP7_75t_L g365 ( 
.A(n_334),
.Y(n_365)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_278),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_335),
.A2(n_289),
.B(n_286),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_337),
.A2(n_329),
.B1(n_335),
.B2(n_327),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_312),
.A2(n_292),
.B(n_283),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_339),
.A2(n_360),
.B(n_333),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_340),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_316),
.B(n_295),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_341),
.B(n_343),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_313),
.B(n_289),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_308),
.B(n_286),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_348),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_363),
.C(n_364),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_305),
.A2(n_299),
.B(n_270),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_311),
.B(n_272),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_306),
.B(n_272),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_353),
.B(n_356),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_302),
.B(n_270),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_330),
.A2(n_324),
.B(n_323),
.Y(n_360)
);

XNOR2x1_ASAP7_75t_L g362 ( 
.A(n_326),
.B(n_270),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_362),
.B(n_367),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_303),
.B(n_270),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_287),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_328),
.A2(n_287),
.B1(n_253),
.B2(n_235),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_366),
.A2(n_208),
.B1(n_176),
.B2(n_179),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_330),
.B(n_222),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_366),
.Y(n_368)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_368),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_338),
.B(n_307),
.Y(n_369)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_369),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_325),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_379),
.Y(n_399)
);

HAxp5_ASAP7_75t_SL g372 ( 
.A(n_339),
.B(n_319),
.CON(n_372),
.SN(n_372)
);

AND2x2_ASAP7_75t_SL g420 ( 
.A(n_372),
.B(n_387),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_349),
.A2(n_305),
.B1(n_314),
.B2(n_321),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_373),
.A2(n_393),
.B1(n_394),
.B2(n_397),
.Y(n_408)
);

XOR2x2_ASAP7_75t_L g422 ( 
.A(n_374),
.B(n_220),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_310),
.C(n_334),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_376),
.B(n_384),
.C(n_346),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_342),
.Y(n_377)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_377),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_378),
.A2(n_386),
.B1(n_390),
.B2(n_392),
.Y(n_407)
);

NAND3xp33_ASAP7_75t_L g379 ( 
.A(n_350),
.B(n_318),
.C(n_315),
.Y(n_379)
);

AOI21xp33_ASAP7_75t_L g380 ( 
.A1(n_336),
.A2(n_309),
.B(n_317),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_380),
.A2(n_391),
.B(n_352),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_253),
.Y(n_381)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_381),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_355),
.B(n_237),
.C(n_222),
.Y(n_384)
);

BUFx12f_ASAP7_75t_L g385 ( 
.A(n_365),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_385),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_361),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_354),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_353),
.B(n_220),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_388),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_364),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_363),
.A2(n_166),
.B(n_222),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_345),
.B(n_235),
.Y(n_392)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_344),
.Y(n_393)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_358),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_422),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_382),
.C(n_376),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_404),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_374),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_385),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_403),
.A2(n_224),
.B(n_120),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_370),
.B(n_341),
.C(n_362),
.Y(n_404)
);

MAJx2_ASAP7_75t_L g409 ( 
.A(n_396),
.B(n_337),
.C(n_352),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_409),
.B(n_417),
.C(n_419),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_375),
.A2(n_360),
.B1(n_359),
.B2(n_356),
.Y(n_410)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_410),
.Y(n_428)
);

FAx1_ASAP7_75t_SL g411 ( 
.A(n_389),
.B(n_343),
.CI(n_348),
.CON(n_411),
.SN(n_411)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_164),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_383),
.B(n_367),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_412),
.B(n_414),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_382),
.B(n_349),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_384),
.B(n_208),
.C(n_220),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_368),
.A2(n_123),
.B1(n_127),
.B2(n_143),
.Y(n_418)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_418),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_383),
.B(n_395),
.C(n_396),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_395),
.B(n_220),
.C(n_96),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_129),
.C(n_110),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_369),
.A2(n_127),
.B1(n_135),
.B2(n_96),
.Y(n_423)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_423),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_391),
.B(n_224),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_224),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_407),
.A2(n_394),
.B1(n_387),
.B2(n_378),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_426),
.A2(n_431),
.B1(n_439),
.B2(n_408),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_429),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_402),
.A2(n_387),
.B1(n_372),
.B2(n_381),
.Y(n_431)
);

FAx1_ASAP7_75t_SL g433 ( 
.A(n_404),
.B(n_385),
.CI(n_393),
.CON(n_433),
.SN(n_433)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_433),
.B(n_443),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_399),
.B(n_206),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_434),
.B(n_447),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_435),
.B(n_424),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_420),
.B(n_97),
.Y(n_436)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_436),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_437),
.A2(n_445),
.B(n_417),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_406),
.A2(n_129),
.B1(n_110),
.B2(n_105),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_398),
.Y(n_440)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_440),
.Y(n_459)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_405),
.Y(n_441)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_441),
.Y(n_462)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_413),
.Y(n_442)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_442),
.Y(n_464)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_416),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_422),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_415),
.B(n_120),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_400),
.B(n_105),
.C(n_140),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_448),
.B(n_401),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_455),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_450),
.A2(n_438),
.B1(n_451),
.B2(n_464),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_453),
.B(n_460),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_419),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_414),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_461),
.Y(n_474)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_458),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_430),
.B(n_409),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_444),
.B(n_421),
.C(n_420),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_463),
.B(n_465),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_444),
.B(n_420),
.C(n_412),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_430),
.B(n_428),
.C(n_425),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_466),
.B(n_429),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_436),
.A2(n_411),
.B1(n_8),
.B2(n_9),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_467),
.B(n_445),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_465),
.B(n_448),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_470),
.B(n_473),
.Y(n_492)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_472),
.Y(n_484)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_456),
.Y(n_475)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_475),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_433),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_476),
.B(n_14),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_477),
.Y(n_496)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_462),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_479),
.A2(n_482),
.B1(n_452),
.B2(n_435),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_466),
.A2(n_431),
.B(n_433),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_480),
.A2(n_463),
.B(n_467),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_426),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_481),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_494)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_459),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_460),
.B(n_436),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_483),
.B(n_478),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_485),
.B(n_487),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_432),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_489),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_478),
.B(n_455),
.Y(n_487)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_488),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_468),
.A2(n_446),
.B1(n_453),
.B2(n_439),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_491),
.A2(n_497),
.B(n_0),
.Y(n_507)
);

BUFx24_ASAP7_75t_SL g493 ( 
.A(n_471),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_493),
.B(n_474),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_494),
.B(n_477),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_495),
.A2(n_5),
.B(n_9),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_471),
.B(n_10),
.Y(n_497)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_499),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_501),
.A2(n_506),
.B(n_507),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_481),
.C(n_483),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_503),
.B(n_487),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_5),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_504),
.B(n_0),
.Y(n_509)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_505),
.Y(n_511)
);

A2O1A1Ixp33_ASAP7_75t_SL g506 ( 
.A1(n_496),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_506)
);

O2A1O1Ixp33_ASAP7_75t_SL g518 ( 
.A1(n_509),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_518)
);

AOI21xp33_ASAP7_75t_L g515 ( 
.A1(n_510),
.A2(n_502),
.B(n_491),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_484),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_512),
.B(n_513),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_498),
.B(n_488),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_515),
.B(n_517),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_506),
.C(n_1),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_518),
.B(n_511),
.C(n_509),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_519),
.B(n_516),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_521),
.B(n_520),
.C(n_514),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_2),
.C(n_3),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_2),
.B(n_4),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_4),
.B1(n_522),
.B2(n_210),
.Y(n_525)
);


endmodule