module fake_jpeg_9168_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_26),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_28),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_0),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_75),
.Y(n_83)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_1),
.B(n_2),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_59),
.B1(n_53),
.B2(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_70),
.B(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_81),
.Y(n_104)
);

INVx5_ASAP7_75t_SL g81 ( 
.A(n_73),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_79),
.A2(n_52),
.B1(n_49),
.B2(n_63),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_93),
.B1(n_85),
.B2(n_16),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_95),
.A2(n_97),
.B1(n_65),
.B2(n_51),
.Y(n_103)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_75),
.A2(n_64),
.B1(n_62),
.B2(n_50),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_112)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_90),
.C(n_98),
.Y(n_100)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_103),
.B1(n_106),
.B2(n_107),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_61),
.B1(n_55),
.B2(n_3),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_3),
.B1(n_4),
.B2(n_48),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_116),
.A2(n_115),
.B1(n_112),
.B2(n_114),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_119),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_104),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_118),
.C(n_116),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_109),
.C(n_108),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_124),
.A2(n_108),
.B(n_17),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_111),
.B1(n_113),
.B2(n_105),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_110),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_15),
.C(n_18),
.Y(n_128)
);

AO21x1_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_22),
.B(n_23),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_24),
.B(n_25),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_29),
.B(n_30),
.C(n_36),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_39),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_133),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_134),
.Y(n_135)
);


endmodule