module real_jpeg_4003_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_1),
.A2(n_83),
.B1(n_87),
.B2(n_88),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_1),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_1),
.A2(n_87),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_2),
.Y(n_86)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_2),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_3),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_3),
.B(n_157),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_3),
.A2(n_69),
.B1(n_144),
.B2(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_3),
.B(n_105),
.C(n_131),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_3),
.B(n_24),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_3),
.B(n_265),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_3),
.B(n_145),
.Y(n_293)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_4),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_4),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_4),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_5),
.A2(n_133),
.B1(n_137),
.B2(n_139),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_5),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_5),
.A2(n_44),
.B1(n_139),
.B2(n_230),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_5),
.A2(n_139),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_6),
.A2(n_100),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_6),
.Y(n_201)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_8),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_8),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_8),
.Y(n_162)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_8),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_8),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_8),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_9),
.A2(n_39),
.B1(n_44),
.B2(n_48),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_9),
.A2(n_48),
.B1(n_138),
.B2(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_9),
.A2(n_48),
.B1(n_285),
.B2(n_288),
.Y(n_284)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_10),
.Y(n_182)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_10),
.Y(n_213)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_12),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_12),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_12),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_12),
.Y(n_216)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_12),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_12),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_13),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_13),
.A2(n_54),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_13),
.A2(n_54),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_13),
.A2(n_54),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_14),
.A2(n_100),
.B1(n_104),
.B2(n_107),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_14),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_242),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_240),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_168),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_19),
.B(n_168),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_110),
.C(n_146),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_20),
.A2(n_21),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_67),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_22),
.B(n_68),
.C(n_81),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_38),
.B(n_49),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_23),
.A2(n_38),
.B1(n_57),
.B2(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_23),
.B(n_51),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_24),
.B(n_58),
.Y(n_57)
);

AO22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_32),
.B2(n_35),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g270 ( 
.A(n_29),
.Y(n_270)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_31),
.Y(n_136)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_31),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_31),
.Y(n_255)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_33),
.Y(n_236)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_37),
.Y(n_155)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_42),
.Y(n_148)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_43),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_43),
.Y(n_176)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_56),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_56),
.A2(n_313),
.B(n_316),
.Y(n_312)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_65),
.Y(n_58)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g158 ( 
.A(n_63),
.B(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_81),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_69),
.B(n_188),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_SL g218 ( 
.A1(n_69),
.A2(n_187),
.B(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_69),
.A2(n_193),
.B(n_263),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_SL g313 ( 
.A1(n_69),
.A2(n_314),
.B(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_71),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_72),
.B(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_75),
.B1(n_77),
.B2(n_79),
.Y(n_72)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_73),
.Y(n_184)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_73),
.Y(n_217)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_93),
.B1(n_99),
.B2(n_108),
.Y(n_81)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_82),
.Y(n_161)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_85),
.Y(n_203)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g279 ( 
.A(n_86),
.Y(n_279)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g262 ( 
.A(n_89),
.Y(n_262)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_93),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_93),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_93),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_99),
.Y(n_194)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_103),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_106),
.Y(n_287)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_110),
.B(n_146),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_132),
.B(n_140),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_111),
.A2(n_140),
.B(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_111),
.A2(n_132),
.B1(n_233),
.B2(n_269),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_112),
.B(n_141),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_123),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_117),
.B1(n_120),
.B2(n_122),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_SL g138 ( 
.A(n_122),
.Y(n_138)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_123),
.A2(n_238),
.B(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_126),
.B1(n_128),
.B2(n_130),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g289 ( 
.A(n_129),
.Y(n_289)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_143),
.Y(n_237)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_145),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_160),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_147),
.B(n_160),
.Y(n_317)
);

AOI32xp33_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.A3(n_153),
.B1(n_156),
.B2(n_158),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_152),
.Y(n_251)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_156),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B(n_163),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_163),
.A2(n_284),
.B(n_290),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_164),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_207),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_169)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_191),
.B2(n_192),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_177),
.A3(n_180),
.B1(n_183),
.B2(n_187),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_176),
.Y(n_231)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_176),
.Y(n_314)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_199),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_193),
.A2(n_259),
.B(n_263),
.Y(n_258)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_198),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_204),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_227),
.B2(n_239),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_218),
.B(n_221),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_211)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_227),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B(n_238),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AO21x1_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_319),
.B(n_324),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_305),
.B(n_318),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_273),
.B(n_304),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_257),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_246),
.B(n_257),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_252),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_247),
.A2(n_252),
.B1(n_253),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_247),
.Y(n_302)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

INVx3_ASAP7_75t_SL g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_266),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_267),
.C(n_272),
.Y(n_306)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_259),
.Y(n_298)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_271),
.B2(n_272),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_295),
.B(n_303),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_282),
.B(n_294),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_293),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_293),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_301),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_301),
.Y(n_303)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_307),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_317),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_311),
.C(n_317),
.Y(n_320)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_320),
.B(n_321),
.Y(n_324)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);


endmodule