module real_aes_5374_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_298;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_914;
wire n_203;
wire n_536;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_653;
wire n_155;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx1_ASAP7_75t_L g547 ( .A(n_0), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_1), .A2(n_13), .B1(n_121), .B2(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g591 ( .A(n_2), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g148 ( .A1(n_3), .A2(n_31), .B1(n_149), .B2(n_152), .Y(n_148) );
INVx1_ASAP7_75t_SL g645 ( .A(n_4), .Y(n_645) );
INVx1_ASAP7_75t_L g521 ( .A(n_5), .Y(n_521) );
INVx1_ASAP7_75t_L g876 ( .A(n_5), .Y(n_876) );
INVxp67_ASAP7_75t_L g893 ( .A(n_5), .Y(n_893) );
BUFx2_ASAP7_75t_L g915 ( .A(n_5), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_6), .A2(n_86), .B1(n_197), .B2(n_198), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_7), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_8), .B(n_143), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_9), .A2(n_33), .B1(n_118), .B2(n_120), .Y(n_117) );
INVx2_ASAP7_75t_L g228 ( .A(n_10), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_11), .A2(n_53), .B1(n_134), .B2(n_553), .Y(n_552) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_12), .A2(n_65), .B(n_139), .Y(n_138) );
OA21x2_ASAP7_75t_L g144 ( .A1(n_12), .A2(n_65), .B(n_139), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_14), .B(n_224), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_15), .A2(n_78), .B1(n_131), .B2(n_153), .Y(n_586) );
INVx2_ASAP7_75t_L g633 ( .A(n_16), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_17), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_SL g225 ( .A(n_18), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_19), .B(n_242), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_20), .A2(n_22), .B1(n_197), .B2(n_198), .Y(n_597) );
BUFx3_ASAP7_75t_L g895 ( .A(n_21), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_23), .A2(n_60), .B1(n_150), .B2(n_589), .Y(n_588) );
O2A1O1Ixp5_ASAP7_75t_L g629 ( .A1(n_24), .A2(n_128), .B(n_149), .C(n_630), .Y(n_629) );
O2A1O1Ixp5_ASAP7_75t_L g246 ( .A1(n_25), .A2(n_127), .B(n_247), .C(n_250), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_26), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_27), .B(n_158), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_28), .A2(n_79), .B1(n_221), .B2(n_254), .Y(n_558) );
INVx1_ASAP7_75t_L g525 ( .A(n_29), .Y(n_525) );
INVx1_ASAP7_75t_L g626 ( .A(n_30), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_32), .A2(n_100), .B1(n_907), .B2(n_916), .Y(n_99) );
AND2x2_ASAP7_75t_L g913 ( .A(n_34), .B(n_914), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_35), .B(n_235), .Y(n_543) );
INVx2_ASAP7_75t_L g631 ( .A(n_36), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_37), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g156 ( .A1(n_38), .A2(n_43), .B1(n_157), .B2(n_159), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_39), .A2(n_64), .B1(n_159), .B2(n_180), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_40), .B(n_153), .Y(n_233) );
INVx2_ASAP7_75t_L g173 ( .A(n_41), .Y(n_173) );
INVx2_ASAP7_75t_L g605 ( .A(n_42), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_44), .B(n_158), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_45), .B(n_137), .Y(n_203) );
INVx1_ASAP7_75t_SL g648 ( .A(n_46), .Y(n_648) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_47), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_48), .A2(n_124), .B(n_221), .C(n_222), .Y(n_220) );
INVx1_ASAP7_75t_L g306 ( .A(n_49), .Y(n_306) );
INVx1_ASAP7_75t_L g570 ( .A(n_50), .Y(n_570) );
INVx2_ASAP7_75t_L g257 ( .A(n_51), .Y(n_257) );
INVx1_ASAP7_75t_L g139 ( .A(n_52), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_54), .B(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g188 ( .A(n_54), .B(n_141), .Y(n_188) );
INVx2_ASAP7_75t_L g182 ( .A(n_55), .Y(n_182) );
INVx1_ASAP7_75t_L g651 ( .A(n_56), .Y(n_651) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_57), .Y(n_125) );
INVx1_ASAP7_75t_SL g251 ( .A(n_58), .Y(n_251) );
AOI221xp5_ASAP7_75t_L g102 ( .A1(n_59), .A2(n_103), .B1(n_104), .B2(n_878), .C(n_881), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_59), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_61), .B(n_610), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_62), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g898 ( .A1(n_63), .A2(n_899), .B1(n_900), .B2(n_901), .Y(n_898) );
CKINVDCx14_ASAP7_75t_R g899 ( .A(n_63), .Y(n_899) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_66), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g887 ( .A(n_67), .Y(n_887) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_68), .A2(n_124), .B(n_149), .C(n_185), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_69), .Y(n_624) );
OR2x6_ASAP7_75t_L g522 ( .A(n_70), .B(n_523), .Y(n_522) );
AND3x1_ASAP7_75t_L g912 ( .A(n_70), .B(n_913), .C(n_915), .Y(n_912) );
CKINVDCx16_ASAP7_75t_R g292 ( .A(n_71), .Y(n_292) );
INVx1_ASAP7_75t_L g302 ( .A(n_72), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_73), .B(n_154), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_74), .B(n_118), .Y(n_240) );
NOR2xp67_ASAP7_75t_L g216 ( .A(n_75), .B(n_217), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_76), .A2(n_177), .B(n_179), .C(n_183), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g282 ( .A1(n_76), .A2(n_177), .B(n_179), .C(n_183), .Y(n_282) );
INVx1_ASAP7_75t_L g524 ( .A(n_77), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g911 ( .A(n_77), .B(n_525), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_80), .A2(n_92), .B1(n_130), .B2(n_134), .Y(n_129) );
INVx1_ASAP7_75t_L g914 ( .A(n_81), .Y(n_914) );
BUFx5_ASAP7_75t_L g119 ( .A(n_82), .Y(n_119) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_82), .Y(n_122) );
INVx1_ASAP7_75t_L g133 ( .A(n_82), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_83), .B(n_297), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_84), .B(n_610), .Y(n_646) );
INVx2_ASAP7_75t_L g608 ( .A(n_85), .Y(n_608) );
INVx1_ASAP7_75t_L g613 ( .A(n_87), .Y(n_613) );
INVx2_ASAP7_75t_L g577 ( .A(n_88), .Y(n_577) );
INVx2_ASAP7_75t_SL g141 ( .A(n_89), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_90), .Y(n_882) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_91), .B(n_242), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_93), .B(n_144), .Y(n_303) );
INVx1_ASAP7_75t_SL g168 ( .A(n_94), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_95), .B(n_189), .Y(n_260) );
AND2x2_ASAP7_75t_L g142 ( .A(n_96), .B(n_143), .Y(n_142) );
INVx1_ASAP7_75t_SL g255 ( .A(n_97), .Y(n_255) );
AO22x2_ASAP7_75t_L g593 ( .A1(n_98), .A2(n_308), .B1(n_594), .B2(n_598), .Y(n_593) );
AO32x2_ASAP7_75t_L g666 ( .A1(n_98), .A2(n_194), .A3(n_309), .B1(n_594), .B2(n_667), .Y(n_666) );
AO21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_894), .B(n_896), .Y(n_100) );
NAND2xp5_ASAP7_75t_SL g101 ( .A(n_102), .B(n_886), .Y(n_101) );
OAI22x1_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_517), .B1(n_526), .B2(n_871), .Y(n_104) );
INVx1_ASAP7_75t_L g900 ( .A(n_105), .Y(n_900) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_106), .A2(n_527), .B1(n_872), .B2(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g901 ( .A(n_106), .Y(n_901) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_429), .Y(n_106) );
NAND3xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_349), .C(n_393), .Y(n_107) );
NOR3xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_319), .C(n_337), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_272), .Y(n_109) );
AOI22xp33_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_204), .B1(n_261), .B2(n_269), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g405 ( .A(n_112), .Y(n_405) );
OR2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_169), .Y(n_112) );
NOR2x1p5_ASAP7_75t_L g420 ( .A(n_113), .B(n_325), .Y(n_420) );
NAND2x1_ASAP7_75t_L g113 ( .A(n_114), .B(n_145), .Y(n_113) );
INVx2_ASAP7_75t_L g264 ( .A(n_114), .Y(n_264) );
INVx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g329 ( .A(n_115), .Y(n_329) );
AO31x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_126), .A3(n_135), .B(n_142), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_123), .Y(n_116) );
A2O1A1Ixp33_ASAP7_75t_L g647 ( .A1(n_118), .A2(n_124), .B(n_648), .C(n_649), .Y(n_647) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g134 ( .A(n_119), .Y(n_134) );
INVx2_ASAP7_75t_L g158 ( .A(n_119), .Y(n_158) );
INVx1_ASAP7_75t_L g178 ( .A(n_119), .Y(n_178) );
INVx2_ASAP7_75t_L g197 ( .A(n_119), .Y(n_197) );
NAND2xp33_ASAP7_75t_L g214 ( .A(n_119), .B(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g627 ( .A(n_120), .Y(n_627) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVxp67_ASAP7_75t_SL g221 ( .A(n_121), .Y(n_221) );
INVx1_ASAP7_75t_L g256 ( .A(n_121), .Y(n_256) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx3_ASAP7_75t_L g154 ( .A(n_122), .Y(n_154) );
INVx2_ASAP7_75t_L g181 ( .A(n_122), .Y(n_181) );
INVx6_ASAP7_75t_L g224 ( .A(n_122), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_123), .A2(n_156), .B(n_160), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_123), .B(n_187), .Y(n_567) );
NOR3xp33_ASAP7_75t_L g569 ( .A(n_123), .B(n_187), .C(n_570), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_123), .A2(n_586), .B1(n_587), .B2(n_588), .Y(n_585) );
INVx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g603 ( .A1(n_124), .A2(n_604), .B(n_605), .C(n_606), .Y(n_603) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_125), .Y(n_128) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_125), .Y(n_183) );
INVxp67_ASAP7_75t_L g200 ( .A(n_125), .Y(n_200) );
INVx4_ASAP7_75t_L g236 ( .A(n_125), .Y(n_236) );
INVx1_ASAP7_75t_L g560 ( .A(n_125), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_127), .B(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_127), .B(n_187), .Y(n_572) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_128), .A2(n_539), .B(n_541), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_128), .A2(n_218), .B1(n_595), .B2(n_597), .Y(n_594) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g159 ( .A(n_132), .Y(n_159) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g151 ( .A(n_133), .Y(n_151) );
INVx2_ASAP7_75t_L g300 ( .A(n_134), .Y(n_300) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_136), .B(n_194), .Y(n_279) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_136), .A2(n_563), .B(n_576), .Y(n_562) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_137), .B(n_259), .Y(n_258) );
BUFx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx4_ASAP7_75t_L g163 ( .A(n_138), .Y(n_163) );
INVx2_ASAP7_75t_L g227 ( .A(n_138), .Y(n_227) );
INVx3_ASAP7_75t_L g165 ( .A(n_140), .Y(n_165) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_140), .Y(n_194) );
INVx1_ASAP7_75t_L g259 ( .A(n_140), .Y(n_259) );
INVx3_ASAP7_75t_L g549 ( .A(n_140), .Y(n_549) );
AND2x2_ASAP7_75t_L g584 ( .A(n_140), .B(n_210), .Y(n_584) );
AND2x2_ASAP7_75t_L g598 ( .A(n_140), .B(n_599), .Y(n_598) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g167 ( .A(n_144), .Y(n_167) );
INVx1_ASAP7_75t_L g174 ( .A(n_144), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_144), .B(n_549), .Y(n_548) );
NOR2xp67_ASAP7_75t_L g555 ( .A(n_144), .B(n_549), .Y(n_555) );
INVx1_ASAP7_75t_L g578 ( .A(n_144), .Y(n_578) );
INVx1_ASAP7_75t_L g599 ( .A(n_144), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_144), .B(n_549), .Y(n_611) );
INVx1_ASAP7_75t_L g614 ( .A(n_144), .Y(n_614) );
NOR2x1_ASAP7_75t_L g330 ( .A(n_145), .B(n_278), .Y(n_330) );
INVx1_ASAP7_75t_L g380 ( .A(n_145), .Y(n_380) );
AND2x2_ASAP7_75t_L g440 ( .A(n_145), .B(n_266), .Y(n_440) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g277 ( .A(n_146), .Y(n_277) );
AOI21x1_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_155), .B(n_166), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_149), .B(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g610 ( .A(n_151), .Y(n_610) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g198 ( .A(n_154), .Y(n_198) );
INVx1_ASAP7_75t_L g217 ( .A(n_154), .Y(n_217) );
INVx1_ASAP7_75t_L g540 ( .A(n_154), .Y(n_540) );
INVx1_ASAP7_75t_L g553 ( .A(n_154), .Y(n_553) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp67_ASAP7_75t_L g565 ( .A(n_159), .B(n_566), .Y(n_565) );
A2O1A1Ixp33_ASAP7_75t_L g607 ( .A1(n_159), .A2(n_183), .B(n_608), .C(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_164), .Y(n_160) );
AOI21x1_ASAP7_75t_L g266 ( .A1(n_161), .A2(n_267), .B(n_268), .Y(n_266) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g211 ( .A(n_163), .Y(n_211) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_164), .A2(n_232), .B(n_237), .Y(n_231) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_165), .A2(n_303), .B(n_308), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx1_ASAP7_75t_L g189 ( .A(n_167), .Y(n_189) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g397 ( .A(n_170), .B(n_328), .Y(n_397) );
NOR2x1_ASAP7_75t_L g170 ( .A(n_171), .B(n_190), .Y(n_170) );
AND2x2_ASAP7_75t_L g353 ( .A(n_171), .B(n_329), .Y(n_353) );
INVx1_ASAP7_75t_L g419 ( .A(n_171), .Y(n_419) );
AND2x4_ASAP7_75t_L g427 ( .A(n_171), .B(n_264), .Y(n_427) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_171), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_171), .B(n_482), .Y(n_481) );
OR2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_175), .Y(n_171) );
INVxp67_ASAP7_75t_SL g284 ( .A(n_172), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
INVx1_ASAP7_75t_L g192 ( .A(n_174), .Y(n_192) );
NOR4xp25_ASAP7_75t_L g175 ( .A(n_176), .B(n_184), .C(n_187), .D(n_189), .Y(n_175) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g544 ( .A(n_178), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_180), .B(n_182), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_180), .B(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g254 ( .A(n_180), .Y(n_254) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g297 ( .A(n_181), .Y(n_297) );
INVx2_ASAP7_75t_SL g202 ( .A(n_183), .Y(n_202) );
INVx1_ASAP7_75t_L g218 ( .A(n_183), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_183), .B(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_183), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_183), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g587 ( .A(n_183), .Y(n_587) );
A2O1A1Ixp33_ASAP7_75t_L g643 ( .A1(n_183), .A2(n_644), .B(n_645), .C(n_646), .Y(n_643) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_184), .Y(n_283) );
NOR2x1_ASAP7_75t_SL g208 ( .A(n_187), .B(n_209), .Y(n_208) );
AOI221x1_ASAP7_75t_L g620 ( .A1(n_187), .A2(n_621), .B1(n_623), .B2(n_625), .C(n_627), .Y(n_620) );
INVx4_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_191), .Y(n_325) );
AND2x2_ASAP7_75t_L g348 ( .A(n_191), .B(n_276), .Y(n_348) );
INVx1_ASAP7_75t_L g476 ( .A(n_191), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_191), .B(n_329), .Y(n_479) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_203), .Y(n_191) );
OAI21x1_ASAP7_75t_L g230 ( .A1(n_192), .A2(n_231), .B(n_241), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_195), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_199), .B1(n_201), .B2(n_202), .Y(n_195) );
OAI22xp33_ASAP7_75t_L g573 ( .A1(n_197), .A2(n_249), .B1(n_574), .B2(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g644 ( .A(n_198), .Y(n_644) );
OAI21xp5_ASAP7_75t_SL g252 ( .A1(n_199), .A2(n_253), .B(n_258), .Y(n_252) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g268 ( .A(n_203), .Y(n_268) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_229), .Y(n_204) );
OR2x6_ASAP7_75t_L g335 ( .A(n_205), .B(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g447 ( .A(n_205), .B(n_357), .Y(n_447) );
INVx2_ASAP7_75t_SL g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g388 ( .A(n_206), .B(n_389), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_206), .B(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g436 ( .A(n_206), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g270 ( .A(n_207), .Y(n_270) );
OR2x2_ASAP7_75t_L g288 ( .A(n_207), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g343 ( .A(n_207), .B(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g362 ( .A(n_207), .B(n_289), .Y(n_362) );
AND2x2_ASAP7_75t_L g412 ( .A(n_207), .B(n_344), .Y(n_412) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_207), .Y(n_490) );
AO31x2_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_212), .A3(n_219), .B(n_226), .Y(n_207) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_211), .B(n_549), .Y(n_642) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_216), .B(n_218), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_218), .A2(n_238), .B(n_240), .Y(n_237) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_225), .Y(n_222) );
INVx1_ASAP7_75t_L g622 ( .A(n_223), .Y(n_622) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g239 ( .A(n_224), .Y(n_239) );
INVx2_ASAP7_75t_L g249 ( .A(n_224), .Y(n_249) );
INVx1_ASAP7_75t_L g295 ( .A(n_224), .Y(n_295) );
INVx1_ASAP7_75t_L g589 ( .A(n_224), .Y(n_589) );
INVx2_ASAP7_75t_SL g596 ( .A(n_224), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
INVx3_ASAP7_75t_L g242 ( .A(n_227), .Y(n_242) );
BUFx3_ASAP7_75t_L g309 ( .A(n_227), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_227), .B(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_227), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_243), .Y(n_229) );
AND2x2_ASAP7_75t_L g271 ( .A(n_230), .B(n_244), .Y(n_271) );
OR2x2_ASAP7_75t_L g395 ( .A(n_230), .B(n_343), .Y(n_395) );
AND2x2_ASAP7_75t_L g437 ( .A(n_230), .B(n_290), .Y(n_437) );
OAI21x1_ASAP7_75t_L g313 ( .A1(n_231), .A2(n_241), .B(n_308), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_235), .Y(n_232) );
AND2x2_ASAP7_75t_L g623 ( .A(n_235), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g625 ( .A(n_235), .B(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
O2A1O1Ixp5_ASAP7_75t_SL g291 ( .A1(n_236), .A2(n_292), .B(n_293), .C(n_296), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_236), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g311 ( .A(n_243), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g487 ( .A(n_243), .B(n_270), .Y(n_487) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_244), .B(n_366), .Y(n_365) );
INVx3_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g318 ( .A(n_245), .Y(n_318) );
INVx1_ASAP7_75t_L g376 ( .A(n_245), .Y(n_376) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_252), .B(n_260), .Y(n_245) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_249), .B(n_546), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B1(n_256), .B2(n_257), .Y(n_253) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g498 ( .A(n_262), .B(n_330), .Y(n_498) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
BUFx2_ASAP7_75t_SL g274 ( .A(n_264), .Y(n_274) );
INVx1_ASAP7_75t_L g341 ( .A(n_264), .Y(n_341) );
AND2x2_ASAP7_75t_L g381 ( .A(n_264), .B(n_278), .Y(n_381) );
AND2x2_ASAP7_75t_L g403 ( .A(n_265), .B(n_392), .Y(n_403) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g383 ( .A(n_266), .B(n_276), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_269), .B(n_422), .Y(n_421) );
INVxp33_ASAP7_75t_L g428 ( .A(n_269), .Y(n_428) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx1_ASAP7_75t_L g366 ( .A(n_270), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_270), .Y(n_369) );
OR2x2_ASAP7_75t_L g448 ( .A(n_270), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g497 ( .A(n_270), .B(n_316), .Y(n_497) );
INVx1_ASAP7_75t_L g389 ( .A(n_271), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_285), .Y(n_272) );
INVx1_ASAP7_75t_L g358 ( .A(n_273), .Y(n_358) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND2x1p5_ASAP7_75t_L g372 ( .A(n_275), .B(n_325), .Y(n_372) );
INVx3_ASAP7_75t_L g474 ( .A(n_275), .Y(n_474) );
AND2x4_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g392 ( .A(n_277), .Y(n_392) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_278), .Y(n_515) );
OA21x2_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_280), .B(n_284), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OAI21xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_310), .B(n_314), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g463 ( .A(n_288), .Y(n_463) );
OR2x2_ASAP7_75t_L g494 ( .A(n_288), .B(n_466), .Y(n_494) );
AND2x2_ASAP7_75t_L g317 ( .A(n_289), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_289), .B(n_316), .Y(n_357) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g450 ( .A(n_290), .B(n_312), .Y(n_450) );
OAI21x1_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_298), .B(n_307), .Y(n_290) );
OAI21xp5_ASAP7_75t_L g344 ( .A1(n_291), .A2(n_298), .B(n_307), .Y(n_344) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_294), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g568 ( .A(n_297), .Y(n_568) );
NAND3x1_ASAP7_75t_L g298 ( .A(n_299), .B(n_303), .C(n_304), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AO31x2_ASAP7_75t_L g619 ( .A1(n_309), .A2(n_620), .A3(n_628), .B(n_632), .Y(n_619) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g387 ( .A(n_311), .B(n_362), .Y(n_387) );
INVxp67_ASAP7_75t_L g400 ( .A(n_311), .Y(n_400) );
INVx2_ASAP7_75t_L g316 ( .A(n_312), .Y(n_316) );
AND2x2_ASAP7_75t_L g370 ( .A(n_312), .B(n_318), .Y(n_370) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g406 ( .A(n_314), .Y(n_406) );
NAND2x1p5_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx2_ASAP7_75t_L g416 ( .A(n_315), .Y(n_416) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_SL g336 ( .A(n_316), .Y(n_336) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_316), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_317), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g384 ( .A(n_317), .Y(n_384) );
INVx2_ASAP7_75t_SL g334 ( .A(n_318), .Y(n_334) );
BUFx2_ASAP7_75t_L g439 ( .A(n_318), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_331), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_326), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_324), .B(n_328), .Y(n_408) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g471 ( .A(n_325), .Y(n_471) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
NOR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g342 ( .A(n_334), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g411 ( .A(n_334), .Y(n_411) );
AND2x2_ASAP7_75t_L g491 ( .A(n_334), .B(n_450), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_334), .B(n_412), .Y(n_495) );
NOR3xp33_ASAP7_75t_L g514 ( .A(n_334), .B(n_340), .C(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g453 ( .A(n_335), .B(n_399), .Y(n_453) );
INVx1_ASAP7_75t_L g361 ( .A(n_336), .Y(n_361) );
O2A1O1Ixp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_342), .B(n_345), .C(n_347), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2x1p5_ASAP7_75t_L g457 ( .A(n_340), .B(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g382 ( .A(n_341), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g402 ( .A(n_341), .B(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g425 ( .A(n_343), .B(n_411), .Y(n_425) );
INVx1_ASAP7_75t_L g503 ( .A(n_343), .Y(n_503) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_344), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g485 ( .A1(n_347), .A2(n_457), .B1(n_486), .B2(n_488), .C(n_492), .Y(n_485) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g352 ( .A(n_348), .B(n_353), .Y(n_352) );
NOR4xp25_ASAP7_75t_L g349 ( .A(n_350), .B(n_363), .C(n_373), .D(n_385), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_354), .B1(n_358), .B2(n_359), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_351), .A2(n_364), .B1(n_367), .B2(n_371), .Y(n_363) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AOI21xp33_ASAP7_75t_SL g432 ( .A1(n_352), .A2(n_433), .B(n_434), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_353), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g409 ( .A(n_353), .Y(n_409) );
AND2x2_ASAP7_75t_L g470 ( .A(n_353), .B(n_471), .Y(n_470) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g465 ( .A(n_356), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI211xp5_ASAP7_75t_L g467 ( .A1(n_359), .A2(n_468), .B(n_469), .C(n_472), .Y(n_467) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_362), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g443 ( .A(n_362), .B(n_416), .Y(n_443) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g483 ( .A(n_369), .B(n_437), .Y(n_483) );
INVx1_ASAP7_75t_L g508 ( .A(n_370), .Y(n_508) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g458 ( .A(n_372), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_377), .B1(n_382), .B2(n_384), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_375), .B(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_R g466 ( .A(n_376), .Y(n_466) );
OAI22xp33_ASAP7_75t_L g424 ( .A1(n_377), .A2(n_425), .B1(n_426), .B2(n_428), .Y(n_424) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
NOR2xp33_ASAP7_75t_SL g516 ( .A(n_379), .B(n_475), .Y(n_516) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g510 ( .A(n_380), .B(n_397), .Y(n_510) );
AND2x4_ASAP7_75t_L g455 ( .A(n_381), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g500 ( .A(n_382), .Y(n_500) );
INVx2_ASAP7_75t_L g456 ( .A(n_383), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_388), .B(n_390), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_388), .A2(n_453), .B1(n_454), .B2(n_457), .C(n_459), .Y(n_452) );
AND2x2_ASAP7_75t_L g464 ( .A(n_391), .B(n_419), .Y(n_464) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_392), .Y(n_445) );
INVx1_ASAP7_75t_L g482 ( .A(n_392), .Y(n_482) );
NOR3xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_413), .C(n_424), .Y(n_393) );
OAI221xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_398), .B2(n_401), .C(n_404), .Y(n_394) );
INVx1_ASAP7_75t_L g499 ( .A(n_395), .Y(n_499) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_399), .A2(n_510), .B1(n_511), .B2(n_512), .Y(n_509) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_403), .B(n_418), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B1(n_407), .B2(n_410), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_414), .B(n_421), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .Y(n_414) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_420), .Y(n_460) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g433 ( .A(n_425), .Y(n_433) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g444 ( .A(n_427), .B(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g451 ( .A(n_427), .B(n_440), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_484), .Y(n_429) );
NOR3xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_452), .C(n_467), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_442), .Y(n_431) );
NOR3xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_438), .C(n_441), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI21xp33_ASAP7_75t_L g469 ( .A1(n_436), .A2(n_444), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g511 ( .A(n_437), .B(n_466), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g462 ( .A(n_439), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_446), .B2(n_451), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_455), .A2(n_503), .B1(n_504), .B2(n_507), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_461), .B1(n_464), .B2(n_465), .Y(n_459) );
INVx1_ASAP7_75t_L g468 ( .A(n_460), .Y(n_468) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
OAI21xp5_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_477), .B(n_483), .Y(n_472) );
NOR2x1_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_479), .B(n_481), .Y(n_506) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_501), .Y(n_484) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
AOI22xp33_ASAP7_75t_SL g492 ( .A1(n_493), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_492) );
NAND3xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .C(n_496), .Y(n_493) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_509), .Y(n_501) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_516), .Y(n_513) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx8_ASAP7_75t_L g880 ( .A(n_520), .Y(n_880) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
OR2x6_ASAP7_75t_L g885 ( .A(n_521), .B(n_522), .Y(n_885) );
INVx8_ASAP7_75t_L g877 ( .A(n_522), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVxp67_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
NOR2x1p5_ASAP7_75t_L g528 ( .A(n_529), .B(n_763), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_731), .Y(n_529) );
NOR4xp25_ASAP7_75t_L g530 ( .A(n_531), .B(n_672), .C(n_698), .D(n_717), .Y(n_530) );
OAI211xp5_ASAP7_75t_SL g531 ( .A1(n_532), .A2(n_579), .B(n_615), .C(n_660), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OAI21xp5_ASAP7_75t_L g729 ( .A1(n_533), .A2(n_654), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_561), .Y(n_533) );
AND2x2_ASAP7_75t_L g775 ( .A(n_534), .B(n_680), .Y(n_775) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_550), .Y(n_534) );
AND2x2_ASAP7_75t_L g639 ( .A(n_535), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g656 ( .A(n_535), .Y(n_656) );
INVx1_ASAP7_75t_L g707 ( .A(n_535), .Y(n_707) );
INVx2_ASAP7_75t_L g735 ( .A(n_535), .Y(n_735) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_535), .Y(n_866) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_542), .B(n_548), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B(n_545), .Y(n_542) );
INVx2_ASAP7_75t_L g637 ( .A(n_550), .Y(n_637) );
INVx1_ASAP7_75t_L g693 ( .A(n_550), .Y(n_693) );
AND2x2_ASAP7_75t_L g734 ( .A(n_550), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g816 ( .A(n_550), .Y(n_816) );
NAND2x1p5_ASAP7_75t_L g550 ( .A(n_551), .B(n_557), .Y(n_550) );
AND2x2_ASAP7_75t_SL g657 ( .A(n_551), .B(n_557), .Y(n_657) );
OA21x2_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_554), .B(n_556), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_555), .B(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx2_ASAP7_75t_L g736 ( .A(n_561), .Y(n_736) );
BUFx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g638 ( .A(n_562), .Y(n_638) );
OR2x2_ASAP7_75t_L g659 ( .A(n_562), .B(n_641), .Y(n_659) );
AND2x2_ASAP7_75t_L g862 ( .A(n_562), .B(n_702), .Y(n_862) );
AO21x2_ASAP7_75t_L g670 ( .A1(n_563), .A2(n_576), .B(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_571), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_567), .B1(n_568), .B2(n_569), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_L g667 ( .A(n_578), .Y(n_667) );
INVxp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_592), .Y(n_580) );
INVx4_ASAP7_75t_L g634 ( .A(n_581), .Y(n_634) );
INVx2_ASAP7_75t_L g677 ( .A(n_581), .Y(n_677) );
AND2x2_ASAP7_75t_L g694 ( .A(n_581), .B(n_695), .Y(n_694) );
BUFx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g665 ( .A(n_582), .Y(n_665) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g653 ( .A(n_583), .Y(n_653) );
INVx1_ASAP7_75t_L g690 ( .A(n_583), .Y(n_690) );
AOI21x1_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B(n_590), .Y(n_583) );
INVx1_ASAP7_75t_L g604 ( .A(n_589), .Y(n_604) );
AND2x4_ASAP7_75t_L g741 ( .A(n_592), .B(n_713), .Y(n_741) );
AND2x4_ASAP7_75t_L g756 ( .A(n_592), .B(n_757), .Y(n_756) );
AND2x4_ASAP7_75t_L g592 ( .A(n_593), .B(n_600), .Y(n_592) );
AND2x2_ASAP7_75t_L g652 ( .A(n_593), .B(n_653), .Y(n_652) );
AND2x4_ASAP7_75t_L g683 ( .A(n_593), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g716 ( .A(n_593), .Y(n_716) );
INVx1_ASAP7_75t_L g813 ( .A(n_593), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_596), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g689 ( .A(n_600), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g695 ( .A(n_600), .B(n_619), .Y(n_695) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g618 ( .A(n_601), .B(n_619), .Y(n_618) );
AND2x4_ASAP7_75t_L g675 ( .A(n_601), .B(n_676), .Y(n_675) );
BUFx3_ASAP7_75t_L g684 ( .A(n_601), .Y(n_684) );
INVx1_ASAP7_75t_L g715 ( .A(n_601), .Y(n_715) );
AND2x4_ASAP7_75t_L g789 ( .A(n_601), .B(n_790), .Y(n_789) );
INVx3_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AO31x2_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_607), .A3(n_611), .B(n_612), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
NOR2xp33_ASAP7_75t_SL g650 ( .A(n_614), .B(n_651), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_635), .B1(n_652), .B2(n_654), .Y(n_615) );
INVx3_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2x1p5_ASAP7_75t_L g617 ( .A(n_618), .B(n_634), .Y(n_617) );
AND2x2_ASAP7_75t_L g727 ( .A(n_618), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g857 ( .A(n_618), .B(n_813), .Y(n_857) );
INVx2_ASAP7_75t_L g663 ( .A(n_619), .Y(n_663) );
OR2x2_ASAP7_75t_L g758 ( .A(n_619), .B(n_653), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_619), .B(n_653), .Y(n_761) );
INVx1_ASAP7_75t_L g790 ( .A(n_619), .Y(n_790) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_639), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
AND2x2_ASAP7_75t_L g669 ( .A(n_637), .B(n_670), .Y(n_669) );
BUFx2_ASAP7_75t_L g681 ( .A(n_637), .Y(n_681) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_637), .Y(n_869) );
OR2x2_ASAP7_75t_L g706 ( .A(n_638), .B(n_707), .Y(n_706) );
AND2x4_ASAP7_75t_L g724 ( .A(n_638), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g668 ( .A(n_639), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g711 ( .A(n_639), .B(n_693), .Y(n_711) );
INVx1_ASAP7_75t_L g725 ( .A(n_640), .Y(n_725) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g680 ( .A(n_641), .B(n_670), .Y(n_680) );
INVx2_ASAP7_75t_L g702 ( .A(n_641), .Y(n_702) );
INVx1_ASAP7_75t_L g720 ( .A(n_641), .Y(n_720) );
INVx1_ASAP7_75t_L g818 ( .A(n_641), .Y(n_818) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_641), .Y(n_822) );
AO31x2_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .A3(n_647), .B(n_650), .Y(n_641) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_653), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_654), .A2(n_741), .B1(n_743), .B2(n_744), .Y(n_742) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_658), .Y(n_654) );
AND2x2_ASAP7_75t_L g751 ( .A(n_655), .B(n_724), .Y(n_751) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
AND2x2_ASAP7_75t_L g687 ( .A(n_656), .B(n_657), .Y(n_687) );
INVx1_ASAP7_75t_L g810 ( .A(n_656), .Y(n_810) );
AOI32xp33_ASAP7_75t_L g699 ( .A1(n_657), .A2(n_683), .A3(n_700), .B1(n_704), .B2(n_705), .Y(n_699) );
INVx2_ASAP7_75t_L g850 ( .A(n_657), .Y(n_850) );
INVx1_ASAP7_75t_L g697 ( .A(n_658), .Y(n_697) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_659), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_668), .Y(n_660) );
AND2x4_ASAP7_75t_SL g661 ( .A(n_662), .B(n_664), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
BUFx3_ASAP7_75t_L g713 ( .A(n_663), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_663), .B(n_676), .Y(n_749) );
AND2x2_ASAP7_75t_L g769 ( .A(n_663), .B(n_690), .Y(n_769) );
INVx2_ASAP7_75t_SL g781 ( .A(n_663), .Y(n_781) );
INVx1_ASAP7_75t_L g787 ( .A(n_664), .Y(n_787) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_665), .B(n_676), .Y(n_835) );
INVx2_ASAP7_75t_L g676 ( .A(n_666), .Y(n_676) );
BUFx8_ASAP7_75t_L g728 ( .A(n_666), .Y(n_728) );
INVxp67_ASAP7_75t_L g671 ( .A(n_667), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_668), .B(n_804), .Y(n_803) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_669), .B(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g746 ( .A(n_670), .B(n_735), .Y(n_746) );
AND2x2_ASAP7_75t_L g819 ( .A(n_670), .B(n_707), .Y(n_819) );
AND2x2_ASAP7_75t_L g849 ( .A(n_670), .B(n_850), .Y(n_849) );
OAI221xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_678), .B1(n_682), .B2(n_686), .C(n_688), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
INVx2_ASAP7_75t_L g779 ( .A(n_675), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_676), .B(n_781), .Y(n_780) );
AND2x2_ASAP7_75t_L g777 ( .A(n_677), .B(n_683), .Y(n_777) );
NOR2x1_ASAP7_75t_L g778 ( .A(n_677), .B(n_779), .Y(n_778) );
OAI21xp33_ASAP7_75t_SL g739 ( .A1(n_678), .A2(n_740), .B(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
AND2x2_ASAP7_75t_L g691 ( .A(n_680), .B(n_692), .Y(n_691) );
INVxp67_ASAP7_75t_L g784 ( .A(n_681), .Y(n_784) );
AND2x2_ASAP7_75t_L g802 ( .A(n_681), .B(n_724), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_685), .Y(n_682) );
INVx2_ASAP7_75t_SL g772 ( .A(n_684), .Y(n_772) );
OR2x2_ASAP7_75t_L g748 ( .A(n_685), .B(n_749), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_686), .B(n_736), .Y(n_762) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_687), .B(n_854), .Y(n_853) );
AOI22x1_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B1(n_694), .B2(n_696), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_689), .B(n_713), .Y(n_796) );
AND2x2_ASAP7_75t_L g804 ( .A(n_689), .B(n_713), .Y(n_804) );
INVx2_ASAP7_75t_L g703 ( .A(n_690), .Y(n_703) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_690), .Y(n_861) );
OAI21xp33_ASAP7_75t_L g708 ( .A1(n_691), .A2(n_709), .B(n_712), .Y(n_708) );
AND2x4_ASAP7_75t_L g744 ( .A(n_692), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g821 ( .A(n_692), .B(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g840 ( .A(n_692), .Y(n_840) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g704 ( .A(n_695), .B(n_703), .Y(n_704) );
AND2x2_ASAP7_75t_L g738 ( .A(n_695), .B(n_728), .Y(n_738) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_695), .Y(n_743) );
AND2x2_ASAP7_75t_L g845 ( .A(n_695), .B(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_708), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_700), .B(n_868), .Y(n_867) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVxp67_ASAP7_75t_SL g827 ( .A(n_702), .Y(n_827) );
AND2x2_ASAP7_75t_L g730 ( .A(n_703), .B(n_714), .Y(n_730) );
INVx1_ASAP7_75t_L g754 ( .A(n_703), .Y(n_754) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g719 ( .A(n_707), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g723 ( .A(n_707), .Y(n_723) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
NAND4xp25_ASAP7_75t_L g814 ( .A(n_713), .B(n_728), .C(n_815), .D(n_819), .Y(n_814) );
AND2x2_ASAP7_75t_L g753 ( .A(n_714), .B(n_754), .Y(n_753) );
AND2x4_ASAP7_75t_SL g714 ( .A(n_715), .B(n_716), .Y(n_714) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_721), .B(n_726), .C(n_729), .Y(n_717) );
OAI221xp5_ASAP7_75t_L g747 ( .A1(n_718), .A2(n_748), .B1(n_750), .B2(n_752), .C(n_755), .Y(n_747) );
AND2x4_ASAP7_75t_L g848 ( .A(n_719), .B(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AND2x4_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
AND2x2_ASAP7_75t_L g782 ( .A(n_724), .B(n_734), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_724), .B(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g759 ( .A(n_728), .B(n_760), .Y(n_759) );
INVxp67_ASAP7_75t_SL g830 ( .A(n_728), .Y(n_830) );
AND2x2_ASAP7_75t_SL g844 ( .A(n_728), .B(n_789), .Y(n_844) );
INVx2_ASAP7_75t_L g846 ( .A(n_728), .Y(n_846) );
NOR3xp33_ASAP7_75t_SL g731 ( .A(n_732), .B(n_739), .C(n_747), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_733), .B(n_737), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_736), .Y(n_733) );
BUFx3_ASAP7_75t_L g823 ( .A(n_734), .Y(n_823) );
AND2x2_ASAP7_75t_L g855 ( .A(n_734), .B(n_736), .Y(n_855) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx3_ASAP7_75t_L g797 ( .A(n_744), .Y(n_797) );
INVxp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OR2x6_ASAP7_75t_L g826 ( .A(n_746), .B(n_827), .Y(n_826) );
INVxp67_ASAP7_75t_SL g870 ( .A(n_746), .Y(n_870) );
INVxp67_ASAP7_75t_SL g774 ( .A(n_749), .Y(n_774) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
A2O1A1Ixp33_ASAP7_75t_L g783 ( .A1(n_753), .A2(n_784), .B(n_785), .C(n_791), .Y(n_783) );
OAI21xp33_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_759), .B(n_762), .Y(n_755) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OAI21xp5_ASAP7_75t_SL g795 ( .A1(n_758), .A2(n_779), .B(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g800 ( .A(n_758), .Y(n_800) );
INVx2_ASAP7_75t_L g836 ( .A(n_759), .Y(n_836) );
AND2x4_ASAP7_75t_L g812 ( .A(n_760), .B(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_831), .Y(n_763) );
NOR3xp33_ASAP7_75t_L g764 ( .A(n_765), .B(n_793), .C(n_805), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_776), .C(n_783), .Y(n_765) );
OAI21xp33_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_770), .B(n_775), .Y(n_766) );
INVxp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVxp67_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_769), .B(n_830), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
AND2x2_ASAP7_75t_L g799 ( .A(n_772), .B(n_800), .Y(n_799) );
OAI32xp33_ASAP7_75t_L g858 ( .A1(n_772), .A2(n_856), .A3(n_859), .B1(n_863), .B2(n_867), .Y(n_858) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OAI31xp33_ASAP7_75t_SL g776 ( .A1(n_777), .A2(n_778), .A3(n_780), .B(n_782), .Y(n_776) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
OR2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVxp67_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
OAI221xp5_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_797), .B1(n_798), .B2(n_801), .C(n_803), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NAND3xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_820), .C(n_824), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
OAI21xp5_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_811), .B(n_814), .Y(n_807) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
OAI21xp33_ASAP7_75t_L g820 ( .A1(n_812), .A2(n_821), .B(n_823), .Y(n_820) );
AND2x2_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_817), .Y(n_854) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_825), .B(n_828), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g841 ( .A(n_826), .Y(n_841) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NOR3xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_842), .C(n_858), .Y(n_831) );
AOI21x1_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_836), .B(n_837), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
AND2x4_ASAP7_75t_L g838 ( .A(n_839), .B(n_841), .Y(n_838) );
INVxp67_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OAI22xp33_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_847), .B1(n_851), .B2(n_856), .Y(n_842) );
NOR2xp33_ASAP7_75t_SL g843 ( .A(n_844), .B(n_845), .Y(n_843) );
INVx2_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
NOR2xp33_ASAP7_75t_SL g851 ( .A(n_852), .B(n_855), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx2_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
AND2x4_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .Y(n_860) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
AND2x4_ASAP7_75t_L g868 ( .A(n_869), .B(n_870), .Y(n_868) );
BUFx3_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
BUFx12f_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
CKINVDCx11_ASAP7_75t_R g873 ( .A(n_874), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
OR2x6_ASAP7_75t_L g875 ( .A(n_876), .B(n_877), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_877), .B(n_893), .Y(n_892) );
INVx2_ASAP7_75t_SL g879 ( .A(n_880), .Y(n_879) );
NOR2xp33_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
BUFx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
BUFx3_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
O2A1O1Ixp33_ASAP7_75t_SL g896 ( .A1(n_886), .A2(n_897), .B(n_902), .C(n_904), .Y(n_896) );
OR2x2_ASAP7_75t_L g886 ( .A(n_887), .B(n_888), .Y(n_886) );
INVx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
CKINVDCx5p33_ASAP7_75t_R g889 ( .A(n_890), .Y(n_889) );
BUFx12f_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
BUFx8_ASAP7_75t_L g903 ( .A(n_891), .Y(n_903) );
BUFx6f_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
BUFx3_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
HB1xp67_ASAP7_75t_L g906 ( .A(n_895), .Y(n_906) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVxp67_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
BUFx2_ASAP7_75t_SL g907 ( .A(n_908), .Y(n_907) );
BUFx3_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
CKINVDCx6p67_ASAP7_75t_R g917 ( .A(n_909), .Y(n_917) );
BUFx5_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_911), .B(n_912), .Y(n_910) );
BUFx2_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
endmodule