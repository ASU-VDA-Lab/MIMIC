module fake_ibex_758_n_2923 (n_151, n_85, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_545, n_194, n_249, n_334, n_312, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_7, n_109, n_127, n_121, n_527, n_465, n_48, n_325, n_57, n_301, n_496, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_13, n_122, n_523, n_116, n_370, n_431, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_490, n_52, n_448, n_99, n_466, n_269, n_156, n_126, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_536, n_352, n_290, n_558, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_514, n_429, n_275, n_541, n_98, n_129, n_267, n_245, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_480, n_416, n_365, n_4, n_6, n_539, n_100, n_179, n_354, n_206, n_392, n_516, n_548, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_546, n_199, n_495, n_410, n_308, n_463, n_411, n_135, n_520, n_512, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_517, n_211, n_218, n_314, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_532, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_476, n_461, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_311, n_406, n_97, n_197, n_528, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_2923);

input n_151;
input n_85;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_194;
input n_249;
input n_334;
input n_312;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_523;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_490;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_126;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_536;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_514;
input n_429;
input n_275;
input n_541;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_480;
input n_416;
input n_365;
input n_4;
input n_6;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_516;
input n_548;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_546;
input n_199;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_520;
input n_512;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_476;
input n_461;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_2923;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_2569;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_1079;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_969;
wire n_678;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_1308;
wire n_1138;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_667;
wire n_884;
wire n_2396;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2724;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_641;
wire n_1937;
wire n_2311;
wire n_893;
wire n_1654;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_852;
wire n_1427;
wire n_1133;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2814;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2922;
wire n_2347;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_1955;
wire n_917;
wire n_2413;
wire n_2249;
wire n_2362;
wire n_968;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_2090;
wire n_666;
wire n_2260;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1960;
wire n_1723;
wire n_2663;
wire n_793;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_2906;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_605;
wire n_2373;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_971;
wire n_1326;
wire n_702;
wire n_1350;
wire n_906;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_2541;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_2723;
wire n_1616;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_2256;
wire n_606;
wire n_737;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2879;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_2573;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_591;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_2838;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_594;
wire n_2361;
wire n_1566;
wire n_1464;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_660;
wire n_2590;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_576;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_607;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2823;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_2010;
wire n_1756;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_2905;
wire n_803;
wire n_2570;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_2095;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2352;
wire n_2212;
wire n_2716;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_2903;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_2654;
wire n_2463;
wire n_717;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_588;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_916;
wire n_2298;
wire n_2771;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_2772;
wire n_2778;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_626;
wire n_1941;
wire n_1707;
wire n_2422;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_2862;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_598;
wire n_2141;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_2920;
wire n_604;
wire n_1598;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_1625;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_636;
wire n_1259;
wire n_2108;
wire n_2535;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2709;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_2665;
wire n_1124;
wire n_611;
wire n_1690;
wire n_2688;
wire n_2881;
wire n_1673;
wire n_2018;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_2758;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_2845;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_2447;
wire n_2818;
wire n_1057;
wire n_1473;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_775;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_2608;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_616;
wire n_1885;
wire n_1989;
wire n_1740;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2861;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2803;
wire n_2816;
wire n_2433;
wire n_1256;
wire n_2798;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_1961;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_688;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_2518;
wire n_2784;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_1029;
wire n_2394;
wire n_770;
wire n_1635;
wire n_1572;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_2323;
wire n_740;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_1986;
wire n_2882;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_2734;
wire n_2870;
wire n_758;
wire n_1166;
wire n_720;
wire n_1390;
wire n_710;
wire n_2775;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_580;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_999;
wire n_2634;
wire n_1092;
wire n_1808;
wire n_560;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_2492;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_1142;
wire n_783;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2357;
wire n_2303;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_924;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_2092;
wire n_566;
wire n_581;
wire n_1365;
wire n_1472;
wire n_2443;
wire n_2802;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2704;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_1736;
wire n_2907;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_2754;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_2673;
wire n_2676;
wire n_921;
wire n_2430;
wire n_1534;
wire n_2912;
wire n_908;
wire n_1346;
wire n_565;
wire n_2834;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_866;

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_102),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_208),
.Y(n_561)
);

BUFx10_ASAP7_75t_L g562 ( 
.A(n_204),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_500),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_156),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_100),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_508),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_276),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_531),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_117),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_370),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_292),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_399),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_232),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_221),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_207),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_12),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_100),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_492),
.Y(n_578)
);

BUFx8_ASAP7_75t_SL g579 ( 
.A(n_39),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_254),
.Y(n_580)
);

CKINVDCx14_ASAP7_75t_R g581 ( 
.A(n_317),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_225),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_175),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_392),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_533),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_284),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_390),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_222),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_476),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_466),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_306),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_538),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_349),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_214),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_219),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_139),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_486),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_541),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_458),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_323),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_301),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_61),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_465),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_537),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_82),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_110),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_37),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_182),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_37),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_331),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_112),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_98),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_3),
.Y(n_613)
);

BUFx10_ASAP7_75t_L g614 ( 
.A(n_471),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_59),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_222),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_130),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_423),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_542),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_407),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_280),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_432),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_158),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_31),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_342),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_308),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_358),
.Y(n_627)
);

CKINVDCx16_ASAP7_75t_R g628 ( 
.A(n_398),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_506),
.Y(n_629)
);

BUFx10_ASAP7_75t_L g630 ( 
.A(n_228),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_280),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_70),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_237),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_186),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_532),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_54),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_148),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_248),
.Y(n_638)
);

BUFx10_ASAP7_75t_L g639 ( 
.A(n_515),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_38),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_443),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_233),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_344),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_539),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_505),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_225),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_128),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_452),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_418),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_315),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_356),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_168),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_289),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_252),
.Y(n_654)
);

CKINVDCx16_ASAP7_75t_R g655 ( 
.A(n_424),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_252),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_76),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_416),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_433),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_297),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_255),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_549),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_341),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_395),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_43),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_263),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_546),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_121),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_28),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_282),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_347),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_298),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_21),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_322),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_497),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_365),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_113),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_220),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_234),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_540),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_259),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_101),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_264),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_359),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_305),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_363),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_385),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_522),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_109),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_350),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_455),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_190),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_302),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_548),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_63),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_111),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_241),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_255),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_467),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_351),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_402),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_62),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_346),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_420),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_85),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_78),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_382),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_551),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_273),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_215),
.Y(n_710)
);

CKINVDCx16_ASAP7_75t_R g711 ( 
.A(n_406),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_85),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_374),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_459),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_534),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_439),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_4),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_447),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_478),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_181),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_545),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_362),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_186),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_435),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_485),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_501),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_232),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_48),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_122),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_101),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_357),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_128),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_184),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_517),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_348),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_326),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_143),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_324),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_45),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_290),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_23),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_131),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_97),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_147),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_277),
.B(n_290),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_38),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_166),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_223),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_507),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_441),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_25),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_72),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_278),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_417),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_431),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_262),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_137),
.Y(n_757)
);

INVx1_ASAP7_75t_SL g758 ( 
.A(n_224),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_105),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_284),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_328),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_144),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_36),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_44),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_314),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_267),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_249),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_391),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_529),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_269),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_553),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_388),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_195),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_451),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_241),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_10),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_150),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_555),
.Y(n_778)
);

CKINVDCx14_ASAP7_75t_R g779 ( 
.A(n_79),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_526),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_151),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_201),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_343),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_400),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_520),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_513),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_170),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_65),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_121),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_224),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_155),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_396),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_256),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_278),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_23),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_136),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_L g797 ( 
.A(n_161),
.B(n_352),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_332),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_94),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_488),
.Y(n_800)
);

NOR2xp67_ASAP7_75t_L g801 ( 
.A(n_68),
.B(n_405),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_335),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_462),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_62),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_519),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_34),
.Y(n_806)
);

NOR2xp67_ASAP7_75t_L g807 ( 
.A(n_368),
.B(n_345),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_387),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_244),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_394),
.Y(n_810)
);

NOR2xp67_ASAP7_75t_L g811 ( 
.A(n_448),
.B(n_487),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_134),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_554),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_208),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_521),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_58),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_248),
.Y(n_817)
);

BUFx10_ASAP7_75t_L g818 ( 
.A(n_360),
.Y(n_818)
);

CKINVDCx14_ASAP7_75t_R g819 ( 
.A(n_414),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_2),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_307),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_96),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_40),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_180),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_299),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_550),
.Y(n_826)
);

BUFx10_ASAP7_75t_L g827 ( 
.A(n_20),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_509),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_143),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_263),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_198),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_355),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_287),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_461),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_250),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_176),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_22),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_474),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_149),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_490),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_376),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_512),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_243),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_523),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_207),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_354),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_293),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_32),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_258),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_25),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_336),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_329),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_211),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_446),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_496),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_8),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_2),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_518),
.Y(n_858)
);

BUFx2_ASAP7_75t_SL g859 ( 
.A(n_91),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_15),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_179),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_473),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_93),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_384),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_194),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_491),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_353),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_214),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_457),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_469),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_176),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_377),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_53),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_291),
.Y(n_874)
);

INVxp67_ASAP7_75t_SL g875 ( 
.A(n_235),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_148),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_238),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_109),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_503),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_6),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_453),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_210),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_48),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_164),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_235),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_456),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_175),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_504),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_70),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_7),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_311),
.Y(n_891)
);

BUFx8_ASAP7_75t_SL g892 ( 
.A(n_552),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_135),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_404),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_91),
.Y(n_895)
);

BUFx10_ASAP7_75t_L g896 ( 
.A(n_481),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_645),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_779),
.A2(n_3),
.B1(n_0),
.B2(n_1),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_605),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_605),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_779),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_579),
.Y(n_902)
);

INVx5_ASAP7_75t_L g903 ( 
.A(n_645),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_562),
.Y(n_904)
);

OAI22x1_ASAP7_75t_SL g905 ( 
.A1(n_564),
.A2(n_4),
.B1(n_0),
.B2(n_1),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_578),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_579),
.Y(n_907)
);

CKINVDCx16_ASAP7_75t_R g908 ( 
.A(n_628),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_707),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_634),
.Y(n_910)
);

INVx6_ASAP7_75t_L g911 ( 
.A(n_614),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_578),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_892),
.Y(n_913)
);

INVx4_ASAP7_75t_L g914 ( 
.A(n_707),
.Y(n_914)
);

OAI21x1_ASAP7_75t_L g915 ( 
.A1(n_707),
.A2(n_310),
.B(n_309),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_562),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_684),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_786),
.B(n_5),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_SL g919 ( 
.A1(n_564),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_602),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_562),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_614),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_634),
.B(n_9),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_630),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_578),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_642),
.Y(n_926)
);

INVx5_ASAP7_75t_L g927 ( 
.A(n_614),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_767),
.B(n_9),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_803),
.B(n_10),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_578),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_625),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_625),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_642),
.B(n_11),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_747),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_747),
.Y(n_935)
);

BUFx12f_ASAP7_75t_L g936 ( 
.A(n_630),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_794),
.Y(n_937)
);

INVxp67_ASAP7_75t_L g938 ( 
.A(n_631),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_625),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_803),
.B(n_11),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_869),
.B(n_13),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_794),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_762),
.B(n_13),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_655),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_895),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_869),
.B(n_14),
.Y(n_946)
);

OA21x2_ASAP7_75t_L g947 ( 
.A1(n_590),
.A2(n_313),
.B(n_312),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_625),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_833),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_861),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_861),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_573),
.B(n_16),
.Y(n_952)
);

OAI21x1_ASAP7_75t_L g953 ( 
.A1(n_590),
.A2(n_318),
.B(n_316),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_699),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_561),
.B(n_17),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_699),
.Y(n_956)
);

OA21x2_ASAP7_75t_L g957 ( 
.A1(n_604),
.A2(n_320),
.B(n_319),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_573),
.B(n_580),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_699),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_647),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_684),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_647),
.Y(n_962)
);

INVx5_ASAP7_75t_L g963 ( 
.A(n_639),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_699),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_892),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_580),
.B(n_17),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_742),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_862),
.Y(n_968)
);

BUFx8_ASAP7_75t_SL g969 ( 
.A(n_594),
.Y(n_969)
);

INVx5_ASAP7_75t_L g970 ( 
.A(n_639),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_742),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_848),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_630),
.B(n_18),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_862),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_717),
.B(n_18),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_711),
.Y(n_976)
);

BUFx8_ASAP7_75t_SL g977 ( 
.A(n_594),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_565),
.B(n_19),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_793),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_647),
.Y(n_980)
);

OA21x2_ASAP7_75t_L g981 ( 
.A1(n_604),
.A2(n_325),
.B(n_321),
.Y(n_981)
);

INVx5_ASAP7_75t_L g982 ( 
.A(n_639),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_848),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_569),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_575),
.B(n_19),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_576),
.Y(n_986)
);

AOI22x1_ASAP7_75t_SL g987 ( 
.A1(n_601),
.A2(n_612),
.B1(n_652),
.B2(n_636),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_588),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_SL g989 ( 
.A1(n_601),
.A2(n_24),
.B1(n_21),
.B2(n_22),
.Y(n_989)
);

OAI21x1_ASAP7_75t_L g990 ( 
.A1(n_651),
.A2(n_330),
.B(n_327),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_560),
.Y(n_991)
);

AOI22x1_ASAP7_75t_SL g992 ( 
.A1(n_612),
.A2(n_27),
.B1(n_24),
.B2(n_26),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_608),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_615),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_862),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_651),
.A2(n_334),
.B(n_333),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_913),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_913),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_908),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_911),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_965),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_965),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_969),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_969),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_977),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_977),
.Y(n_1006)
);

BUFx10_ASAP7_75t_L g1007 ( 
.A(n_911),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_976),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_976),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_R g1010 ( 
.A(n_904),
.B(n_581),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_902),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_936),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_R g1013 ( 
.A(n_904),
.B(n_581),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_902),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_907),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_907),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_901),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_991),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_901),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_987),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_935),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_920),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_922),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_922),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_920),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_945),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_917),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_945),
.Y(n_1028)
);

CKINVDCx20_ASAP7_75t_R g1029 ( 
.A(n_938),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_933),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_979),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_911),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_952),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_938),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_R g1035 ( 
.A(n_916),
.B(n_819),
.Y(n_1035)
);

CKINVDCx14_ASAP7_75t_R g1036 ( 
.A(n_927),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_R g1037 ( 
.A(n_916),
.B(n_921),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_927),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_927),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_906),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_952),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_927),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_963),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_963),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_973),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_963),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_963),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_970),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_906),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_970),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_970),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_970),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_921),
.B(n_571),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_982),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_949),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_982),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_966),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_949),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_961),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_966),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_982),
.Y(n_1061)
);

AND3x2_ASAP7_75t_L g1062 ( 
.A(n_918),
.B(n_875),
.C(n_586),
.Y(n_1062)
);

CKINVDCx20_ASAP7_75t_R g1063 ( 
.A(n_928),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_958),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_899),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_900),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_R g1067 ( 
.A(n_924),
.B(n_819),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_982),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_909),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_924),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_897),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_992),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_910),
.Y(n_1073)
);

INVx2_ASAP7_75t_SL g1074 ( 
.A(n_909),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_905),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_906),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_943),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_989),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_985),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_985),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_919),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_R g1082 ( 
.A(n_926),
.B(n_618),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_914),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_897),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_898),
.Y(n_1085)
);

OR2x2_ASAP7_75t_L g1086 ( 
.A(n_984),
.B(n_574),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_944),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_918),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_R g1089 ( 
.A(n_914),
.B(n_618),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_986),
.B(n_736),
.Y(n_1090)
);

AND2x6_ASAP7_75t_L g1091 ( 
.A(n_929),
.B(n_718),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_923),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_929),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_988),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_903),
.B(n_585),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_934),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_937),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_942),
.Y(n_1098)
);

BUFx10_ASAP7_75t_L g1099 ( 
.A(n_975),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_950),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_940),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_951),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_903),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_940),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_941),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_993),
.B(n_774),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_903),
.B(n_585),
.Y(n_1107)
);

INVxp33_ASAP7_75t_SL g1108 ( 
.A(n_975),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_994),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_946),
.Y(n_1110)
);

OR2x2_ASAP7_75t_L g1111 ( 
.A(n_967),
.B(n_577),
.Y(n_1111)
);

CKINVDCx16_ASAP7_75t_R g1112 ( 
.A(n_946),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_903),
.B(n_818),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_971),
.B(n_774),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_955),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_955),
.Y(n_1116)
);

NOR2xp67_ASAP7_75t_L g1117 ( 
.A(n_972),
.B(n_563),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_978),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_983),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_960),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_915),
.Y(n_1121)
);

CKINVDCx16_ASAP7_75t_R g1122 ( 
.A(n_962),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_953),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_947),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_980),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_912),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_990),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_996),
.Y(n_1128)
);

INVx4_ASAP7_75t_L g1129 ( 
.A(n_947),
.Y(n_1129)
);

OAI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_957),
.A2(n_652),
.B1(n_766),
.B2(n_636),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_957),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_981),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_912),
.B(n_583),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_925),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_925),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_925),
.B(n_587),
.Y(n_1136)
);

INVxp33_ASAP7_75t_SL g1137 ( 
.A(n_981),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_930),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_930),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_930),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_931),
.Y(n_1141)
);

CKINVDCx20_ASAP7_75t_R g1142 ( 
.A(n_931),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_931),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_R g1144 ( 
.A(n_932),
.B(n_641),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_932),
.Y(n_1145)
);

CKINVDCx16_ASAP7_75t_R g1146 ( 
.A(n_932),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_939),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_939),
.Y(n_1148)
);

NAND2xp33_ASAP7_75t_R g1149 ( 
.A(n_939),
.B(n_883),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_948),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_948),
.B(n_818),
.Y(n_1151)
);

CKINVDCx16_ASAP7_75t_R g1152 ( 
.A(n_954),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_995),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_954),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_956),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_956),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_956),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_959),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_959),
.B(n_587),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_964),
.Y(n_1160)
);

AOI21x1_ASAP7_75t_L g1161 ( 
.A1(n_964),
.A2(n_872),
.B(n_785),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_968),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_968),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_968),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_974),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_974),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_995),
.Y(n_1167)
);

CKINVDCx20_ASAP7_75t_R g1168 ( 
.A(n_995),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_911),
.B(n_785),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_R g1170 ( 
.A(n_913),
.B(n_641),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_R g1171 ( 
.A(n_913),
.B(n_644),
.Y(n_1171)
);

AOI21x1_ASAP7_75t_L g1172 ( 
.A1(n_953),
.A2(n_872),
.B(n_591),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_913),
.Y(n_1173)
);

AND3x1_ASAP7_75t_L g1174 ( 
.A(n_944),
.B(n_633),
.C(n_632),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_922),
.B(n_818),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1069),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1092),
.B(n_896),
.Y(n_1177)
);

OR2x6_ASAP7_75t_L g1178 ( 
.A(n_1012),
.B(n_859),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_L g1179 ( 
.A(n_1105),
.B(n_745),
.C(n_600),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1112),
.B(n_566),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1069),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1142),
.Y(n_1182)
);

NAND2xp33_ASAP7_75t_L g1183 ( 
.A(n_1010),
.B(n_568),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1065),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_SL g1185 ( 
.A1(n_1089),
.A2(n_820),
.B1(n_823),
.B2(n_766),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1175),
.B(n_896),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1059),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1022),
.B(n_827),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1168),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1022),
.B(n_827),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1121),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1110),
.B(n_570),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1108),
.B(n_598),
.Y(n_1193)
);

OR2x2_ASAP7_75t_L g1194 ( 
.A(n_1025),
.B(n_606),
.Y(n_1194)
);

INVxp33_ASAP7_75t_L g1195 ( 
.A(n_1170),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1066),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1115),
.B(n_1116),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1094),
.B(n_572),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1118),
.B(n_589),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1073),
.Y(n_1200)
);

NAND3xp33_ASAP7_75t_L g1201 ( 
.A(n_1129),
.B(n_626),
.C(n_610),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1023),
.B(n_1024),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_1017),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1030),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1055),
.B(n_584),
.Y(n_1205)
);

INVxp67_ASAP7_75t_L g1206 ( 
.A(n_1034),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1096),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1109),
.B(n_592),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1026),
.B(n_567),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1021),
.Y(n_1210)
);

NAND2xp33_ASAP7_75t_L g1211 ( 
.A(n_1013),
.B(n_593),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1169),
.B(n_597),
.Y(n_1212)
);

NOR2xp67_ASAP7_75t_L g1213 ( 
.A(n_1028),
.B(n_27),
.Y(n_1213)
);

INVx4_ASAP7_75t_L g1214 ( 
.A(n_1146),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1000),
.B(n_721),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1093),
.B(n_599),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1097),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1013),
.B(n_603),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1058),
.B(n_582),
.Y(n_1219)
);

INVxp67_ASAP7_75t_L g1220 ( 
.A(n_1031),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1070),
.B(n_724),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1098),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1100),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1102),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1119),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1071),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1133),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1033),
.B(n_627),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1083),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_SL g1230 ( 
.A(n_1124),
.B(n_644),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1064),
.B(n_826),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1090),
.B(n_619),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1084),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1172),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1079),
.B(n_858),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1080),
.B(n_864),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1035),
.B(n_620),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1099),
.B(n_622),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1041),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1103),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1099),
.B(n_629),
.Y(n_1241)
);

INVxp67_ASAP7_75t_SL g1242 ( 
.A(n_1029),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1154),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1074),
.B(n_643),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1057),
.B(n_648),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1060),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1117),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1131),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1114),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1036),
.B(n_649),
.Y(n_1250)
);

NOR3xp33_ASAP7_75t_L g1251 ( 
.A(n_1130),
.B(n_737),
.C(n_609),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1114),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1106),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1106),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1054),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1111),
.Y(n_1256)
);

INVxp33_ASAP7_75t_L g1257 ( 
.A(n_1170),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1131),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1086),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1136),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1067),
.B(n_659),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1122),
.B(n_664),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1019),
.B(n_671),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1161),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1159),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1037),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1091),
.B(n_674),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1120),
.Y(n_1268)
);

NOR3xp33_ASAP7_75t_L g1269 ( 
.A(n_1130),
.B(n_758),
.C(n_746),
.Y(n_1269)
);

BUFx8_ASAP7_75t_L g1270 ( 
.A(n_1053),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1132),
.B(n_1137),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1091),
.B(n_687),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1125),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1091),
.B(n_635),
.Y(n_1274)
);

BUFx5_ASAP7_75t_L g1275 ( 
.A(n_1123),
.Y(n_1275)
);

NOR2x1p5_ASAP7_75t_L g1276 ( 
.A(n_1004),
.B(n_595),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1032),
.B(n_688),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1127),
.B(n_650),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1128),
.B(n_658),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1095),
.B(n_667),
.Y(n_1280)
);

NAND2x1p5_ASAP7_75t_L g1281 ( 
.A(n_1113),
.B(n_640),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1151),
.Y(n_1282)
);

INVx4_ASAP7_75t_L g1283 ( 
.A(n_1152),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1068),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1107),
.B(n_675),
.Y(n_1285)
);

INVxp67_ASAP7_75t_L g1286 ( 
.A(n_1018),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1038),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1039),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1088),
.B(n_691),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1077),
.B(n_596),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_SL g1291 ( 
.A(n_1006),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1042),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1067),
.B(n_676),
.Y(n_1293)
);

INVx1_ASAP7_75t_SL g1294 ( 
.A(n_1089),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1082),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_997),
.Y(n_1296)
);

INVxp33_ASAP7_75t_L g1297 ( 
.A(n_1171),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_SL g1298 ( 
.A(n_1008),
.B(n_662),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1043),
.B(n_680),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1044),
.B(n_1046),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1126),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1047),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1048),
.B(n_1050),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1148),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1134),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1051),
.B(n_690),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1052),
.B(n_694),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1144),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1101),
.B(n_701),
.Y(n_1309)
);

INVx8_ASAP7_75t_L g1310 ( 
.A(n_1056),
.Y(n_1310)
);

NOR3xp33_ASAP7_75t_L g1311 ( 
.A(n_1081),
.B(n_795),
.C(n_611),
.Y(n_1311)
);

NOR3xp33_ASAP7_75t_L g1312 ( 
.A(n_1078),
.B(n_613),
.C(n_607),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1062),
.B(n_662),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1061),
.B(n_713),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1045),
.B(n_714),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1082),
.B(n_715),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1062),
.B(n_716),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1009),
.B(n_719),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_R g1319 ( 
.A(n_999),
.B(n_663),
.Y(n_1319)
);

OAI21xp33_ASAP7_75t_L g1320 ( 
.A1(n_1144),
.A2(n_666),
.B(n_657),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1171),
.Y(n_1321)
);

NOR2xp67_ASAP7_75t_L g1322 ( 
.A(n_998),
.B(n_29),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1135),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1138),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1063),
.B(n_722),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1001),
.B(n_725),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1139),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1174),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1002),
.B(n_726),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1173),
.B(n_734),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1143),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1145),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1147),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1156),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1157),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1167),
.B(n_755),
.Y(n_1336)
);

NOR2xp67_ASAP7_75t_L g1337 ( 
.A(n_1072),
.B(n_29),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1085),
.B(n_771),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1158),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1164),
.Y(n_1340)
);

NAND3xp33_ASAP7_75t_L g1341 ( 
.A(n_1149),
.B(n_703),
.C(n_700),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1165),
.B(n_783),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1166),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1087),
.B(n_792),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1141),
.Y(n_1345)
);

NAND3xp33_ASAP7_75t_L g1346 ( 
.A(n_1149),
.B(n_731),
.C(n_708),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1153),
.B(n_735),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1153),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1003),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1011),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1160),
.B(n_798),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1162),
.B(n_738),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1163),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1014),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1040),
.B(n_800),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1140),
.B(n_802),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1075),
.B(n_805),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1155),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1040),
.Y(n_1359)
);

INVxp67_ASAP7_75t_SL g1360 ( 
.A(n_1005),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1150),
.B(n_808),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1015),
.B(n_616),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1016),
.B(n_813),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1150),
.B(n_821),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1040),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1040),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1049),
.B(n_828),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1076),
.Y(n_1368)
);

NAND2xp33_ASAP7_75t_L g1369 ( 
.A(n_1049),
.B(n_832),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1020),
.B(n_834),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1049),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1049),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1076),
.B(n_617),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1076),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1069),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1092),
.B(n_838),
.Y(n_1376)
);

A2O1A1Ixp33_ASAP7_75t_L g1377 ( 
.A1(n_1104),
.A2(n_672),
.B(n_677),
.C(n_669),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1069),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_L g1379 ( 
.A(n_1104),
.B(n_754),
.C(n_750),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1007),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1069),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1069),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1104),
.B(n_840),
.Y(n_1383)
);

NAND3xp33_ASAP7_75t_L g1384 ( 
.A(n_1104),
.B(n_765),
.C(n_761),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1069),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1104),
.B(n_841),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1069),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1069),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1069),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1112),
.B(n_846),
.Y(n_1390)
);

AND2x2_ASAP7_75t_SL g1391 ( 
.A(n_1174),
.B(n_663),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1069),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1069),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1112),
.B(n_851),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1112),
.B(n_852),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1112),
.B(n_854),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1104),
.B(n_768),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1104),
.B(n_769),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1104),
.B(n_772),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1092),
.A2(n_681),
.B1(n_685),
.B2(n_678),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1069),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1112),
.B(n_855),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1092),
.B(n_879),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1069),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1092),
.B(n_881),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1027),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1069),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1104),
.B(n_778),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1069),
.Y(n_1409)
);

NOR2xp67_ASAP7_75t_L g1410 ( 
.A(n_1012),
.B(n_30),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1069),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1104),
.B(n_780),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1184),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1191),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1214),
.B(n_686),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1197),
.A2(n_704),
.B1(n_749),
.B2(n_686),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1270),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1191),
.Y(n_1418)
);

OR2x4_ASAP7_75t_L g1419 ( 
.A(n_1338),
.B(n_820),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1196),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1200),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1229),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1251),
.A2(n_837),
.B1(n_845),
.B2(n_823),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1182),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1248),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1256),
.B(n_621),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1242),
.Y(n_1427)
);

NAND3xp33_ASAP7_75t_SL g1428 ( 
.A(n_1269),
.B(n_749),
.C(n_704),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1197),
.B(n_837),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1294),
.B(n_886),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1397),
.B(n_623),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1259),
.B(n_845),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1397),
.B(n_624),
.Y(n_1433)
);

NAND2x1p5_ASAP7_75t_L g1434 ( 
.A(n_1214),
.B(n_689),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1270),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1398),
.B(n_637),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_SL g1437 ( 
.A1(n_1391),
.A2(n_877),
.B1(n_889),
.B2(n_876),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1398),
.B(n_1399),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1283),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1203),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1191),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1325),
.B(n_876),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1271),
.A2(n_889),
.B1(n_877),
.B2(n_702),
.Y(n_1443)
);

AND2x6_ASAP7_75t_SL g1444 ( 
.A(n_1178),
.B(n_698),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1207),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1188),
.B(n_638),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1253),
.A2(n_712),
.B(n_720),
.C(n_709),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1319),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_1189),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1399),
.B(n_646),
.Y(n_1450)
);

INVx5_ASAP7_75t_L g1451 ( 
.A(n_1310),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1217),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1284),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1222),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1230),
.A2(n_654),
.B1(n_656),
.B2(n_653),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1278),
.A2(n_1279),
.B(n_1274),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1408),
.B(n_660),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1227),
.B(n_727),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1220),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1408),
.B(n_661),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1291),
.Y(n_1461)
);

AND2x6_ASAP7_75t_L g1462 ( 
.A(n_1258),
.B(n_718),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1412),
.B(n_665),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1243),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1296),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1412),
.B(n_673),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1258),
.Y(n_1467)
);

BUFx4f_ASAP7_75t_L g1468 ( 
.A(n_1178),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1178),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1199),
.B(n_679),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1179),
.A2(n_1176),
.B1(n_1375),
.B2(n_1181),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1199),
.B(n_682),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1304),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1223),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1380),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1224),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1206),
.B(n_683),
.Y(n_1477)
);

AOI21xp33_ASAP7_75t_L g1478 ( 
.A1(n_1193),
.A2(n_1289),
.B(n_1190),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1219),
.B(n_1180),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1271),
.A2(n_732),
.B1(n_739),
.B2(n_728),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1194),
.Y(n_1481)
);

INVx2_ASAP7_75t_SL g1482 ( 
.A(n_1310),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1390),
.B(n_692),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_1310),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1287),
.B(n_740),
.Y(n_1485)
);

O2A1O1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1377),
.A2(n_751),
.B(n_752),
.C(n_741),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1179),
.A2(n_756),
.B1(n_759),
.B2(n_753),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1298),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1286),
.B(n_693),
.Y(n_1489)
);

OR2x4_ASAP7_75t_L g1490 ( 
.A(n_1344),
.B(n_760),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1378),
.B(n_695),
.Y(n_1491)
);

AOI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1204),
.A2(n_770),
.B1(n_775),
.B2(n_764),
.Y(n_1492)
);

INVx5_ASAP7_75t_L g1493 ( 
.A(n_1304),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1239),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1381),
.A2(n_788),
.B1(n_789),
.B2(n_777),
.Y(n_1495)
);

AOI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1246),
.A2(n_791),
.B1(n_804),
.B2(n_796),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1382),
.B(n_696),
.Y(n_1497)
);

BUFx6f_ASAP7_75t_L g1498 ( 
.A(n_1304),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1385),
.B(n_697),
.Y(n_1499)
);

INVx4_ASAP7_75t_L g1500 ( 
.A(n_1295),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1209),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1321),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1387),
.B(n_705),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1254),
.A2(n_814),
.B1(n_817),
.B2(n_812),
.Y(n_1504)
);

NOR2x1p5_ASAP7_75t_L g1505 ( 
.A(n_1313),
.B(n_706),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1185),
.B(n_710),
.Y(n_1506)
);

NAND2x1p5_ASAP7_75t_L g1507 ( 
.A(n_1266),
.B(n_822),
.Y(n_1507)
);

NAND2x1p5_ASAP7_75t_L g1508 ( 
.A(n_1308),
.B(n_825),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1210),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1394),
.B(n_1395),
.Y(n_1510)
);

AOI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1278),
.A2(n_811),
.B(n_807),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1225),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1288),
.B(n_839),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1290),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1234),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1292),
.B(n_843),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1388),
.B(n_723),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1396),
.B(n_729),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1389),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1402),
.B(n_730),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1392),
.Y(n_1521)
);

BUFx6f_ASAP7_75t_L g1522 ( 
.A(n_1234),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1393),
.B(n_733),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1234),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1401),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1350),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1404),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1313),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1309),
.B(n_743),
.Y(n_1529)
);

OR2x6_ASAP7_75t_L g1530 ( 
.A(n_1354),
.B(n_856),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1411),
.A2(n_1409),
.B1(n_1407),
.B2(n_1379),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1315),
.B(n_744),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1260),
.Y(n_1533)
);

INVxp67_ASAP7_75t_L g1534 ( 
.A(n_1230),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1349),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1265),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1263),
.B(n_748),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1291),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1281),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1379),
.A2(n_871),
.B1(n_878),
.B2(n_865),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1177),
.B(n_757),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1376),
.B(n_763),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1255),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1362),
.B(n_1328),
.Y(n_1544)
);

BUFx4f_ASAP7_75t_L g1545 ( 
.A(n_1281),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1403),
.B(n_773),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1405),
.B(n_776),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1347),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1249),
.B(n_781),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1205),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1252),
.B(n_782),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1373),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1349),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1360),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1187),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1384),
.A2(n_884),
.B1(n_810),
.B2(n_815),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1240),
.Y(n_1557)
);

AND2x6_ASAP7_75t_L g1558 ( 
.A(n_1274),
.B(n_784),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1247),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1301),
.Y(n_1560)
);

BUFx12f_ASAP7_75t_L g1561 ( 
.A(n_1276),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1279),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1383),
.B(n_787),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1386),
.B(n_790),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1213),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1262),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1384),
.A2(n_670),
.B1(n_836),
.B2(n_668),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1228),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1341),
.A2(n_894),
.B1(n_842),
.B2(n_844),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1208),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1235),
.B(n_799),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_SL g1572 ( 
.A1(n_1238),
.A2(n_809),
.B1(n_816),
.B2(n_806),
.Y(n_1572)
);

INVxp67_ASAP7_75t_SL g1573 ( 
.A(n_1275),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1236),
.B(n_824),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_SL g1575 ( 
.A(n_1202),
.B(n_893),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1192),
.B(n_829),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1400),
.B(n_830),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1228),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1241),
.B(n_831),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1406),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1226),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1341),
.A2(n_670),
.B1(n_836),
.B2(n_668),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1233),
.Y(n_1583)
);

INVx1_ASAP7_75t_SL g1584 ( 
.A(n_1250),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1293),
.B(n_835),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1352),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1264),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1302),
.B(n_1268),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1410),
.Y(n_1589)
);

NOR2x1p5_ASAP7_75t_L g1590 ( 
.A(n_1317),
.B(n_847),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1198),
.B(n_849),
.Y(n_1591)
);

O2A1O1Ixp33_ASAP7_75t_L g1592 ( 
.A1(n_1311),
.A2(n_870),
.B(n_888),
.C(n_866),
.Y(n_1592)
);

NOR3xp33_ASAP7_75t_SL g1593 ( 
.A(n_1357),
.B(n_853),
.C(n_850),
.Y(n_1593)
);

AND2x6_ASAP7_75t_SL g1594 ( 
.A(n_1370),
.B(n_891),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1221),
.A2(n_860),
.B1(n_863),
.B2(n_857),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1231),
.B(n_868),
.Y(n_1596)
);

O2A1O1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1320),
.A2(n_801),
.B(n_797),
.C(n_873),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1346),
.A2(n_882),
.B1(n_885),
.B2(n_874),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1245),
.B(n_890),
.Y(n_1599)
);

BUFx2_ASAP7_75t_SL g1600 ( 
.A(n_1322),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1293),
.B(n_887),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1300),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1273),
.B(n_670),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1346),
.A2(n_836),
.B1(n_880),
.B2(n_670),
.Y(n_1604)
);

NAND2x1p5_ASAP7_75t_L g1605 ( 
.A(n_1316),
.B(n_836),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1299),
.Y(n_1606)
);

AND2x6_ASAP7_75t_SL g1607 ( 
.A(n_1363),
.B(n_26),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1280),
.A2(n_880),
.B1(n_867),
.B2(n_862),
.Y(n_1608)
);

O2A1O1Ixp5_ASAP7_75t_L g1609 ( 
.A1(n_1201),
.A2(n_867),
.B(n_880),
.C(n_338),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1352),
.Y(n_1610)
);

AND2x6_ASAP7_75t_SL g1611 ( 
.A(n_1326),
.B(n_30),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1280),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1267),
.B(n_867),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1285),
.Y(n_1614)
);

OR2x2_ASAP7_75t_SL g1615 ( 
.A(n_1195),
.B(n_867),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1285),
.Y(n_1616)
);

BUFx4f_ASAP7_75t_L g1617 ( 
.A(n_1333),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1232),
.B(n_31),
.Y(n_1618)
);

INVx2_ASAP7_75t_SL g1619 ( 
.A(n_1305),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1216),
.B(n_32),
.Y(n_1620)
);

NAND3xp33_ASAP7_75t_L g1621 ( 
.A(n_1299),
.B(n_33),
.C(n_34),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1272),
.B(n_35),
.Y(n_1622)
);

INVx5_ASAP7_75t_L g1623 ( 
.A(n_1323),
.Y(n_1623)
);

OR2x6_ASAP7_75t_L g1624 ( 
.A(n_1337),
.B(n_35),
.Y(n_1624)
);

AND3x2_ASAP7_75t_SL g1625 ( 
.A(n_1257),
.B(n_36),
.C(n_39),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1297),
.B(n_40),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1244),
.B(n_41),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1282),
.B(n_42),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1324),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1306),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1327),
.Y(n_1631)
);

NAND2x1p5_ASAP7_75t_L g1632 ( 
.A(n_1218),
.B(n_1237),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1331),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1318),
.B(n_1329),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_1330),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1332),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1300),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1340),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1303),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1312),
.B(n_43),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1186),
.B(n_44),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1334),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1345),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1335),
.Y(n_1644)
);

AOI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1212),
.A2(n_49),
.B1(n_46),
.B2(n_47),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1277),
.B(n_46),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1339),
.A2(n_50),
.B1(n_47),
.B2(n_49),
.Y(n_1647)
);

INVx1_ASAP7_75t_SL g1648 ( 
.A(n_1303),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1215),
.B(n_51),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1343),
.B(n_1261),
.Y(n_1650)
);

OR2x6_ASAP7_75t_L g1651 ( 
.A(n_1342),
.B(n_51),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1355),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1351),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1307),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1183),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1211),
.B(n_52),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1314),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1336),
.B(n_55),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1361),
.Y(n_1659)
);

INVx4_ASAP7_75t_L g1660 ( 
.A(n_1264),
.Y(n_1660)
);

BUFx4f_ASAP7_75t_L g1661 ( 
.A(n_1264),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1364),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1353),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1356),
.B(n_56),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1367),
.B(n_57),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1369),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1358),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1348),
.A2(n_63),
.B1(n_60),
.B2(n_61),
.Y(n_1668)
);

OAI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1359),
.A2(n_339),
.B(n_337),
.Y(n_1669)
);

INVx5_ASAP7_75t_L g1670 ( 
.A(n_1365),
.Y(n_1670)
);

BUFx4f_ASAP7_75t_L g1671 ( 
.A(n_1372),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1366),
.Y(n_1672)
);

NAND2x1p5_ASAP7_75t_L g1673 ( 
.A(n_1374),
.B(n_64),
.Y(n_1673)
);

INVx4_ASAP7_75t_L g1674 ( 
.A(n_1368),
.Y(n_1674)
);

NOR2xp67_ASAP7_75t_L g1675 ( 
.A(n_1371),
.B(n_340),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1197),
.B(n_64),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1184),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1256),
.B(n_65),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1270),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1271),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1680)
);

INVx5_ASAP7_75t_L g1681 ( 
.A(n_1214),
.Y(n_1681)
);

CKINVDCx20_ASAP7_75t_R g1682 ( 
.A(n_1319),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1256),
.B(n_66),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1242),
.Y(n_1684)
);

INVx3_ASAP7_75t_L g1685 ( 
.A(n_1243),
.Y(n_1685)
);

NOR2x2_ASAP7_75t_L g1686 ( 
.A(n_1178),
.B(n_67),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1319),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1197),
.B(n_69),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1191),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1319),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1191),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1197),
.B(n_69),
.Y(n_1692)
);

A2O1A1Ixp33_ASAP7_75t_L g1693 ( 
.A1(n_1184),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1606),
.B(n_71),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1438),
.B(n_73),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1562),
.A2(n_76),
.B(n_74),
.C(n_75),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_SL g1697 ( 
.A(n_1451),
.B(n_74),
.Y(n_1697)
);

BUFx6f_ASAP7_75t_L g1698 ( 
.A(n_1467),
.Y(n_1698)
);

BUFx6f_ASAP7_75t_L g1699 ( 
.A(n_1467),
.Y(n_1699)
);

O2A1O1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1447),
.A2(n_78),
.B(n_75),
.C(n_77),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1429),
.A2(n_80),
.B1(n_77),
.B2(n_79),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1461),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1481),
.B(n_80),
.Y(n_1703)
);

OAI22x1_ASAP7_75t_L g1704 ( 
.A1(n_1443),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1440),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1612),
.B(n_83),
.Y(n_1706)
);

A2O1A1Ixp33_ASAP7_75t_L g1707 ( 
.A1(n_1614),
.A2(n_87),
.B(n_84),
.C(n_86),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1514),
.B(n_84),
.Y(n_1708)
);

NOR2x1_ASAP7_75t_L g1709 ( 
.A(n_1530),
.B(n_86),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1616),
.B(n_87),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1568),
.A2(n_1578),
.B1(n_1610),
.B2(n_1586),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1442),
.B(n_88),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1467),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1519),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1451),
.B(n_88),
.Y(n_1715)
);

INVxp67_ASAP7_75t_SL g1716 ( 
.A(n_1416),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1630),
.B(n_89),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1548),
.A2(n_364),
.B(n_361),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1533),
.B(n_89),
.Y(n_1719)
);

A2O1A1Ixp33_ASAP7_75t_L g1720 ( 
.A1(n_1676),
.A2(n_93),
.B(n_90),
.C(n_92),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1432),
.B(n_90),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1521),
.Y(n_1722)
);

A2O1A1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1688),
.A2(n_95),
.B(n_92),
.C(n_94),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1639),
.B(n_95),
.Y(n_1724)
);

O2A1O1Ixp33_ASAP7_75t_L g1725 ( 
.A1(n_1486),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_1725)
);

AO21x2_ASAP7_75t_L g1726 ( 
.A1(n_1669),
.A2(n_367),
.B(n_366),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1525),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1451),
.B(n_99),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1648),
.B(n_99),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1575),
.B(n_102),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1536),
.B(n_1527),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1478),
.B(n_103),
.Y(n_1732)
);

OAI22x1_ASAP7_75t_L g1733 ( 
.A1(n_1443),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1468),
.B(n_104),
.Y(n_1734)
);

AOI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1573),
.A2(n_371),
.B(n_369),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1661),
.A2(n_373),
.B(n_372),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1661),
.A2(n_378),
.B(n_375),
.Y(n_1737)
);

BUFx12f_ASAP7_75t_L g1738 ( 
.A(n_1538),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1428),
.A2(n_1506),
.B1(n_1437),
.B2(n_1501),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1468),
.B(n_106),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1563),
.A2(n_1564),
.B(n_1433),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1431),
.A2(n_380),
.B(n_379),
.Y(n_1742)
);

INVx3_ASAP7_75t_SL g1743 ( 
.A(n_1686),
.Y(n_1743)
);

AOI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1436),
.A2(n_383),
.B(n_381),
.Y(n_1744)
);

NAND3xp33_ASAP7_75t_SL g1745 ( 
.A(n_1448),
.B(n_106),
.C(n_107),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1681),
.B(n_107),
.Y(n_1746)
);

BUFx2_ASAP7_75t_L g1747 ( 
.A(n_1530),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1413),
.Y(n_1748)
);

O2A1O1Ixp33_ASAP7_75t_L g1749 ( 
.A1(n_1678),
.A2(n_113),
.B(n_108),
.C(n_112),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1450),
.A2(n_389),
.B(n_386),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1420),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1471),
.B(n_114),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1479),
.B(n_115),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1457),
.A2(n_397),
.B(n_393),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1421),
.Y(n_1755)
);

INVx4_ASAP7_75t_L g1756 ( 
.A(n_1681),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1445),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1452),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1454),
.B(n_116),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1460),
.A2(n_1466),
.B(n_1463),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1459),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1681),
.B(n_117),
.Y(n_1762)
);

INVx4_ASAP7_75t_L g1763 ( 
.A(n_1493),
.Y(n_1763)
);

BUFx2_ASAP7_75t_L g1764 ( 
.A(n_1427),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1615),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_1765)
);

AO21x1_ASAP7_75t_L g1766 ( 
.A1(n_1673),
.A2(n_403),
.B(n_401),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1550),
.B(n_118),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1474),
.B(n_119),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1684),
.B(n_120),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1476),
.B(n_123),
.Y(n_1770)
);

INVx4_ASAP7_75t_L g1771 ( 
.A(n_1493),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1480),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1437),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1677),
.Y(n_1774)
);

O2A1O1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1683),
.A2(n_129),
.B(n_126),
.C(n_127),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1528),
.B(n_127),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1570),
.B(n_129),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1602),
.B(n_130),
.Y(n_1778)
);

NAND2x1p5_ASAP7_75t_L g1779 ( 
.A(n_1493),
.B(n_1545),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1422),
.Y(n_1780)
);

O2A1O1Ixp33_ASAP7_75t_L g1781 ( 
.A1(n_1592),
.A2(n_133),
.B(n_131),
.C(n_132),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1637),
.B(n_132),
.Y(n_1782)
);

OAI21x1_ASAP7_75t_L g1783 ( 
.A1(n_1609),
.A2(n_409),
.B(n_408),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1535),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1494),
.B(n_134),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_R g1786 ( 
.A(n_1682),
.B(n_135),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1487),
.B(n_136),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1415),
.B(n_137),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1415),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_1789)
);

A2O1A1Ixp33_ASAP7_75t_L g1790 ( 
.A1(n_1659),
.A2(n_141),
.B(n_138),
.C(n_140),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1434),
.B(n_141),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1482),
.B(n_142),
.Y(n_1792)
);

OR2x2_ASAP7_75t_SL g1793 ( 
.A(n_1489),
.B(n_142),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_SL g1794 ( 
.A1(n_1419),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_1794)
);

OAI221xp5_ASAP7_75t_L g1795 ( 
.A1(n_1423),
.A2(n_145),
.B1(n_146),
.B2(n_149),
.C(n_150),
.Y(n_1795)
);

O2A1O1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1692),
.A2(n_1693),
.B(n_1470),
.C(n_1472),
.Y(n_1796)
);

AOI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1515),
.A2(n_411),
.B(n_410),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1446),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1515),
.A2(n_413),
.B(n_412),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1531),
.B(n_152),
.Y(n_1800)
);

O2A1O1Ixp33_ASAP7_75t_L g1801 ( 
.A1(n_1618),
.A2(n_155),
.B(n_153),
.C(n_154),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1544),
.B(n_154),
.Y(n_1802)
);

BUFx2_ASAP7_75t_L g1803 ( 
.A(n_1553),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1515),
.A2(n_419),
.B(n_415),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1571),
.B(n_1574),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1512),
.B(n_156),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1480),
.B(n_157),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1552),
.B(n_157),
.Y(n_1808)
);

BUFx2_ASAP7_75t_L g1809 ( 
.A(n_1554),
.Y(n_1809)
);

AO22x1_ASAP7_75t_L g1810 ( 
.A1(n_1687),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1685),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_SL g1812 ( 
.A1(n_1490),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_1812)
);

BUFx12f_ASAP7_75t_L g1813 ( 
.A(n_1417),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1526),
.B(n_162),
.Y(n_1814)
);

OAI21xp33_ASAP7_75t_L g1815 ( 
.A1(n_1541),
.A2(n_162),
.B(n_163),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1680),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1505),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_1817)
);

NAND2x1p5_ASAP7_75t_L g1818 ( 
.A(n_1545),
.B(n_167),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1495),
.B(n_168),
.Y(n_1819)
);

NOR2xp33_ASAP7_75t_R g1820 ( 
.A(n_1690),
.B(n_169),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1484),
.B(n_1654),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1584),
.B(n_169),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_SL g1823 ( 
.A(n_1455),
.B(n_170),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1642),
.Y(n_1824)
);

A2O1A1Ixp33_ASAP7_75t_L g1825 ( 
.A1(n_1621),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_1825)
);

CKINVDCx8_ASAP7_75t_R g1826 ( 
.A(n_1444),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1522),
.A2(n_422),
.B(n_421),
.Y(n_1827)
);

A2O1A1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1620),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_1828)
);

BUFx12f_ASAP7_75t_L g1829 ( 
.A(n_1435),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1508),
.B(n_174),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1458),
.B(n_174),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1458),
.B(n_177),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1465),
.Y(n_1833)
);

O2A1O1Ixp33_ASAP7_75t_L g1834 ( 
.A1(n_1658),
.A2(n_179),
.B(n_177),
.C(n_178),
.Y(n_1834)
);

BUFx12f_ASAP7_75t_L g1835 ( 
.A(n_1679),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_R g1836 ( 
.A(n_1444),
.B(n_178),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1644),
.B(n_180),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1643),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1549),
.B(n_182),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1680),
.A2(n_183),
.B1(n_185),
.B2(n_187),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1488),
.B(n_185),
.Y(n_1841)
);

BUFx6f_ASAP7_75t_L g1842 ( 
.A(n_1414),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1551),
.B(n_187),
.Y(n_1843)
);

INVxp67_ASAP7_75t_L g1844 ( 
.A(n_1651),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1588),
.B(n_188),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1655),
.A2(n_188),
.B1(n_189),
.B2(n_191),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1566),
.B(n_191),
.Y(n_1847)
);

BUFx2_ASAP7_75t_L g1848 ( 
.A(n_1424),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1492),
.B(n_192),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1509),
.Y(n_1850)
);

AOI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1522),
.A2(n_426),
.B(n_425),
.Y(n_1851)
);

A2O1A1Ixp33_ASAP7_75t_L g1852 ( 
.A1(n_1569),
.A2(n_192),
.B(n_193),
.C(n_194),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1522),
.A2(n_428),
.B(n_427),
.Y(n_1853)
);

NOR2xp67_ASAP7_75t_SL g1854 ( 
.A(n_1561),
.B(n_193),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1655),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_1855)
);

A2O1A1Ixp33_ASAP7_75t_L g1856 ( 
.A1(n_1569),
.A2(n_196),
.B(n_197),
.C(n_198),
.Y(n_1856)
);

A2O1A1Ixp33_ASAP7_75t_L g1857 ( 
.A1(n_1556),
.A2(n_199),
.B(n_200),
.C(n_201),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1492),
.B(n_199),
.Y(n_1858)
);

A2O1A1Ixp33_ASAP7_75t_L g1859 ( 
.A1(n_1556),
.A2(n_1597),
.B(n_1641),
.C(n_1645),
.Y(n_1859)
);

NOR3xp33_ASAP7_75t_SL g1860 ( 
.A(n_1635),
.B(n_200),
.C(n_202),
.Y(n_1860)
);

O2A1O1Ixp33_ASAP7_75t_L g1861 ( 
.A1(n_1426),
.A2(n_202),
.B(n_203),
.C(n_204),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1496),
.B(n_203),
.Y(n_1862)
);

AOI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1534),
.A2(n_205),
.B1(n_206),
.B2(n_209),
.Y(n_1863)
);

AOI21x1_ASAP7_75t_L g1864 ( 
.A1(n_1511),
.A2(n_430),
.B(n_429),
.Y(n_1864)
);

OAI21x1_ASAP7_75t_L g1865 ( 
.A1(n_1675),
.A2(n_436),
.B(n_434),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1588),
.B(n_205),
.Y(n_1866)
);

INVxp67_ASAP7_75t_L g1867 ( 
.A(n_1651),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1477),
.B(n_212),
.Y(n_1868)
);

OAI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1608),
.A2(n_213),
.B(n_215),
.Y(n_1869)
);

BUFx12f_ASAP7_75t_L g1870 ( 
.A(n_1453),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_SL g1871 ( 
.A(n_1657),
.B(n_213),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1581),
.Y(n_1872)
);

OAI21xp33_ASAP7_75t_SL g1873 ( 
.A1(n_1668),
.A2(n_216),
.B(n_217),
.Y(n_1873)
);

AOI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1524),
.A2(n_438),
.B(n_437),
.Y(n_1874)
);

INVx2_ASAP7_75t_SL g1875 ( 
.A(n_1449),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1583),
.Y(n_1876)
);

A2O1A1Ixp33_ASAP7_75t_L g1877 ( 
.A1(n_1626),
.A2(n_216),
.B(n_217),
.C(n_218),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1500),
.B(n_1475),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1500),
.B(n_218),
.Y(n_1879)
);

A2O1A1Ixp33_ASAP7_75t_L g1880 ( 
.A1(n_1608),
.A2(n_219),
.B(n_220),
.C(n_221),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1668),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_1881)
);

INVx4_ASAP7_75t_L g1882 ( 
.A(n_1418),
.Y(n_1882)
);

AOI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1505),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1469),
.B(n_229),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1667),
.Y(n_1885)
);

BUFx2_ASAP7_75t_L g1886 ( 
.A(n_1507),
.Y(n_1886)
);

HB1xp67_ASAP7_75t_L g1887 ( 
.A(n_1603),
.Y(n_1887)
);

OAI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1496),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_SL g1889 ( 
.A(n_1595),
.B(n_230),
.Y(n_1889)
);

BUFx8_ASAP7_75t_SL g1890 ( 
.A(n_1502),
.Y(n_1890)
);

AOI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1613),
.A2(n_442),
.B(n_440),
.Y(n_1891)
);

AOI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1585),
.A2(n_445),
.B(n_444),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1636),
.B(n_231),
.Y(n_1893)
);

OAI221xp5_ASAP7_75t_L g1894 ( 
.A1(n_1504),
.A2(n_233),
.B1(n_234),
.B2(n_236),
.C(n_237),
.Y(n_1894)
);

BUFx6f_ASAP7_75t_L g1895 ( 
.A(n_1441),
.Y(n_1895)
);

OAI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1649),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_1896)
);

AOI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1601),
.A2(n_460),
.B(n_558),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1439),
.Y(n_1898)
);

CKINVDCx20_ASAP7_75t_R g1899 ( 
.A(n_1593),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1638),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1529),
.B(n_239),
.Y(n_1901)
);

OAI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1540),
.A2(n_240),
.B(n_242),
.Y(n_1902)
);

BUFx3_ASAP7_75t_L g1903 ( 
.A(n_1623),
.Y(n_1903)
);

BUFx6f_ASAP7_75t_L g1904 ( 
.A(n_1441),
.Y(n_1904)
);

BUFx12f_ASAP7_75t_L g1905 ( 
.A(n_1611),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1485),
.B(n_240),
.Y(n_1906)
);

INVx5_ASAP7_75t_L g1907 ( 
.A(n_1462),
.Y(n_1907)
);

AOI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1650),
.A2(n_464),
.B(n_557),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1532),
.B(n_243),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1559),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1599),
.A2(n_463),
.B(n_556),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_R g1912 ( 
.A(n_1617),
.B(n_244),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1580),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1510),
.B(n_245),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1560),
.B(n_245),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1485),
.B(n_246),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1537),
.B(n_246),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1513),
.B(n_247),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1483),
.B(n_247),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1513),
.B(n_249),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1518),
.B(n_250),
.Y(n_1921)
);

A2O1A1Ixp33_ASAP7_75t_L g1922 ( 
.A1(n_1646),
.A2(n_251),
.B(n_253),
.C(n_254),
.Y(n_1922)
);

O2A1O1Ixp33_ASAP7_75t_L g1923 ( 
.A1(n_1627),
.A2(n_251),
.B(n_253),
.C(n_256),
.Y(n_1923)
);

NAND2x1p5_ASAP7_75t_L g1924 ( 
.A(n_1671),
.B(n_257),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1663),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1520),
.B(n_257),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_1607),
.Y(n_1927)
);

A2O1A1Ixp33_ASAP7_75t_L g1928 ( 
.A1(n_1656),
.A2(n_258),
.B(n_259),
.C(n_260),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_1607),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_1611),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1516),
.B(n_260),
.Y(n_1931)
);

O2A1O1Ixp33_ASAP7_75t_L g1932 ( 
.A1(n_1664),
.A2(n_261),
.B(n_262),
.C(n_265),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_1594),
.Y(n_1933)
);

A2O1A1Ixp33_ASAP7_75t_L g1934 ( 
.A1(n_1628),
.A2(n_1665),
.B(n_1622),
.C(n_1542),
.Y(n_1934)
);

BUFx8_ASAP7_75t_L g1935 ( 
.A(n_1640),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1587),
.A2(n_477),
.B(n_547),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_R g1937 ( 
.A(n_1617),
.B(n_261),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1543),
.B(n_265),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1516),
.B(n_266),
.Y(n_1939)
);

BUFx2_ASAP7_75t_L g1940 ( 
.A(n_1662),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1587),
.A2(n_479),
.B(n_544),
.Y(n_1941)
);

BUFx4_ASAP7_75t_SL g1942 ( 
.A(n_1624),
.Y(n_1942)
);

NAND3xp33_ASAP7_75t_SL g1943 ( 
.A(n_1572),
.B(n_266),
.C(n_267),
.Y(n_1943)
);

OR2x6_ASAP7_75t_L g1944 ( 
.A(n_1539),
.B(n_268),
.Y(n_1944)
);

NOR3xp33_ASAP7_75t_SL g1945 ( 
.A(n_1634),
.B(n_268),
.C(n_269),
.Y(n_1945)
);

A2O1A1Ixp33_ASAP7_75t_L g1946 ( 
.A1(n_1546),
.A2(n_270),
.B(n_271),
.C(n_272),
.Y(n_1946)
);

O2A1O1Ixp33_ASAP7_75t_L g1947 ( 
.A1(n_1577),
.A2(n_270),
.B(n_271),
.C(n_272),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1671),
.B(n_273),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_SL g1949 ( 
.A1(n_1689),
.A2(n_483),
.B(n_543),
.Y(n_1949)
);

BUFx6f_ASAP7_75t_L g1950 ( 
.A(n_1691),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1504),
.B(n_1491),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1497),
.B(n_274),
.Y(n_1952)
);

AO22x1_ASAP7_75t_L g1953 ( 
.A1(n_1625),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1499),
.B(n_275),
.Y(n_1954)
);

O2A1O1Ixp33_ASAP7_75t_L g1955 ( 
.A1(n_1547),
.A2(n_277),
.B(n_279),
.C(n_281),
.Y(n_1955)
);

INVx3_ASAP7_75t_L g1956 ( 
.A(n_1691),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1503),
.B(n_1517),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1473),
.Y(n_1958)
);

INVxp67_ASAP7_75t_L g1959 ( 
.A(n_1523),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_SL g1960 ( 
.A(n_1473),
.B(n_281),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1543),
.B(n_282),
.Y(n_1961)
);

HB1xp67_ASAP7_75t_L g1962 ( 
.A(n_1473),
.Y(n_1962)
);

BUFx2_ASAP7_75t_L g1963 ( 
.A(n_1558),
.Y(n_1963)
);

INVx3_ASAP7_75t_L g1964 ( 
.A(n_1498),
.Y(n_1964)
);

A2O1A1Ixp33_ASAP7_75t_L g1965 ( 
.A1(n_1598),
.A2(n_283),
.B(n_285),
.C(n_286),
.Y(n_1965)
);

OAI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1647),
.A2(n_283),
.B1(n_285),
.B2(n_286),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1498),
.B(n_288),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1631),
.B(n_288),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1633),
.B(n_289),
.Y(n_1969)
);

BUFx6f_ASAP7_75t_SL g1970 ( 
.A(n_1619),
.Y(n_1970)
);

A2O1A1Ixp33_ASAP7_75t_L g1971 ( 
.A1(n_1598),
.A2(n_291),
.B(n_292),
.C(n_293),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1633),
.B(n_294),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_SL g1973 ( 
.A(n_1660),
.B(n_494),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1629),
.B(n_294),
.Y(n_1974)
);

INVx4_ASAP7_75t_L g1975 ( 
.A(n_1498),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1579),
.B(n_295),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1576),
.B(n_295),
.Y(n_1977)
);

AOI21xp5_ASAP7_75t_L g1978 ( 
.A1(n_1425),
.A2(n_493),
.B(n_536),
.Y(n_1978)
);

O2A1O1Ixp33_ASAP7_75t_L g1979 ( 
.A1(n_1596),
.A2(n_296),
.B(n_297),
.C(n_298),
.Y(n_1979)
);

BUFx4f_ASAP7_75t_L g1980 ( 
.A(n_1632),
.Y(n_1980)
);

BUFx3_ASAP7_75t_L g1981 ( 
.A(n_1623),
.Y(n_1981)
);

INVx4_ASAP7_75t_L g1982 ( 
.A(n_1557),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1591),
.B(n_300),
.Y(n_1983)
);

NOR2xp33_ASAP7_75t_R g1984 ( 
.A(n_1594),
.B(n_301),
.Y(n_1984)
);

HB1xp67_ASAP7_75t_L g1985 ( 
.A(n_1555),
.Y(n_1985)
);

INVx2_ASAP7_75t_SL g1986 ( 
.A(n_1590),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1660),
.A2(n_498),
.B(n_535),
.Y(n_1987)
);

OR2x6_ASAP7_75t_L g1988 ( 
.A(n_1600),
.B(n_302),
.Y(n_1988)
);

BUFx8_ASAP7_75t_L g1989 ( 
.A(n_1652),
.Y(n_1989)
);

O2A1O1Ixp33_ASAP7_75t_L g1990 ( 
.A1(n_1565),
.A2(n_303),
.B(n_304),
.C(n_305),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1653),
.B(n_1589),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1605),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1558),
.B(n_303),
.Y(n_1993)
);

NOR2xp33_ASAP7_75t_L g1994 ( 
.A(n_1430),
.B(n_304),
.Y(n_1994)
);

O2A1O1Ixp33_ASAP7_75t_L g1995 ( 
.A1(n_1590),
.A2(n_449),
.B(n_450),
.C(n_454),
.Y(n_1995)
);

O2A1O1Ixp33_ASAP7_75t_L g1996 ( 
.A1(n_1666),
.A2(n_468),
.B(n_470),
.C(n_472),
.Y(n_1996)
);

OAI21x1_ASAP7_75t_L g1997 ( 
.A1(n_1582),
.A2(n_475),
.B(n_480),
.Y(n_1997)
);

A2O1A1Ixp33_ASAP7_75t_L g1998 ( 
.A1(n_1604),
.A2(n_482),
.B(n_484),
.C(n_489),
.Y(n_1998)
);

OAI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1557),
.A2(n_495),
.B1(n_499),
.B2(n_502),
.Y(n_1999)
);

AOI21xp5_ASAP7_75t_L g2000 ( 
.A1(n_1674),
.A2(n_510),
.B(n_511),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1567),
.B(n_514),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1670),
.B(n_516),
.Y(n_2002)
);

AND2x2_ASAP7_75t_SL g2003 ( 
.A(n_1672),
.B(n_524),
.Y(n_2003)
);

AOI22xp33_ASAP7_75t_L g2004 ( 
.A1(n_1670),
.A2(n_525),
.B1(n_527),
.B2(n_528),
.Y(n_2004)
);

AOI21xp5_ASAP7_75t_L g2005 ( 
.A1(n_1672),
.A2(n_530),
.B(n_559),
.Y(n_2005)
);

OAI22x1_ASAP7_75t_L g2006 ( 
.A1(n_1443),
.A2(n_1680),
.B1(n_1242),
.B2(n_1505),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1606),
.B(n_1197),
.Y(n_2007)
);

INVxp33_ASAP7_75t_SL g2008 ( 
.A(n_1416),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_1440),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1464),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1606),
.B(n_1112),
.Y(n_2011)
);

BUFx4f_ASAP7_75t_L g2012 ( 
.A(n_1417),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1606),
.B(n_1112),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1519),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1519),
.Y(n_2015)
);

INVx5_ASAP7_75t_L g2016 ( 
.A(n_1467),
.Y(n_2016)
);

OAI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_1438),
.A2(n_1612),
.B1(n_1616),
.B2(n_1614),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1606),
.B(n_1197),
.Y(n_2018)
);

AOI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_1438),
.A2(n_1137),
.B(n_1456),
.Y(n_2019)
);

AOI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1438),
.A2(n_1137),
.B(n_1456),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1606),
.B(n_1197),
.Y(n_2021)
);

CKINVDCx14_ASAP7_75t_R g2022 ( 
.A(n_1682),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1438),
.B(n_1562),
.Y(n_2023)
);

BUFx12f_ASAP7_75t_L g2024 ( 
.A(n_1461),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1606),
.B(n_1112),
.Y(n_2025)
);

BUFx2_ASAP7_75t_L g2026 ( 
.A(n_1440),
.Y(n_2026)
);

OAI22xp5_ASAP7_75t_SL g2027 ( 
.A1(n_1437),
.A2(n_1185),
.B1(n_1005),
.B2(n_1003),
.Y(n_2027)
);

INVx4_ASAP7_75t_L g2028 ( 
.A(n_1779),
.Y(n_2028)
);

BUFx10_ASAP7_75t_L g2029 ( 
.A(n_1970),
.Y(n_2029)
);

BUFx2_ASAP7_75t_L g2030 ( 
.A(n_1747),
.Y(n_2030)
);

AOI22x1_ASAP7_75t_L g2031 ( 
.A1(n_1741),
.A2(n_1760),
.B1(n_2006),
.B2(n_1911),
.Y(n_2031)
);

INVx4_ASAP7_75t_L g2032 ( 
.A(n_1779),
.Y(n_2032)
);

INVx1_ASAP7_75t_SL g2033 ( 
.A(n_2023),
.Y(n_2033)
);

CKINVDCx6p67_ASAP7_75t_R g2034 ( 
.A(n_1813),
.Y(n_2034)
);

OR2x6_ASAP7_75t_L g2035 ( 
.A(n_1944),
.B(n_2017),
.Y(n_2035)
);

INVx6_ASAP7_75t_SL g2036 ( 
.A(n_1988),
.Y(n_2036)
);

INVx4_ASAP7_75t_L g2037 ( 
.A(n_1870),
.Y(n_2037)
);

BUFx4f_ASAP7_75t_SL g2038 ( 
.A(n_1829),
.Y(n_2038)
);

BUFx8_ASAP7_75t_SL g2039 ( 
.A(n_1738),
.Y(n_2039)
);

BUFx8_ASAP7_75t_L g2040 ( 
.A(n_1835),
.Y(n_2040)
);

AO21x2_ASAP7_75t_L g2041 ( 
.A1(n_1859),
.A2(n_1726),
.B(n_1934),
.Y(n_2041)
);

AOI22x1_ASAP7_75t_L g2042 ( 
.A1(n_1742),
.A2(n_1744),
.B1(n_1754),
.B2(n_1750),
.Y(n_2042)
);

BUFx12f_ASAP7_75t_L g2043 ( 
.A(n_2024),
.Y(n_2043)
);

AO21x2_ASAP7_75t_L g2044 ( 
.A1(n_1726),
.A2(n_1961),
.B(n_1938),
.Y(n_2044)
);

AO21x1_ASAP7_75t_L g2045 ( 
.A1(n_1765),
.A2(n_2017),
.B(n_1855),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1838),
.Y(n_2046)
);

AO21x2_ASAP7_75t_L g2047 ( 
.A1(n_1938),
.A2(n_1961),
.B(n_1800),
.Y(n_2047)
);

INVx1_ASAP7_75t_SL g2048 ( 
.A(n_1940),
.Y(n_2048)
);

HB1xp67_ASAP7_75t_L g2049 ( 
.A(n_1711),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_1942),
.Y(n_2050)
);

NOR2xp67_ASAP7_75t_SL g2051 ( 
.A(n_1826),
.B(n_1907),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2011),
.B(n_2013),
.Y(n_2052)
);

BUFx3_ASAP7_75t_L g2053 ( 
.A(n_2016),
.Y(n_2053)
);

AO21x1_ASAP7_75t_L g2054 ( 
.A1(n_1765),
.A2(n_1855),
.B(n_1846),
.Y(n_2054)
);

NAND3xp33_ASAP7_75t_SL g2055 ( 
.A(n_1912),
.B(n_1937),
.C(n_1984),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1714),
.Y(n_2056)
);

INVx4_ASAP7_75t_L g2057 ( 
.A(n_2016),
.Y(n_2057)
);

AO21x2_ASAP7_75t_L g2058 ( 
.A1(n_1800),
.A2(n_1864),
.B(n_1869),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1722),
.Y(n_2059)
);

BUFx12f_ASAP7_75t_L g2060 ( 
.A(n_1702),
.Y(n_2060)
);

AO21x2_ASAP7_75t_L g2061 ( 
.A1(n_1869),
.A2(n_1825),
.B(n_1711),
.Y(n_2061)
);

HB1xp67_ASAP7_75t_L g2062 ( 
.A(n_2016),
.Y(n_2062)
);

INVx2_ASAP7_75t_SL g2063 ( 
.A(n_2012),
.Y(n_2063)
);

OAI21x1_ASAP7_75t_L g2064 ( 
.A1(n_1956),
.A2(n_1964),
.B(n_1799),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_L g2065 ( 
.A(n_2008),
.B(n_2025),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1951),
.B(n_1748),
.Y(n_2066)
);

CKINVDCx12_ASAP7_75t_R g2067 ( 
.A(n_1988),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1925),
.Y(n_2068)
);

BUFx3_ASAP7_75t_L g2069 ( 
.A(n_1848),
.Y(n_2069)
);

OAI21x1_ASAP7_75t_L g2070 ( 
.A1(n_1797),
.A2(n_1827),
.B(n_1804),
.Y(n_2070)
);

INVx5_ASAP7_75t_L g2071 ( 
.A(n_1699),
.Y(n_2071)
);

OAI21x1_ASAP7_75t_L g2072 ( 
.A1(n_1851),
.A2(n_1874),
.B(n_1853),
.Y(n_2072)
);

INVx2_ASAP7_75t_SL g2073 ( 
.A(n_2012),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1751),
.B(n_1755),
.Y(n_2074)
);

AO21x2_ASAP7_75t_L g2075 ( 
.A1(n_1766),
.A2(n_1806),
.B(n_1993),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_1890),
.Y(n_2076)
);

OAI21x1_ASAP7_75t_SL g2077 ( 
.A1(n_1902),
.A2(n_1993),
.B(n_1717),
.Y(n_2077)
);

INVx1_ASAP7_75t_SL g2078 ( 
.A(n_1764),
.Y(n_2078)
);

HB1xp67_ASAP7_75t_L g2079 ( 
.A(n_1944),
.Y(n_2079)
);

AO21x2_ASAP7_75t_L g2080 ( 
.A1(n_1806),
.A2(n_1710),
.B(n_1717),
.Y(n_2080)
);

AOI22xp33_ASAP7_75t_SL g2081 ( 
.A1(n_1881),
.A2(n_1846),
.B1(n_1816),
.B2(n_1840),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1727),
.Y(n_2082)
);

NAND2x1p5_ASAP7_75t_L g2083 ( 
.A(n_1907),
.B(n_1763),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_2014),
.B(n_2015),
.Y(n_2084)
);

INVx4_ASAP7_75t_L g2085 ( 
.A(n_1771),
.Y(n_2085)
);

CKINVDCx16_ASAP7_75t_R g2086 ( 
.A(n_1836),
.Y(n_2086)
);

INVx3_ASAP7_75t_L g2087 ( 
.A(n_1771),
.Y(n_2087)
);

INVx2_ASAP7_75t_SL g2088 ( 
.A(n_1886),
.Y(n_2088)
);

OA21x2_ASAP7_75t_L g2089 ( 
.A1(n_1997),
.A2(n_1815),
.B(n_1718),
.Y(n_2089)
);

AO21x2_ASAP7_75t_L g2090 ( 
.A1(n_1710),
.A2(n_1752),
.B(n_1719),
.Y(n_2090)
);

AO21x2_ASAP7_75t_L g2091 ( 
.A1(n_1719),
.A2(n_1967),
.B(n_1960),
.Y(n_2091)
);

CKINVDCx16_ASAP7_75t_R g2092 ( 
.A(n_1786),
.Y(n_2092)
);

INVx8_ASAP7_75t_L g2093 ( 
.A(n_1944),
.Y(n_2093)
);

INVx8_ASAP7_75t_L g2094 ( 
.A(n_1988),
.Y(n_2094)
);

BUFx3_ASAP7_75t_L g2095 ( 
.A(n_1903),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1757),
.Y(n_2096)
);

INVx6_ASAP7_75t_L g2097 ( 
.A(n_1989),
.Y(n_2097)
);

OAI21x1_ASAP7_75t_L g2098 ( 
.A1(n_1936),
.A2(n_1941),
.B(n_2005),
.Y(n_2098)
);

CKINVDCx20_ASAP7_75t_R g2099 ( 
.A(n_2022),
.Y(n_2099)
);

HB1xp67_ASAP7_75t_L g2100 ( 
.A(n_1969),
.Y(n_2100)
);

BUFx3_ASAP7_75t_L g2101 ( 
.A(n_1981),
.Y(n_2101)
);

NAND2x1p5_ASAP7_75t_L g2102 ( 
.A(n_1907),
.B(n_1746),
.Y(n_2102)
);

INVx6_ASAP7_75t_SL g2103 ( 
.A(n_1746),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1731),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1805),
.B(n_1809),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1758),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1774),
.Y(n_2107)
);

OR2x6_ASAP7_75t_L g2108 ( 
.A(n_1818),
.B(n_1915),
.Y(n_2108)
);

OAI21xp5_ASAP7_75t_L g2109 ( 
.A1(n_1796),
.A2(n_1695),
.B(n_1957),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_1705),
.B(n_2026),
.Y(n_2110)
);

AND2x4_ASAP7_75t_L g2111 ( 
.A(n_1821),
.B(n_1780),
.Y(n_2111)
);

CKINVDCx16_ASAP7_75t_R g2112 ( 
.A(n_2027),
.Y(n_2112)
);

INVx3_ASAP7_75t_SL g2113 ( 
.A(n_1762),
.Y(n_2113)
);

INVx1_ASAP7_75t_SL g2114 ( 
.A(n_1761),
.Y(n_2114)
);

INVx1_ASAP7_75t_SL g2115 ( 
.A(n_1784),
.Y(n_2115)
);

AO21x2_ASAP7_75t_L g2116 ( 
.A1(n_1759),
.A2(n_1770),
.B(n_1768),
.Y(n_2116)
);

INVxp67_ASAP7_75t_SL g2117 ( 
.A(n_1842),
.Y(n_2117)
);

AO21x2_ASAP7_75t_L g2118 ( 
.A1(n_1785),
.A2(n_1972),
.B(n_1968),
.Y(n_2118)
);

INVx4_ASAP7_75t_L g2119 ( 
.A(n_1762),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1885),
.B(n_1824),
.Y(n_2120)
);

AOI22xp33_ASAP7_75t_L g2121 ( 
.A1(n_1732),
.A2(n_1716),
.B1(n_1795),
.B2(n_1753),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_1782),
.B(n_2009),
.Y(n_2122)
);

BUFx5_ASAP7_75t_L g2123 ( 
.A(n_2003),
.Y(n_2123)
);

AOI21xp5_ASAP7_75t_L g2124 ( 
.A1(n_1839),
.A2(n_1843),
.B(n_1952),
.Y(n_2124)
);

INVx2_ASAP7_75t_SL g2125 ( 
.A(n_1803),
.Y(n_2125)
);

OAI21xp5_ASAP7_75t_L g2126 ( 
.A1(n_1706),
.A2(n_1808),
.B(n_1996),
.Y(n_2126)
);

AOI22xp5_ASAP7_75t_L g2127 ( 
.A1(n_2007),
.A2(n_2018),
.B1(n_2021),
.B2(n_1739),
.Y(n_2127)
);

AND2x4_ASAP7_75t_L g2128 ( 
.A(n_1872),
.B(n_1876),
.Y(n_2128)
);

INVx4_ASAP7_75t_SL g2129 ( 
.A(n_1699),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_1939),
.B(n_1703),
.Y(n_2130)
);

INVx3_ASAP7_75t_L g2131 ( 
.A(n_1882),
.Y(n_2131)
);

OAI21x1_ASAP7_75t_L g2132 ( 
.A1(n_1987),
.A2(n_1978),
.B(n_2000),
.Y(n_2132)
);

INVx4_ASAP7_75t_L g2133 ( 
.A(n_1970),
.Y(n_2133)
);

OAI21x1_ASAP7_75t_L g2134 ( 
.A1(n_1908),
.A2(n_1735),
.B(n_1736),
.Y(n_2134)
);

OAI21x1_ASAP7_75t_L g2135 ( 
.A1(n_1737),
.A2(n_1891),
.B(n_1892),
.Y(n_2135)
);

OAI21x1_ASAP7_75t_L g2136 ( 
.A1(n_1897),
.A2(n_1999),
.B(n_1949),
.Y(n_2136)
);

BUFx3_ASAP7_75t_L g2137 ( 
.A(n_1713),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1900),
.Y(n_2138)
);

INVx2_ASAP7_75t_SL g2139 ( 
.A(n_1980),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1808),
.Y(n_2140)
);

INVx2_ASAP7_75t_SL g2141 ( 
.A(n_1980),
.Y(n_2141)
);

INVx2_ASAP7_75t_SL g2142 ( 
.A(n_1915),
.Y(n_2142)
);

NAND2x1p5_ASAP7_75t_L g2143 ( 
.A(n_1882),
.B(n_1975),
.Y(n_2143)
);

BUFx3_ASAP7_75t_L g2144 ( 
.A(n_1713),
.Y(n_2144)
);

NAND2x1p5_ASAP7_75t_L g2145 ( 
.A(n_1975),
.B(n_1963),
.Y(n_2145)
);

BUFx4f_ASAP7_75t_SL g2146 ( 
.A(n_1905),
.Y(n_2146)
);

INVx2_ASAP7_75t_SL g2147 ( 
.A(n_1833),
.Y(n_2147)
);

BUFx8_ASAP7_75t_L g2148 ( 
.A(n_1875),
.Y(n_2148)
);

OAI21x1_ASAP7_75t_L g2149 ( 
.A1(n_1999),
.A2(n_1995),
.B(n_2002),
.Y(n_2149)
);

OR2x6_ASAP7_75t_L g2150 ( 
.A(n_1818),
.B(n_1924),
.Y(n_2150)
);

BUFx3_ASAP7_75t_L g2151 ( 
.A(n_1842),
.Y(n_2151)
);

INVxp67_ASAP7_75t_SL g2152 ( 
.A(n_1842),
.Y(n_2152)
);

BUFx8_ASAP7_75t_L g2153 ( 
.A(n_1791),
.Y(n_2153)
);

HB1xp67_ASAP7_75t_L g2154 ( 
.A(n_1969),
.Y(n_2154)
);

BUFx2_ASAP7_75t_SL g2155 ( 
.A(n_1792),
.Y(n_2155)
);

AO21x2_ASAP7_75t_L g2156 ( 
.A1(n_1954),
.A2(n_1971),
.B(n_1965),
.Y(n_2156)
);

OAI21x1_ASAP7_75t_L g2157 ( 
.A1(n_1811),
.A2(n_1962),
.B(n_1992),
.Y(n_2157)
);

BUFx2_ASAP7_75t_SL g2158 ( 
.A(n_1792),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_1721),
.B(n_1959),
.Y(n_2159)
);

BUFx2_ASAP7_75t_L g2160 ( 
.A(n_1844),
.Y(n_2160)
);

AO21x2_ASAP7_75t_L g2161 ( 
.A1(n_1893),
.A2(n_1723),
.B(n_1720),
.Y(n_2161)
);

NOR2xp67_ASAP7_75t_L g2162 ( 
.A(n_1867),
.B(n_1986),
.Y(n_2162)
);

CKINVDCx11_ASAP7_75t_R g2163 ( 
.A(n_1743),
.Y(n_2163)
);

CKINVDCx20_ASAP7_75t_R g2164 ( 
.A(n_1820),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1850),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1913),
.B(n_1910),
.Y(n_2166)
);

OAI21xp5_ASAP7_75t_L g2167 ( 
.A1(n_1787),
.A2(n_1873),
.B(n_1819),
.Y(n_2167)
);

NAND2x1p5_ASAP7_75t_L g2168 ( 
.A(n_1895),
.B(n_1904),
.Y(n_2168)
);

CKINVDCx6p67_ASAP7_75t_R g2169 ( 
.A(n_1899),
.Y(n_2169)
);

NAND2x1p5_ASAP7_75t_L g2170 ( 
.A(n_1895),
.B(n_1904),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1837),
.Y(n_2171)
);

INVx2_ASAP7_75t_SL g2172 ( 
.A(n_1989),
.Y(n_2172)
);

INVx3_ASAP7_75t_L g2173 ( 
.A(n_1982),
.Y(n_2173)
);

OA21x2_ASAP7_75t_L g2174 ( 
.A1(n_1696),
.A2(n_1922),
.B(n_1880),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1888),
.Y(n_2175)
);

AO21x2_ASAP7_75t_L g2176 ( 
.A1(n_1707),
.A2(n_1790),
.B(n_1946),
.Y(n_2176)
);

BUFx10_ASAP7_75t_L g2177 ( 
.A(n_1778),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_1847),
.B(n_1814),
.Y(n_2178)
);

AO21x1_ASAP7_75t_L g2179 ( 
.A1(n_1816),
.A2(n_1840),
.B(n_1896),
.Y(n_2179)
);

INVx3_ASAP7_75t_SL g2180 ( 
.A(n_1933),
.Y(n_2180)
);

INVx5_ASAP7_75t_SL g2181 ( 
.A(n_1950),
.Y(n_2181)
);

CKINVDCx11_ASAP7_75t_R g2182 ( 
.A(n_1772),
.Y(n_2182)
);

AO21x1_ASAP7_75t_L g2183 ( 
.A1(n_1896),
.A2(n_1973),
.B(n_1966),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1950),
.Y(n_2184)
);

INVx2_ASAP7_75t_SL g2185 ( 
.A(n_1898),
.Y(n_2185)
);

NAND2x1p5_ASAP7_75t_L g2186 ( 
.A(n_1950),
.B(n_1958),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1849),
.Y(n_2187)
);

INVx4_ASAP7_75t_L g2188 ( 
.A(n_1958),
.Y(n_2188)
);

INVx3_ASAP7_75t_L g2189 ( 
.A(n_1982),
.Y(n_2189)
);

INVx3_ASAP7_75t_L g2190 ( 
.A(n_2010),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1849),
.Y(n_2191)
);

INVx8_ASAP7_75t_L g2192 ( 
.A(n_1724),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1858),
.Y(n_2193)
);

AOI22x1_ASAP7_75t_L g2194 ( 
.A1(n_1704),
.A2(n_1733),
.B1(n_1868),
.B2(n_1887),
.Y(n_2194)
);

OA21x2_ASAP7_75t_L g2195 ( 
.A1(n_1877),
.A2(n_1928),
.B(n_1998),
.Y(n_2195)
);

INVx1_ASAP7_75t_SL g2196 ( 
.A(n_1729),
.Y(n_2196)
);

INVx3_ASAP7_75t_L g2197 ( 
.A(n_1935),
.Y(n_2197)
);

NAND2x1p5_ASAP7_75t_L g2198 ( 
.A(n_1709),
.B(n_1878),
.Y(n_2198)
);

AO21x2_ASAP7_75t_L g2199 ( 
.A1(n_1841),
.A2(n_1856),
.B(n_1852),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1976),
.B(n_1917),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_1802),
.B(n_1767),
.Y(n_2201)
);

OAI21xp5_ASAP7_75t_L g2202 ( 
.A1(n_1858),
.A2(n_1862),
.B(n_1807),
.Y(n_2202)
);

AND2x4_ASAP7_75t_L g2203 ( 
.A(n_1845),
.B(n_1866),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1862),
.Y(n_2204)
);

HB1xp67_ASAP7_75t_L g2205 ( 
.A(n_1985),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1807),
.Y(n_2206)
);

OAI21x1_ASAP7_75t_L g2207 ( 
.A1(n_2004),
.A2(n_1749),
.B(n_1775),
.Y(n_2207)
);

BUFx6f_ASAP7_75t_L g2208 ( 
.A(n_1697),
.Y(n_2208)
);

INVx3_ASAP7_75t_SL g2209 ( 
.A(n_1793),
.Y(n_2209)
);

OA21x2_ASAP7_75t_L g2210 ( 
.A1(n_1857),
.A2(n_1828),
.B(n_1945),
.Y(n_2210)
);

OAI21x1_ASAP7_75t_L g2211 ( 
.A1(n_2001),
.A2(n_1801),
.B(n_1728),
.Y(n_2211)
);

AO21x2_ASAP7_75t_L g2212 ( 
.A1(n_1830),
.A2(n_1947),
.B(n_1879),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1831),
.Y(n_2213)
);

NAND2x1p5_ASAP7_75t_L g2214 ( 
.A(n_1948),
.B(n_1715),
.Y(n_2214)
);

NAND2x1p5_ASAP7_75t_L g2215 ( 
.A(n_1734),
.B(n_1740),
.Y(n_2215)
);

HB1xp67_ASAP7_75t_L g2216 ( 
.A(n_1772),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_1822),
.B(n_1777),
.Y(n_2217)
);

BUFx3_ASAP7_75t_L g2218 ( 
.A(n_1935),
.Y(n_2218)
);

INVx5_ASAP7_75t_L g2219 ( 
.A(n_1973),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1974),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_1708),
.B(n_1773),
.Y(n_2221)
);

INVx4_ASAP7_75t_L g2222 ( 
.A(n_1927),
.Y(n_2222)
);

INVx2_ASAP7_75t_SL g2223 ( 
.A(n_1788),
.Y(n_2223)
);

NOR2xp33_ASAP7_75t_L g2224 ( 
.A(n_1712),
.B(n_1991),
.Y(n_2224)
);

OAI21xp5_ASAP7_75t_L g2225 ( 
.A1(n_1725),
.A2(n_1700),
.B(n_1914),
.Y(n_2225)
);

INVx6_ASAP7_75t_SL g2226 ( 
.A(n_1854),
.Y(n_2226)
);

BUFx2_ASAP7_75t_R g2227 ( 
.A(n_1929),
.Y(n_2227)
);

OAI21x1_ASAP7_75t_L g2228 ( 
.A1(n_1932),
.A2(n_1923),
.B(n_1834),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1832),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1860),
.B(n_1930),
.Y(n_2230)
);

BUFx3_ASAP7_75t_L g2231 ( 
.A(n_1906),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1694),
.Y(n_2232)
);

OA21x2_ASAP7_75t_L g2233 ( 
.A1(n_1916),
.A2(n_1918),
.B(n_1931),
.Y(n_2233)
);

INVx3_ASAP7_75t_SL g2234 ( 
.A(n_1871),
.Y(n_2234)
);

OAI21x1_ASAP7_75t_L g2235 ( 
.A1(n_1979),
.A2(n_1861),
.B(n_1955),
.Y(n_2235)
);

BUFx2_ASAP7_75t_R g2236 ( 
.A(n_1889),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1920),
.Y(n_2237)
);

BUFx8_ASAP7_75t_SL g2238 ( 
.A(n_1953),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1789),
.Y(n_2239)
);

OAI21x1_ASAP7_75t_L g2240 ( 
.A1(n_1990),
.A2(n_1966),
.B(n_1781),
.Y(n_2240)
);

INVx2_ASAP7_75t_SL g2241 ( 
.A(n_1823),
.Y(n_2241)
);

BUFx4f_ASAP7_75t_SL g2242 ( 
.A(n_1730),
.Y(n_2242)
);

INVx4_ASAP7_75t_L g2243 ( 
.A(n_1812),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1798),
.Y(n_2244)
);

AO21x2_ASAP7_75t_L g2245 ( 
.A1(n_1943),
.A2(n_1863),
.B(n_1883),
.Y(n_2245)
);

BUFx2_ASAP7_75t_SL g2246 ( 
.A(n_1810),
.Y(n_2246)
);

OAI21x1_ASAP7_75t_L g2247 ( 
.A1(n_1817),
.A2(n_1701),
.B(n_1994),
.Y(n_2247)
);

AO21x2_ASAP7_75t_L g2248 ( 
.A1(n_1745),
.A2(n_1909),
.B(n_1901),
.Y(n_2248)
);

OAI21x1_ASAP7_75t_L g2249 ( 
.A1(n_1884),
.A2(n_1983),
.B(n_1977),
.Y(n_2249)
);

INVx3_ASAP7_75t_L g2250 ( 
.A(n_1769),
.Y(n_2250)
);

AO21x2_ASAP7_75t_L g2251 ( 
.A1(n_1894),
.A2(n_1919),
.B(n_1921),
.Y(n_2251)
);

BUFx2_ASAP7_75t_L g2252 ( 
.A(n_1776),
.Y(n_2252)
);

BUFx2_ASAP7_75t_R g2253 ( 
.A(n_1794),
.Y(n_2253)
);

AOI22x1_ASAP7_75t_L g2254 ( 
.A1(n_1926),
.A2(n_1741),
.B1(n_1760),
.B2(n_2006),
.Y(n_2254)
);

NAND2x1p5_ASAP7_75t_L g2255 ( 
.A(n_1756),
.B(n_1451),
.Y(n_2255)
);

BUFx3_ASAP7_75t_L g2256 ( 
.A(n_1779),
.Y(n_2256)
);

INVx8_ASAP7_75t_L g2257 ( 
.A(n_1870),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2023),
.B(n_2017),
.Y(n_2258)
);

NAND2x1p5_ASAP7_75t_L g2259 ( 
.A(n_1756),
.B(n_1451),
.Y(n_2259)
);

NAND2x1p5_ASAP7_75t_L g2260 ( 
.A(n_1756),
.B(n_1451),
.Y(n_2260)
);

INVx1_ASAP7_75t_SL g2261 ( 
.A(n_2023),
.Y(n_2261)
);

AO21x1_ASAP7_75t_L g2262 ( 
.A1(n_1765),
.A2(n_2017),
.B(n_1855),
.Y(n_2262)
);

HB1xp67_ASAP7_75t_L g2263 ( 
.A(n_2017),
.Y(n_2263)
);

OAI21x1_ASAP7_75t_L g2264 ( 
.A1(n_1865),
.A2(n_1783),
.B(n_1172),
.Y(n_2264)
);

OAI21x1_ASAP7_75t_L g2265 ( 
.A1(n_1865),
.A2(n_1783),
.B(n_1172),
.Y(n_2265)
);

AND2x4_ASAP7_75t_L g2266 ( 
.A(n_2023),
.B(n_1451),
.Y(n_2266)
);

BUFx3_ASAP7_75t_L g2267 ( 
.A(n_1779),
.Y(n_2267)
);

BUFx3_ASAP7_75t_L g2268 ( 
.A(n_1779),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_2011),
.B(n_1112),
.Y(n_2269)
);

AOI22x1_ASAP7_75t_L g2270 ( 
.A1(n_1741),
.A2(n_1760),
.B1(n_2006),
.B2(n_1911),
.Y(n_2270)
);

NOR2xp33_ASAP7_75t_SL g2271 ( 
.A(n_2003),
.B(n_2017),
.Y(n_2271)
);

OAI21xp5_ASAP7_75t_L g2272 ( 
.A1(n_2019),
.A2(n_2020),
.B(n_2017),
.Y(n_2272)
);

AOI22x1_ASAP7_75t_L g2273 ( 
.A1(n_1741),
.A2(n_1760),
.B1(n_2006),
.B2(n_1911),
.Y(n_2273)
);

NAND2x1p5_ASAP7_75t_L g2274 ( 
.A(n_1756),
.B(n_1451),
.Y(n_2274)
);

OAI21x1_ASAP7_75t_L g2275 ( 
.A1(n_1865),
.A2(n_1783),
.B(n_1172),
.Y(n_2275)
);

OR2x2_ASAP7_75t_L g2276 ( 
.A(n_2011),
.B(n_2013),
.Y(n_2276)
);

CKINVDCx6p67_ASAP7_75t_R g2277 ( 
.A(n_1813),
.Y(n_2277)
);

INVx2_ASAP7_75t_SL g2278 ( 
.A(n_1942),
.Y(n_2278)
);

OAI21xp5_ASAP7_75t_L g2279 ( 
.A1(n_2019),
.A2(n_2020),
.B(n_2017),
.Y(n_2279)
);

AND2x4_ASAP7_75t_L g2280 ( 
.A(n_2023),
.B(n_1451),
.Y(n_2280)
);

BUFx6f_ASAP7_75t_L g2281 ( 
.A(n_1698),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2023),
.Y(n_2282)
);

AOI21xp5_ASAP7_75t_L g2283 ( 
.A1(n_2017),
.A2(n_1137),
.B(n_1711),
.Y(n_2283)
);

OAI21x1_ASAP7_75t_L g2284 ( 
.A1(n_1865),
.A2(n_1783),
.B(n_1172),
.Y(n_2284)
);

CKINVDCx11_ASAP7_75t_R g2285 ( 
.A(n_1813),
.Y(n_2285)
);

AOI22xp33_ASAP7_75t_L g2286 ( 
.A1(n_2017),
.A2(n_1251),
.B1(n_1269),
.B2(n_1951),
.Y(n_2286)
);

AND2x4_ASAP7_75t_L g2287 ( 
.A(n_2023),
.B(n_1451),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2023),
.Y(n_2288)
);

INVx4_ASAP7_75t_L g2289 ( 
.A(n_1779),
.Y(n_2289)
);

CKINVDCx11_ASAP7_75t_R g2290 ( 
.A(n_2285),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2074),
.Y(n_2291)
);

OR2x6_ASAP7_75t_L g2292 ( 
.A(n_2035),
.B(n_2093),
.Y(n_2292)
);

BUFx6f_ASAP7_75t_L g2293 ( 
.A(n_2256),
.Y(n_2293)
);

AOI22xp5_ASAP7_75t_L g2294 ( 
.A1(n_2081),
.A2(n_2182),
.B1(n_2035),
.B2(n_2179),
.Y(n_2294)
);

AOI22xp33_ASAP7_75t_L g2295 ( 
.A1(n_2182),
.A2(n_2081),
.B1(n_2054),
.B2(n_2243),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2120),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2120),
.Y(n_2297)
);

AOI21x1_ASAP7_75t_L g2298 ( 
.A1(n_2283),
.A2(n_2077),
.B(n_2183),
.Y(n_2298)
);

HB1xp67_ASAP7_75t_L g2299 ( 
.A(n_2263),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2056),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2059),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2082),
.Y(n_2302)
);

OA21x2_ASAP7_75t_L g2303 ( 
.A1(n_2254),
.A2(n_2283),
.B(n_2279),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2258),
.B(n_2187),
.Y(n_2304)
);

INVx3_ASAP7_75t_L g2305 ( 
.A(n_2028),
.Y(n_2305)
);

BUFx6f_ASAP7_75t_L g2306 ( 
.A(n_2267),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2106),
.Y(n_2307)
);

BUFx8_ASAP7_75t_L g2308 ( 
.A(n_2043),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2107),
.Y(n_2309)
);

CKINVDCx20_ASAP7_75t_R g2310 ( 
.A(n_2040),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2084),
.Y(n_2311)
);

AOI222xp33_ASAP7_75t_L g2312 ( 
.A1(n_2055),
.A2(n_2243),
.B1(n_2209),
.B2(n_2216),
.C1(n_2094),
.C2(n_2065),
.Y(n_2312)
);

INVx1_ASAP7_75t_SL g2313 ( 
.A(n_2033),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2084),
.Y(n_2314)
);

OA21x2_ASAP7_75t_L g2315 ( 
.A1(n_2272),
.A2(n_2279),
.B(n_2270),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2138),
.Y(n_2316)
);

AOI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_2045),
.A2(n_2262),
.B1(n_2271),
.B2(n_2216),
.Y(n_2317)
);

OAI21x1_ASAP7_75t_L g2318 ( 
.A1(n_2264),
.A2(n_2275),
.B(n_2265),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2269),
.B(n_2105),
.Y(n_2319)
);

AOI22xp5_ASAP7_75t_L g2320 ( 
.A1(n_2271),
.A2(n_2261),
.B1(n_2033),
.B2(n_2055),
.Y(n_2320)
);

AOI21x1_ASAP7_75t_L g2321 ( 
.A1(n_2124),
.A2(n_2089),
.B(n_2284),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2191),
.B(n_2193),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2096),
.Y(n_2323)
);

INVx5_ASAP7_75t_L g2324 ( 
.A(n_2257),
.Y(n_2324)
);

OR2x6_ASAP7_75t_L g2325 ( 
.A(n_2093),
.B(n_2155),
.Y(n_2325)
);

BUFx4f_ASAP7_75t_SL g2326 ( 
.A(n_2040),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2282),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2288),
.Y(n_2328)
);

OAI22xp33_ASAP7_75t_R g2329 ( 
.A1(n_2278),
.A2(n_2172),
.B1(n_2065),
.B2(n_2114),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2052),
.B(n_2261),
.Y(n_2330)
);

AND2x4_ASAP7_75t_L g2331 ( 
.A(n_2150),
.B(n_2266),
.Y(n_2331)
);

BUFx8_ASAP7_75t_L g2332 ( 
.A(n_2060),
.Y(n_2332)
);

INVx3_ASAP7_75t_L g2333 ( 
.A(n_2028),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_2159),
.B(n_2104),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2166),
.Y(n_2335)
);

BUFx12f_ASAP7_75t_L g2336 ( 
.A(n_2285),
.Y(n_2336)
);

OAI21x1_ASAP7_75t_L g2337 ( 
.A1(n_2272),
.A2(n_2064),
.B(n_2031),
.Y(n_2337)
);

INVx1_ASAP7_75t_SL g2338 ( 
.A(n_2115),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2128),
.Y(n_2339)
);

BUFx2_ASAP7_75t_L g2340 ( 
.A(n_2267),
.Y(n_2340)
);

INVx1_ASAP7_75t_SL g2341 ( 
.A(n_2115),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2128),
.Y(n_2342)
);

BUFx3_ASAP7_75t_L g2343 ( 
.A(n_2257),
.Y(n_2343)
);

BUFx3_ASAP7_75t_L g2344 ( 
.A(n_2257),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2046),
.Y(n_2345)
);

AOI22xp33_ASAP7_75t_L g2346 ( 
.A1(n_2224),
.A2(n_2175),
.B1(n_2244),
.B2(n_2221),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2068),
.Y(n_2347)
);

INVx6_ASAP7_75t_L g2348 ( 
.A(n_2148),
.Y(n_2348)
);

INVx1_ASAP7_75t_SL g2349 ( 
.A(n_2158),
.Y(n_2349)
);

INVx3_ASAP7_75t_L g2350 ( 
.A(n_2032),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2122),
.B(n_2110),
.Y(n_2351)
);

BUFx3_ASAP7_75t_L g2352 ( 
.A(n_2148),
.Y(n_2352)
);

AOI22xp33_ASAP7_75t_L g2353 ( 
.A1(n_2094),
.A2(n_2239),
.B1(n_2246),
.B2(n_2036),
.Y(n_2353)
);

OA21x2_ASAP7_75t_L g2354 ( 
.A1(n_2273),
.A2(n_2126),
.B(n_2149),
.Y(n_2354)
);

AOI22xp33_ASAP7_75t_L g2355 ( 
.A1(n_2036),
.A2(n_2217),
.B1(n_2251),
.B2(n_2200),
.Y(n_2355)
);

BUFx2_ASAP7_75t_L g2356 ( 
.A(n_2268),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2165),
.Y(n_2357)
);

INVx6_ASAP7_75t_L g2358 ( 
.A(n_2032),
.Y(n_2358)
);

OAI22xp5_ASAP7_75t_L g2359 ( 
.A1(n_2049),
.A2(n_2219),
.B1(n_2108),
.B2(n_2286),
.Y(n_2359)
);

CKINVDCx11_ASAP7_75t_R g2360 ( 
.A(n_2034),
.Y(n_2360)
);

HB1xp67_ASAP7_75t_L g2361 ( 
.A(n_2100),
.Y(n_2361)
);

BUFx6f_ASAP7_75t_L g2362 ( 
.A(n_2268),
.Y(n_2362)
);

BUFx3_ASAP7_75t_L g2363 ( 
.A(n_2038),
.Y(n_2363)
);

INVx3_ASAP7_75t_L g2364 ( 
.A(n_2289),
.Y(n_2364)
);

AOI21x1_ASAP7_75t_L g2365 ( 
.A1(n_2124),
.A2(n_2089),
.B(n_2079),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2276),
.B(n_2130),
.Y(n_2366)
);

OAI22xp33_ASAP7_75t_SL g2367 ( 
.A1(n_2150),
.A2(n_2108),
.B1(n_2194),
.B2(n_2079),
.Y(n_2367)
);

HB1xp67_ASAP7_75t_L g2368 ( 
.A(n_2100),
.Y(n_2368)
);

CKINVDCx20_ASAP7_75t_R g2369 ( 
.A(n_2038),
.Y(n_2369)
);

AOI21x1_ASAP7_75t_L g2370 ( 
.A1(n_2136),
.A2(n_2150),
.B(n_2206),
.Y(n_2370)
);

BUFx12f_ASAP7_75t_L g2371 ( 
.A(n_2050),
.Y(n_2371)
);

AOI22xp33_ASAP7_75t_SL g2372 ( 
.A1(n_2154),
.A2(n_2123),
.B1(n_2219),
.B2(n_2119),
.Y(n_2372)
);

INVx5_ASAP7_75t_L g2373 ( 
.A(n_2289),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2111),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2266),
.B(n_2280),
.Y(n_2375)
);

NOR2xp33_ASAP7_75t_L g2376 ( 
.A(n_2112),
.B(n_2253),
.Y(n_2376)
);

AOI22xp33_ASAP7_75t_L g2377 ( 
.A1(n_2251),
.A2(n_2200),
.B1(n_2238),
.B2(n_2286),
.Y(n_2377)
);

INVx6_ASAP7_75t_L g2378 ( 
.A(n_2037),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2204),
.B(n_2202),
.Y(n_2379)
);

INVx4_ASAP7_75t_L g2380 ( 
.A(n_2050),
.Y(n_2380)
);

CKINVDCx5p33_ASAP7_75t_R g2381 ( 
.A(n_2039),
.Y(n_2381)
);

AOI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_2067),
.A2(n_2121),
.B1(n_2287),
.B2(n_2201),
.Y(n_2382)
);

OAI21x1_ASAP7_75t_L g2383 ( 
.A1(n_2098),
.A2(n_2072),
.B(n_2070),
.Y(n_2383)
);

AO21x1_ASAP7_75t_SL g2384 ( 
.A1(n_2062),
.A2(n_2103),
.B(n_2219),
.Y(n_2384)
);

AO21x2_ASAP7_75t_L g2385 ( 
.A1(n_2041),
.A2(n_2058),
.B(n_2044),
.Y(n_2385)
);

NAND2x1p5_ASAP7_75t_L g2386 ( 
.A(n_2219),
.B(n_2057),
.Y(n_2386)
);

HB1xp67_ASAP7_75t_L g2387 ( 
.A(n_2062),
.Y(n_2387)
);

BUFx2_ASAP7_75t_SL g2388 ( 
.A(n_2037),
.Y(n_2388)
);

INVx2_ASAP7_75t_SL g2389 ( 
.A(n_2029),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2205),
.Y(n_2390)
);

BUFx2_ASAP7_75t_L g2391 ( 
.A(n_2103),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2205),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2066),
.Y(n_2393)
);

OR2x2_ASAP7_75t_L g2394 ( 
.A(n_2114),
.B(n_2048),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2198),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_2078),
.B(n_2113),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2198),
.Y(n_2397)
);

INVx5_ASAP7_75t_L g2398 ( 
.A(n_2097),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2108),
.Y(n_2399)
);

AOI22xp33_ASAP7_75t_L g2400 ( 
.A1(n_2238),
.A2(n_2250),
.B1(n_2252),
.B2(n_2241),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2140),
.Y(n_2401)
);

BUFx3_ASAP7_75t_L g2402 ( 
.A(n_2277),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2127),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2185),
.Y(n_2404)
);

BUFx3_ASAP7_75t_L g2405 ( 
.A(n_2069),
.Y(n_2405)
);

INVx4_ASAP7_75t_L g2406 ( 
.A(n_2255),
.Y(n_2406)
);

INVx1_ASAP7_75t_SL g2407 ( 
.A(n_2078),
.Y(n_2407)
);

BUFx8_ASAP7_75t_L g2408 ( 
.A(n_2218),
.Y(n_2408)
);

AOI21x1_ASAP7_75t_L g2409 ( 
.A1(n_2235),
.A2(n_2126),
.B(n_2109),
.Y(n_2409)
);

OAI22xp5_ASAP7_75t_L g2410 ( 
.A1(n_2113),
.A2(n_2102),
.B1(n_2142),
.B2(n_2196),
.Y(n_2410)
);

BUFx12f_ASAP7_75t_L g2411 ( 
.A(n_2163),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_2039),
.Y(n_2412)
);

OAI22xp33_ASAP7_75t_L g2413 ( 
.A1(n_2086),
.A2(n_2234),
.B1(n_2092),
.B2(n_2242),
.Y(n_2413)
);

INVx2_ASAP7_75t_SL g2414 ( 
.A(n_2029),
.Y(n_2414)
);

OAI22xp5_ASAP7_75t_L g2415 ( 
.A1(n_2196),
.A2(n_2253),
.B1(n_2236),
.B2(n_2109),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2095),
.B(n_2101),
.Y(n_2416)
);

BUFx3_ASAP7_75t_L g2417 ( 
.A(n_2095),
.Y(n_2417)
);

BUFx8_ASAP7_75t_L g2418 ( 
.A(n_2218),
.Y(n_2418)
);

OAI21x1_ASAP7_75t_L g2419 ( 
.A1(n_2132),
.A2(n_2134),
.B(n_2135),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2101),
.B(n_2088),
.Y(n_2420)
);

BUFx3_ASAP7_75t_L g2421 ( 
.A(n_2097),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2255),
.Y(n_2422)
);

BUFx3_ASAP7_75t_L g2423 ( 
.A(n_2097),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2259),
.Y(n_2424)
);

AOI21x1_ASAP7_75t_L g2425 ( 
.A1(n_2207),
.A2(n_2211),
.B(n_2195),
.Y(n_2425)
);

NAND2x1p5_ASAP7_75t_L g2426 ( 
.A(n_2051),
.B(n_2053),
.Y(n_2426)
);

BUFx3_ASAP7_75t_L g2427 ( 
.A(n_2099),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2259),
.Y(n_2428)
);

AND2x2_ASAP7_75t_SL g2429 ( 
.A(n_2133),
.B(n_2085),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2260),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2260),
.Y(n_2431)
);

HB1xp67_ASAP7_75t_L g2432 ( 
.A(n_2117),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2274),
.Y(n_2433)
);

AO21x2_ASAP7_75t_L g2434 ( 
.A1(n_2041),
.A2(n_2058),
.B(n_2044),
.Y(n_2434)
);

OAI22xp33_ASAP7_75t_L g2435 ( 
.A1(n_2234),
.A2(n_2242),
.B1(n_2178),
.B2(n_2197),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2080),
.B(n_2237),
.Y(n_2436)
);

HB1xp67_ASAP7_75t_L g2437 ( 
.A(n_2117),
.Y(n_2437)
);

CKINVDCx20_ASAP7_75t_R g2438 ( 
.A(n_2099),
.Y(n_2438)
);

OR2x2_ASAP7_75t_L g2439 ( 
.A(n_2125),
.B(n_2147),
.Y(n_2439)
);

AOI22xp33_ASAP7_75t_L g2440 ( 
.A1(n_2203),
.A2(n_2231),
.B1(n_2248),
.B2(n_2245),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2274),
.Y(n_2441)
);

OAI22xp33_ASAP7_75t_L g2442 ( 
.A1(n_2164),
.A2(n_2197),
.B1(n_2192),
.B2(n_2133),
.Y(n_2442)
);

AOI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2075),
.A2(n_2225),
.B(n_2042),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2232),
.Y(n_2444)
);

AOI22xp33_ASAP7_75t_L g2445 ( 
.A1(n_2248),
.A2(n_2245),
.B1(n_2225),
.B2(n_2223),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2171),
.Y(n_2446)
);

BUFx2_ASAP7_75t_SL g2447 ( 
.A(n_2164),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2080),
.B(n_2237),
.Y(n_2448)
);

HB1xp67_ASAP7_75t_L g2449 ( 
.A(n_2152),
.Y(n_2449)
);

BUFx6f_ASAP7_75t_SL g2450 ( 
.A(n_2222),
.Y(n_2450)
);

AND2x2_ASAP7_75t_L g2451 ( 
.A(n_2230),
.B(n_2030),
.Y(n_2451)
);

BUFx2_ASAP7_75t_L g2452 ( 
.A(n_2153),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2213),
.Y(n_2453)
);

INVx2_ASAP7_75t_SL g2454 ( 
.A(n_2139),
.Y(n_2454)
);

BUFx10_ASAP7_75t_L g2455 ( 
.A(n_2076),
.Y(n_2455)
);

AOI21x1_ASAP7_75t_L g2456 ( 
.A1(n_2195),
.A2(n_2240),
.B(n_2228),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2229),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2446),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2366),
.B(n_2160),
.Y(n_2459)
);

NOR2xp33_ASAP7_75t_R g2460 ( 
.A(n_2326),
.B(n_2310),
.Y(n_2460)
);

BUFx2_ASAP7_75t_L g2461 ( 
.A(n_2405),
.Y(n_2461)
);

HB1xp67_ASAP7_75t_L g2462 ( 
.A(n_2387),
.Y(n_2462)
);

INVx3_ASAP7_75t_L g2463 ( 
.A(n_2324),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2300),
.Y(n_2464)
);

NOR2xp67_ASAP7_75t_L g2465 ( 
.A(n_2324),
.B(n_2222),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2351),
.B(n_2087),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_SL g2467 ( 
.A(n_2367),
.B(n_2123),
.Y(n_2467)
);

INVx6_ASAP7_75t_L g2468 ( 
.A(n_2324),
.Y(n_2468)
);

OAI21xp33_ASAP7_75t_L g2469 ( 
.A1(n_2295),
.A2(n_2294),
.B(n_2317),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_2360),
.Y(n_2470)
);

BUFx2_ASAP7_75t_L g2471 ( 
.A(n_2406),
.Y(n_2471)
);

AND2x2_ASAP7_75t_L g2472 ( 
.A(n_2330),
.B(n_2087),
.Y(n_2472)
);

NOR2xp33_ASAP7_75t_R g2473 ( 
.A(n_2369),
.B(n_2076),
.Y(n_2473)
);

CKINVDCx5p33_ASAP7_75t_R g2474 ( 
.A(n_2308),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2301),
.Y(n_2475)
);

CKINVDCx16_ASAP7_75t_R g2476 ( 
.A(n_2343),
.Y(n_2476)
);

HB1xp67_ASAP7_75t_L g2477 ( 
.A(n_2387),
.Y(n_2477)
);

CKINVDCx16_ASAP7_75t_R g2478 ( 
.A(n_2344),
.Y(n_2478)
);

NAND2xp33_ASAP7_75t_R g2479 ( 
.A(n_2452),
.B(n_2210),
.Y(n_2479)
);

NOR3xp33_ASAP7_75t_SL g2480 ( 
.A(n_2413),
.B(n_2226),
.C(n_2146),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2319),
.B(n_2131),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2302),
.Y(n_2482)
);

BUFx2_ASAP7_75t_L g2483 ( 
.A(n_2406),
.Y(n_2483)
);

AOI22xp33_ASAP7_75t_L g2484 ( 
.A1(n_2294),
.A2(n_2210),
.B1(n_2123),
.B2(n_2167),
.Y(n_2484)
);

CKINVDCx12_ASAP7_75t_R g2485 ( 
.A(n_2325),
.Y(n_2485)
);

NOR2xp33_ASAP7_75t_R g2486 ( 
.A(n_2290),
.B(n_2146),
.Y(n_2486)
);

AO31x2_ASAP7_75t_L g2487 ( 
.A1(n_2443),
.A2(n_2184),
.A3(n_2220),
.B(n_2188),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_2308),
.Y(n_2488)
);

AO31x2_ASAP7_75t_L g2489 ( 
.A1(n_2443),
.A2(n_2184),
.A3(n_2188),
.B(n_2075),
.Y(n_2489)
);

HB1xp67_ASAP7_75t_L g2490 ( 
.A(n_2313),
.Y(n_2490)
);

OAI22xp5_ASAP7_75t_L g2491 ( 
.A1(n_2415),
.A2(n_2236),
.B1(n_2215),
.B2(n_2214),
.Y(n_2491)
);

OR2x6_ASAP7_75t_L g2492 ( 
.A(n_2388),
.B(n_2141),
.Y(n_2492)
);

INVx11_ASAP7_75t_L g2493 ( 
.A(n_2408),
.Y(n_2493)
);

INVxp33_ASAP7_75t_SL g2494 ( 
.A(n_2352),
.Y(n_2494)
);

CKINVDCx5p33_ASAP7_75t_R g2495 ( 
.A(n_2336),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2334),
.B(n_2190),
.Y(n_2496)
);

O2A1O1Ixp33_ASAP7_75t_SL g2497 ( 
.A1(n_2413),
.A2(n_2073),
.B(n_2063),
.C(n_2173),
.Y(n_2497)
);

AOI22xp33_ASAP7_75t_SL g2498 ( 
.A1(n_2415),
.A2(n_2123),
.B1(n_2153),
.B2(n_2192),
.Y(n_2498)
);

NOR2x1_ASAP7_75t_SL g2499 ( 
.A(n_2384),
.B(n_2325),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2307),
.Y(n_2500)
);

CKINVDCx20_ASAP7_75t_R g2501 ( 
.A(n_2332),
.Y(n_2501)
);

XOR2xp5_ASAP7_75t_L g2502 ( 
.A(n_2381),
.B(n_2227),
.Y(n_2502)
);

NAND2xp33_ASAP7_75t_R g2503 ( 
.A(n_2305),
.B(n_2226),
.Y(n_2503)
);

OR2x6_ASAP7_75t_L g2504 ( 
.A(n_2348),
.B(n_2192),
.Y(n_2504)
);

OR2x2_ASAP7_75t_L g2505 ( 
.A(n_2394),
.B(n_2338),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2393),
.B(n_2167),
.Y(n_2506)
);

NAND3xp33_ASAP7_75t_SL g2507 ( 
.A(n_2312),
.B(n_2215),
.C(n_2214),
.Y(n_2507)
);

BUFx12f_ASAP7_75t_L g2508 ( 
.A(n_2332),
.Y(n_2508)
);

INVx4_ASAP7_75t_L g2509 ( 
.A(n_2348),
.Y(n_2509)
);

NOR2xp33_ASAP7_75t_L g2510 ( 
.A(n_2427),
.B(n_2180),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2309),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2416),
.B(n_2190),
.Y(n_2512)
);

NOR2xp33_ASAP7_75t_R g2513 ( 
.A(n_2363),
.B(n_2163),
.Y(n_2513)
);

NAND3xp33_ASAP7_75t_SL g2514 ( 
.A(n_2312),
.B(n_2145),
.C(n_2083),
.Y(n_2514)
);

NAND2xp33_ASAP7_75t_SL g2515 ( 
.A(n_2410),
.B(n_2180),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2346),
.B(n_2233),
.Y(n_2516)
);

CKINVDCx8_ASAP7_75t_R g2517 ( 
.A(n_2398),
.Y(n_2517)
);

OAI22xp5_ASAP7_75t_L g2518 ( 
.A1(n_2382),
.A2(n_2145),
.B1(n_2083),
.B2(n_2162),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2316),
.Y(n_2519)
);

BUFx4f_ASAP7_75t_L g2520 ( 
.A(n_2411),
.Y(n_2520)
);

AOI22xp33_ASAP7_75t_SL g2521 ( 
.A1(n_2359),
.A2(n_2123),
.B1(n_2061),
.B2(n_2208),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2444),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2291),
.B(n_2233),
.Y(n_2523)
);

BUFx3_ASAP7_75t_L g2524 ( 
.A(n_2408),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2453),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2457),
.Y(n_2526)
);

NAND2xp33_ASAP7_75t_R g2527 ( 
.A(n_2305),
.B(n_2189),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2323),
.Y(n_2528)
);

INVx2_ASAP7_75t_SL g2529 ( 
.A(n_2418),
.Y(n_2529)
);

CKINVDCx16_ASAP7_75t_R g2530 ( 
.A(n_2402),
.Y(n_2530)
);

CKINVDCx5p33_ASAP7_75t_R g2531 ( 
.A(n_2412),
.Y(n_2531)
);

AOI22xp33_ASAP7_75t_L g2532 ( 
.A1(n_2377),
.A2(n_2123),
.B1(n_2177),
.B2(n_2249),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2296),
.B(n_2116),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2420),
.B(n_2177),
.Y(n_2534)
);

AND2x4_ASAP7_75t_L g2535 ( 
.A(n_2292),
.B(n_2071),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2390),
.Y(n_2536)
);

OR2x6_ASAP7_75t_L g2537 ( 
.A(n_2325),
.B(n_2143),
.Y(n_2537)
);

AND2x4_ASAP7_75t_SL g2538 ( 
.A(n_2333),
.B(n_2169),
.Y(n_2538)
);

NOR2xp33_ASAP7_75t_R g2539 ( 
.A(n_2438),
.B(n_2071),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2392),
.Y(n_2540)
);

CKINVDCx5p33_ASAP7_75t_R g2541 ( 
.A(n_2418),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2375),
.B(n_2247),
.Y(n_2542)
);

HB1xp67_ASAP7_75t_L g2543 ( 
.A(n_2313),
.Y(n_2543)
);

BUFx3_ASAP7_75t_L g2544 ( 
.A(n_2417),
.Y(n_2544)
);

AOI22xp33_ASAP7_75t_L g2545 ( 
.A1(n_2382),
.A2(n_2161),
.B1(n_2199),
.B2(n_2176),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2297),
.B(n_2116),
.Y(n_2546)
);

NAND3xp33_ASAP7_75t_SL g2547 ( 
.A(n_2349),
.B(n_2227),
.C(n_2168),
.Y(n_2547)
);

NAND2xp33_ASAP7_75t_R g2548 ( 
.A(n_2333),
.B(n_2174),
.Y(n_2548)
);

NAND2xp33_ASAP7_75t_R g2549 ( 
.A(n_2350),
.B(n_2174),
.Y(n_2549)
);

INVx2_ASAP7_75t_SL g2550 ( 
.A(n_2358),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2335),
.B(n_2090),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2338),
.B(n_2199),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2327),
.B(n_2090),
.Y(n_2553)
);

AND2x2_ASAP7_75t_L g2554 ( 
.A(n_2341),
.B(n_2176),
.Y(n_2554)
);

INVxp67_ASAP7_75t_SL g2555 ( 
.A(n_2432),
.Y(n_2555)
);

NOR2x1_ASAP7_75t_L g2556 ( 
.A(n_2435),
.B(n_2212),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2328),
.B(n_2156),
.Y(n_2557)
);

INVx1_ASAP7_75t_SL g2558 ( 
.A(n_2358),
.Y(n_2558)
);

NAND2xp33_ASAP7_75t_R g2559 ( 
.A(n_2350),
.B(n_2157),
.Y(n_2559)
);

HB1xp67_ASAP7_75t_L g2560 ( 
.A(n_2407),
.Y(n_2560)
);

AND2x2_ASAP7_75t_SL g2561 ( 
.A(n_2429),
.B(n_2281),
.Y(n_2561)
);

INVx4_ASAP7_75t_SL g2562 ( 
.A(n_2378),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_2401),
.B(n_2156),
.Y(n_2563)
);

CKINVDCx16_ASAP7_75t_R g2564 ( 
.A(n_2371),
.Y(n_2564)
);

OR2x2_ASAP7_75t_L g2565 ( 
.A(n_2341),
.B(n_2047),
.Y(n_2565)
);

AOI22xp33_ASAP7_75t_L g2566 ( 
.A1(n_2403),
.A2(n_2212),
.B1(n_2091),
.B2(n_2118),
.Y(n_2566)
);

OR2x6_ASAP7_75t_L g2567 ( 
.A(n_2447),
.B(n_2170),
.Y(n_2567)
);

AND2x2_ASAP7_75t_L g2568 ( 
.A(n_2407),
.B(n_2181),
.Y(n_2568)
);

BUFx3_ASAP7_75t_L g2569 ( 
.A(n_2378),
.Y(n_2569)
);

OR2x6_ASAP7_75t_L g2570 ( 
.A(n_2380),
.B(n_2170),
.Y(n_2570)
);

AND2x4_ASAP7_75t_L g2571 ( 
.A(n_2331),
.B(n_2129),
.Y(n_2571)
);

NOR3xp33_ASAP7_75t_SL g2572 ( 
.A(n_2435),
.B(n_2442),
.C(n_2376),
.Y(n_2572)
);

OR2x6_ASAP7_75t_L g2573 ( 
.A(n_2380),
.B(n_2168),
.Y(n_2573)
);

CKINVDCx5p33_ASAP7_75t_R g2574 ( 
.A(n_2455),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2396),
.B(n_2181),
.Y(n_2575)
);

NOR2xp33_ASAP7_75t_R g2576 ( 
.A(n_2364),
.B(n_2144),
.Y(n_2576)
);

AND2x2_ASAP7_75t_SL g2577 ( 
.A(n_2353),
.B(n_2281),
.Y(n_2577)
);

BUFx12f_ASAP7_75t_L g2578 ( 
.A(n_2455),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2345),
.Y(n_2579)
);

HB1xp67_ASAP7_75t_L g2580 ( 
.A(n_2432),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2347),
.Y(n_2581)
);

NOR2xp33_ASAP7_75t_R g2582 ( 
.A(n_2373),
.B(n_2137),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2322),
.B(n_2047),
.Y(n_2583)
);

OR2x6_ASAP7_75t_L g2584 ( 
.A(n_2421),
.B(n_2186),
.Y(n_2584)
);

INVx4_ASAP7_75t_L g2585 ( 
.A(n_2373),
.Y(n_2585)
);

INVx4_ASAP7_75t_L g2586 ( 
.A(n_2398),
.Y(n_2586)
);

BUFx3_ASAP7_75t_L g2587 ( 
.A(n_2423),
.Y(n_2587)
);

INVx3_ASAP7_75t_L g2588 ( 
.A(n_2373),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2357),
.Y(n_2589)
);

BUFx3_ASAP7_75t_L g2590 ( 
.A(n_2398),
.Y(n_2590)
);

OR2x6_ASAP7_75t_L g2591 ( 
.A(n_2340),
.B(n_2356),
.Y(n_2591)
);

NOR2xp33_ASAP7_75t_L g2592 ( 
.A(n_2454),
.B(n_2151),
.Y(n_2592)
);

INVxp67_ASAP7_75t_L g2593 ( 
.A(n_2439),
.Y(n_2593)
);

INVxp67_ASAP7_75t_L g2594 ( 
.A(n_2461),
.Y(n_2594)
);

AOI22xp33_ASAP7_75t_SL g2595 ( 
.A1(n_2499),
.A2(n_2367),
.B1(n_2410),
.B2(n_2359),
.Y(n_2595)
);

AND2x4_ASAP7_75t_L g2596 ( 
.A(n_2554),
.B(n_2370),
.Y(n_2596)
);

HB1xp67_ASAP7_75t_L g2597 ( 
.A(n_2580),
.Y(n_2597)
);

OR2x2_ASAP7_75t_L g2598 ( 
.A(n_2555),
.B(n_2490),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2542),
.B(n_2299),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2552),
.B(n_2299),
.Y(n_2600)
);

INVxp67_ASAP7_75t_SL g2601 ( 
.A(n_2462),
.Y(n_2601)
);

HB1xp67_ASAP7_75t_L g2602 ( 
.A(n_2477),
.Y(n_2602)
);

OR2x2_ASAP7_75t_SL g2603 ( 
.A(n_2547),
.B(n_2303),
.Y(n_2603)
);

INVx2_ASAP7_75t_SL g2604 ( 
.A(n_2576),
.Y(n_2604)
);

AND2x4_ASAP7_75t_L g2605 ( 
.A(n_2487),
.B(n_2365),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2458),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2522),
.Y(n_2607)
);

HB1xp67_ASAP7_75t_L g2608 ( 
.A(n_2543),
.Y(n_2608)
);

AND2x2_ASAP7_75t_L g2609 ( 
.A(n_2557),
.B(n_2436),
.Y(n_2609)
);

HB1xp67_ASAP7_75t_L g2610 ( 
.A(n_2560),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2525),
.Y(n_2611)
);

AND2x2_ASAP7_75t_L g2612 ( 
.A(n_2563),
.B(n_2436),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2526),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2583),
.B(n_2448),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2533),
.B(n_2448),
.Y(n_2615)
);

NOR2xp67_ASAP7_75t_L g2616 ( 
.A(n_2585),
.B(n_2389),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2546),
.B(n_2303),
.Y(n_2617)
);

OAI21xp5_ASAP7_75t_L g2618 ( 
.A1(n_2491),
.A2(n_2445),
.B(n_2355),
.Y(n_2618)
);

AND2x2_ASAP7_75t_L g2619 ( 
.A(n_2551),
.B(n_2298),
.Y(n_2619)
);

HB1xp67_ASAP7_75t_L g2620 ( 
.A(n_2472),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2464),
.Y(n_2621)
);

NAND3xp33_ASAP7_75t_L g2622 ( 
.A(n_2479),
.B(n_2440),
.C(n_2320),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2475),
.Y(n_2623)
);

AND2x2_ASAP7_75t_L g2624 ( 
.A(n_2553),
.B(n_2315),
.Y(n_2624)
);

BUFx2_ASAP7_75t_L g2625 ( 
.A(n_2471),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2523),
.B(n_2315),
.Y(n_2626)
);

HB1xp67_ASAP7_75t_L g2627 ( 
.A(n_2466),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2565),
.B(n_2482),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2500),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2511),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2519),
.B(n_2385),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2536),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2540),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2545),
.B(n_2434),
.Y(n_2634)
);

AND2x2_ASAP7_75t_L g2635 ( 
.A(n_2516),
.B(n_2434),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2505),
.B(n_2437),
.Y(n_2636)
);

NOR2xp33_ASAP7_75t_L g2637 ( 
.A(n_2494),
.B(n_2451),
.Y(n_2637)
);

AOI221xp5_ASAP7_75t_L g2638 ( 
.A1(n_2469),
.A2(n_2311),
.B1(n_2314),
.B2(n_2339),
.C(n_2342),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2528),
.Y(n_2639)
);

INVxp67_ASAP7_75t_SL g2640 ( 
.A(n_2527),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2579),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2581),
.Y(n_2642)
);

BUFx2_ASAP7_75t_L g2643 ( 
.A(n_2483),
.Y(n_2643)
);

BUFx2_ASAP7_75t_L g2644 ( 
.A(n_2591),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2589),
.Y(n_2645)
);

NOR2x1_ASAP7_75t_SL g2646 ( 
.A(n_2537),
.B(n_2422),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2506),
.B(n_2449),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2484),
.B(n_2449),
.Y(n_2648)
);

INVx3_ASAP7_75t_L g2649 ( 
.A(n_2585),
.Y(n_2649)
);

AND2x2_ASAP7_75t_L g2650 ( 
.A(n_2496),
.B(n_2379),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2489),
.Y(n_2651)
);

OR2x2_ASAP7_75t_L g2652 ( 
.A(n_2593),
.B(n_2379),
.Y(n_2652)
);

INVxp67_ASAP7_75t_L g2653 ( 
.A(n_2544),
.Y(n_2653)
);

HB1xp67_ASAP7_75t_L g2654 ( 
.A(n_2591),
.Y(n_2654)
);

INVx5_ASAP7_75t_L g2655 ( 
.A(n_2537),
.Y(n_2655)
);

AND2x2_ASAP7_75t_L g2656 ( 
.A(n_2489),
.B(n_2304),
.Y(n_2656)
);

HB1xp67_ASAP7_75t_L g2657 ( 
.A(n_2481),
.Y(n_2657)
);

AND2x2_ASAP7_75t_L g2658 ( 
.A(n_2489),
.B(n_2304),
.Y(n_2658)
);

INVx2_ASAP7_75t_SL g2659 ( 
.A(n_2468),
.Y(n_2659)
);

NOR2xp33_ASAP7_75t_L g2660 ( 
.A(n_2476),
.B(n_2414),
.Y(n_2660)
);

NAND3xp33_ASAP7_75t_L g2661 ( 
.A(n_2572),
.B(n_2400),
.C(n_2404),
.Y(n_2661)
);

BUFx3_ASAP7_75t_L g2662 ( 
.A(n_2468),
.Y(n_2662)
);

BUFx3_ASAP7_75t_L g2663 ( 
.A(n_2517),
.Y(n_2663)
);

INVxp67_ASAP7_75t_L g2664 ( 
.A(n_2459),
.Y(n_2664)
);

INVx2_ASAP7_75t_SL g2665 ( 
.A(n_2561),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2556),
.Y(n_2666)
);

CKINVDCx5p33_ASAP7_75t_R g2667 ( 
.A(n_2460),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2512),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2568),
.Y(n_2669)
);

AOI22xp33_ASAP7_75t_L g2670 ( 
.A1(n_2498),
.A2(n_2329),
.B1(n_2399),
.B2(n_2374),
.Y(n_2670)
);

INVxp67_ASAP7_75t_L g2671 ( 
.A(n_2492),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2534),
.Y(n_2672)
);

BUFx3_ASAP7_75t_L g2673 ( 
.A(n_2590),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2624),
.Y(n_2674)
);

AND2x4_ASAP7_75t_L g2675 ( 
.A(n_2596),
.B(n_2419),
.Y(n_2675)
);

CKINVDCx20_ASAP7_75t_R g2676 ( 
.A(n_2667),
.Y(n_2676)
);

BUFx2_ASAP7_75t_L g2677 ( 
.A(n_2625),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2614),
.B(n_2566),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2614),
.B(n_2521),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2631),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2615),
.B(n_2361),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2599),
.B(n_2456),
.Y(n_2682)
);

AND2x2_ASAP7_75t_L g2683 ( 
.A(n_2599),
.B(n_2409),
.Y(n_2683)
);

AOI21xp5_ASAP7_75t_SL g2684 ( 
.A1(n_2604),
.A2(n_2514),
.B(n_2507),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2615),
.B(n_2361),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2609),
.B(n_2321),
.Y(n_2686)
);

AND2x4_ASAP7_75t_L g2687 ( 
.A(n_2596),
.B(n_2383),
.Y(n_2687)
);

INVxp67_ASAP7_75t_SL g2688 ( 
.A(n_2625),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2609),
.B(n_2354),
.Y(n_2689)
);

AOI22xp33_ASAP7_75t_L g2690 ( 
.A1(n_2661),
.A2(n_2515),
.B1(n_2532),
.B2(n_2577),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2617),
.Y(n_2691)
);

INVxp67_ASAP7_75t_SL g2692 ( 
.A(n_2597),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2628),
.B(n_2368),
.Y(n_2693)
);

AND2x2_ASAP7_75t_L g2694 ( 
.A(n_2612),
.B(n_2425),
.Y(n_2694)
);

HB1xp67_ASAP7_75t_L g2695 ( 
.A(n_2643),
.Y(n_2695)
);

AND2x4_ASAP7_75t_L g2696 ( 
.A(n_2596),
.B(n_2337),
.Y(n_2696)
);

NOR2xp33_ASAP7_75t_R g2697 ( 
.A(n_2667),
.B(n_2501),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2635),
.B(n_2467),
.Y(n_2698)
);

BUFx3_ASAP7_75t_L g2699 ( 
.A(n_2673),
.Y(n_2699)
);

AND2x2_ASAP7_75t_L g2700 ( 
.A(n_2635),
.B(n_2600),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2626),
.Y(n_2701)
);

AND2x2_ASAP7_75t_L g2702 ( 
.A(n_2600),
.B(n_2650),
.Y(n_2702)
);

INVxp33_ASAP7_75t_L g2703 ( 
.A(n_2660),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2626),
.B(n_2656),
.Y(n_2704)
);

NAND4xp25_ASAP7_75t_L g2705 ( 
.A(n_2670),
.B(n_2503),
.C(n_2524),
.D(n_2465),
.Y(n_2705)
);

AND2x2_ASAP7_75t_L g2706 ( 
.A(n_2658),
.B(n_2318),
.Y(n_2706)
);

INVx3_ASAP7_75t_L g2707 ( 
.A(n_2605),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2651),
.Y(n_2708)
);

AND2x2_ASAP7_75t_L g2709 ( 
.A(n_2704),
.B(n_2619),
.Y(n_2709)
);

OR2x2_ASAP7_75t_L g2710 ( 
.A(n_2674),
.B(n_2608),
.Y(n_2710)
);

AND2x4_ASAP7_75t_L g2711 ( 
.A(n_2707),
.B(n_2605),
.Y(n_2711)
);

OR2x2_ASAP7_75t_L g2712 ( 
.A(n_2674),
.B(n_2610),
.Y(n_2712)
);

INVx1_ASAP7_75t_SL g2713 ( 
.A(n_2677),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2680),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2704),
.B(n_2634),
.Y(n_2715)
);

INVx2_ASAP7_75t_SL g2716 ( 
.A(n_2699),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2674),
.B(n_2634),
.Y(n_2717)
);

INVx5_ASAP7_75t_L g2718 ( 
.A(n_2699),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2702),
.B(n_2602),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2702),
.B(n_2601),
.Y(n_2720)
);

INVx1_ASAP7_75t_SL g2721 ( 
.A(n_2697),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2708),
.Y(n_2722)
);

HB1xp67_ASAP7_75t_L g2723 ( 
.A(n_2677),
.Y(n_2723)
);

INVx1_ASAP7_75t_SL g2724 ( 
.A(n_2699),
.Y(n_2724)
);

HB1xp67_ASAP7_75t_L g2725 ( 
.A(n_2695),
.Y(n_2725)
);

OR2x2_ASAP7_75t_L g2726 ( 
.A(n_2701),
.B(n_2598),
.Y(n_2726)
);

AND2x2_ASAP7_75t_L g2727 ( 
.A(n_2691),
.B(n_2647),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2680),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2700),
.B(n_2636),
.Y(n_2729)
);

INVx3_ASAP7_75t_L g2730 ( 
.A(n_2707),
.Y(n_2730)
);

INVx2_ASAP7_75t_SL g2731 ( 
.A(n_2707),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2700),
.B(n_2648),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_SL g2733 ( 
.A(n_2707),
.B(n_2604),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2678),
.B(n_2636),
.Y(n_2734)
);

OR2x2_ASAP7_75t_L g2735 ( 
.A(n_2681),
.B(n_2598),
.Y(n_2735)
);

OR2x2_ASAP7_75t_L g2736 ( 
.A(n_2681),
.B(n_2652),
.Y(n_2736)
);

AND2x2_ASAP7_75t_L g2737 ( 
.A(n_2698),
.B(n_2669),
.Y(n_2737)
);

AND2x2_ASAP7_75t_L g2738 ( 
.A(n_2698),
.B(n_2668),
.Y(n_2738)
);

AND2x2_ASAP7_75t_L g2739 ( 
.A(n_2706),
.B(n_2666),
.Y(n_2739)
);

INVx3_ASAP7_75t_L g2740 ( 
.A(n_2696),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2714),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2714),
.Y(n_2742)
);

AOI22xp5_ASAP7_75t_L g2743 ( 
.A1(n_2721),
.A2(n_2705),
.B1(n_2679),
.B2(n_2640),
.Y(n_2743)
);

OR2x2_ASAP7_75t_L g2744 ( 
.A(n_2735),
.B(n_2685),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2728),
.Y(n_2745)
);

A2O1A1Ixp33_ASAP7_75t_L g2746 ( 
.A1(n_2733),
.A2(n_2705),
.B(n_2663),
.C(n_2616),
.Y(n_2746)
);

OR2x2_ASAP7_75t_L g2747 ( 
.A(n_2735),
.B(n_2685),
.Y(n_2747)
);

OR2x2_ASAP7_75t_L g2748 ( 
.A(n_2726),
.B(n_2693),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2710),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2728),
.Y(n_2750)
);

OR2x2_ASAP7_75t_L g2751 ( 
.A(n_2726),
.B(n_2693),
.Y(n_2751)
);

NAND2x2_ASAP7_75t_L g2752 ( 
.A(n_2731),
.B(n_2529),
.Y(n_2752)
);

INVxp67_ASAP7_75t_L g2753 ( 
.A(n_2725),
.Y(n_2753)
);

OAI22xp5_ASAP7_75t_L g2754 ( 
.A1(n_2718),
.A2(n_2595),
.B1(n_2684),
.B2(n_2690),
.Y(n_2754)
);

AND2x4_ASAP7_75t_L g2755 ( 
.A(n_2718),
.B(n_2675),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2710),
.Y(n_2756)
);

OAI22xp5_ASAP7_75t_L g2757 ( 
.A1(n_2718),
.A2(n_2684),
.B1(n_2644),
.B2(n_2655),
.Y(n_2757)
);

AND2x4_ASAP7_75t_L g2758 ( 
.A(n_2718),
.B(n_2675),
.Y(n_2758)
);

INVx1_ASAP7_75t_SL g2759 ( 
.A(n_2724),
.Y(n_2759)
);

AOI22xp33_ASAP7_75t_L g2760 ( 
.A1(n_2736),
.A2(n_2679),
.B1(n_2618),
.B2(n_2678),
.Y(n_2760)
);

OR2x2_ASAP7_75t_L g2761 ( 
.A(n_2736),
.B(n_2692),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2709),
.B(n_2683),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2709),
.B(n_2686),
.Y(n_2763)
);

AOI22xp5_ASAP7_75t_L g2764 ( 
.A1(n_2718),
.A2(n_2485),
.B1(n_2657),
.B2(n_2627),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2732),
.B(n_2686),
.Y(n_2765)
);

AOI22xp33_ASAP7_75t_L g2766 ( 
.A1(n_2738),
.A2(n_2622),
.B1(n_2683),
.B2(n_2644),
.Y(n_2766)
);

INVx1_ASAP7_75t_SL g2767 ( 
.A(n_2724),
.Y(n_2767)
);

NOR2xp67_ASAP7_75t_L g2768 ( 
.A(n_2718),
.B(n_2655),
.Y(n_2768)
);

OAI21xp33_ASAP7_75t_L g2769 ( 
.A1(n_2715),
.A2(n_2688),
.B(n_2703),
.Y(n_2769)
);

HB1xp67_ASAP7_75t_L g2770 ( 
.A(n_2723),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2732),
.B(n_2694),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2712),
.Y(n_2772)
);

AND2x4_ASAP7_75t_L g2773 ( 
.A(n_2711),
.B(n_2675),
.Y(n_2773)
);

INVx2_ASAP7_75t_SL g2774 ( 
.A(n_2716),
.Y(n_2774)
);

INVxp67_ASAP7_75t_L g2775 ( 
.A(n_2716),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2715),
.B(n_2682),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2712),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2722),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2734),
.B(n_2694),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2717),
.B(n_2689),
.Y(n_2780)
);

OAI21xp33_ASAP7_75t_L g2781 ( 
.A1(n_2743),
.A2(n_2713),
.B(n_2739),
.Y(n_2781)
);

XOR2x2_ASAP7_75t_L g2782 ( 
.A(n_2743),
.B(n_2502),
.Y(n_2782)
);

INVx2_ASAP7_75t_SL g2783 ( 
.A(n_2752),
.Y(n_2783)
);

AOI22xp5_ASAP7_75t_L g2784 ( 
.A1(n_2754),
.A2(n_2739),
.B1(n_2719),
.B2(n_2717),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2741),
.Y(n_2785)
);

AOI22xp33_ASAP7_75t_SL g2786 ( 
.A1(n_2757),
.A2(n_2755),
.B1(n_2758),
.B2(n_2740),
.Y(n_2786)
);

NAND2xp33_ASAP7_75t_L g2787 ( 
.A(n_2746),
.B(n_2486),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2742),
.Y(n_2788)
);

AO22x1_ASAP7_75t_L g2789 ( 
.A1(n_2755),
.A2(n_2655),
.B1(n_2541),
.B2(n_2730),
.Y(n_2789)
);

AOI21xp33_ASAP7_75t_L g2790 ( 
.A1(n_2753),
.A2(n_2654),
.B(n_2671),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2778),
.Y(n_2791)
);

OAI22xp33_ASAP7_75t_L g2792 ( 
.A1(n_2764),
.A2(n_2768),
.B1(n_2774),
.B2(n_2730),
.Y(n_2792)
);

O2A1O1Ixp33_ASAP7_75t_L g2793 ( 
.A1(n_2770),
.A2(n_2653),
.B(n_2594),
.C(n_2713),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2749),
.Y(n_2794)
);

INVxp67_ASAP7_75t_L g2795 ( 
.A(n_2759),
.Y(n_2795)
);

OAI21xp5_ASAP7_75t_L g2796 ( 
.A1(n_2760),
.A2(n_2637),
.B(n_2731),
.Y(n_2796)
);

INVx1_ASAP7_75t_SL g2797 ( 
.A(n_2767),
.Y(n_2797)
);

NAND4xp25_ASAP7_75t_L g2798 ( 
.A(n_2766),
.B(n_2663),
.C(n_2509),
.D(n_2510),
.Y(n_2798)
);

OAI22xp33_ASAP7_75t_L g2799 ( 
.A1(n_2764),
.A2(n_2730),
.B1(n_2655),
.B2(n_2720),
.Y(n_2799)
);

OAI22xp5_ASAP7_75t_L g2800 ( 
.A1(n_2769),
.A2(n_2655),
.B1(n_2730),
.B2(n_2729),
.Y(n_2800)
);

OAI22xp5_ASAP7_75t_L g2801 ( 
.A1(n_2768),
.A2(n_2711),
.B1(n_2665),
.B2(n_2620),
.Y(n_2801)
);

INVxp67_ASAP7_75t_L g2802 ( 
.A(n_2761),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2745),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2756),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2802),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2785),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2797),
.Y(n_2807)
);

OAI21xp5_ASAP7_75t_SL g2808 ( 
.A1(n_2786),
.A2(n_2538),
.B(n_2493),
.Y(n_2808)
);

OAI21xp33_ASAP7_75t_L g2809 ( 
.A1(n_2784),
.A2(n_2775),
.B(n_2772),
.Y(n_2809)
);

NOR2xp33_ASAP7_75t_L g2810 ( 
.A(n_2783),
.B(n_2676),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2797),
.B(n_2762),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2788),
.Y(n_2812)
);

NOR2xp33_ASAP7_75t_L g2813 ( 
.A(n_2795),
.B(n_2508),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2803),
.B(n_2750),
.Y(n_2814)
);

AOI22xp5_ASAP7_75t_L g2815 ( 
.A1(n_2787),
.A2(n_2711),
.B1(n_2758),
.B2(n_2773),
.Y(n_2815)
);

AOI21xp33_ASAP7_75t_L g2816 ( 
.A1(n_2793),
.A2(n_2574),
.B(n_2495),
.Y(n_2816)
);

INVx2_ASAP7_75t_SL g2817 ( 
.A(n_2782),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2796),
.B(n_2773),
.Y(n_2818)
);

AND2x2_ASAP7_75t_SL g2819 ( 
.A(n_2789),
.B(n_2520),
.Y(n_2819)
);

AND2x4_ASAP7_75t_L g2820 ( 
.A(n_2794),
.B(n_2711),
.Y(n_2820)
);

OAI322xp33_ASAP7_75t_L g2821 ( 
.A1(n_2792),
.A2(n_2744),
.A3(n_2747),
.B1(n_2664),
.B2(n_2777),
.C1(n_2751),
.C2(n_2748),
.Y(n_2821)
);

OAI31xp33_ASAP7_75t_L g2822 ( 
.A1(n_2781),
.A2(n_2673),
.A3(n_2518),
.B(n_2349),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2804),
.Y(n_2823)
);

INVx2_ASAP7_75t_SL g2824 ( 
.A(n_2801),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2791),
.Y(n_2825)
);

OAI22xp33_ASAP7_75t_L g2826 ( 
.A1(n_2798),
.A2(n_2763),
.B1(n_2740),
.B2(n_2765),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2798),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2800),
.Y(n_2828)
);

NAND2xp33_ASAP7_75t_SL g2829 ( 
.A(n_2799),
.B(n_2474),
.Y(n_2829)
);

NOR2xp33_ASAP7_75t_L g2830 ( 
.A(n_2790),
.B(n_2530),
.Y(n_2830)
);

AOI22xp33_ASAP7_75t_SL g2831 ( 
.A1(n_2783),
.A2(n_2740),
.B1(n_2646),
.B2(n_2665),
.Y(n_2831)
);

NOR2x1_ASAP7_75t_L g2832 ( 
.A(n_2808),
.B(n_2827),
.Y(n_2832)
);

OAI21xp5_ASAP7_75t_L g2833 ( 
.A1(n_2808),
.A2(n_2480),
.B(n_2492),
.Y(n_2833)
);

NAND3xp33_ASAP7_75t_SL g2834 ( 
.A(n_2822),
.B(n_2513),
.C(n_2488),
.Y(n_2834)
);

NOR2xp67_ASAP7_75t_L g2835 ( 
.A(n_2824),
.B(n_2578),
.Y(n_2835)
);

NOR3xp33_ASAP7_75t_SL g2836 ( 
.A(n_2829),
.B(n_2470),
.C(n_2564),
.Y(n_2836)
);

NOR3xp33_ASAP7_75t_L g2837 ( 
.A(n_2817),
.B(n_2478),
.C(n_2463),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2807),
.B(n_2776),
.Y(n_2838)
);

INVx1_ASAP7_75t_SL g2839 ( 
.A(n_2819),
.Y(n_2839)
);

AOI21xp33_ASAP7_75t_L g2840 ( 
.A1(n_2813),
.A2(n_2659),
.B(n_2558),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2805),
.B(n_2738),
.Y(n_2841)
);

INVxp67_ASAP7_75t_SL g2842 ( 
.A(n_2810),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2811),
.Y(n_2843)
);

NOR3xp33_ASAP7_75t_SL g2844 ( 
.A(n_2826),
.B(n_2531),
.C(n_2559),
.Y(n_2844)
);

OAI21xp5_ASAP7_75t_SL g2845 ( 
.A1(n_2822),
.A2(n_2391),
.B(n_2638),
.Y(n_2845)
);

NAND3xp33_ASAP7_75t_L g2846 ( 
.A(n_2828),
.B(n_2592),
.C(n_2666),
.Y(n_2846)
);

AOI221xp5_ASAP7_75t_L g2847 ( 
.A1(n_2821),
.A2(n_2672),
.B1(n_2771),
.B2(n_2779),
.C(n_2740),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2806),
.B(n_2812),
.Y(n_2848)
);

AOI22xp5_ASAP7_75t_L g2849 ( 
.A1(n_2809),
.A2(n_2687),
.B1(n_2675),
.B2(n_2737),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2814),
.Y(n_2850)
);

NAND3xp33_ASAP7_75t_L g2851 ( 
.A(n_2832),
.B(n_2816),
.C(n_2830),
.Y(n_2851)
);

NOR3x1_ASAP7_75t_L g2852 ( 
.A(n_2834),
.B(n_2816),
.C(n_2823),
.Y(n_2852)
);

NAND3xp33_ASAP7_75t_L g2853 ( 
.A(n_2837),
.B(n_2831),
.C(n_2818),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2838),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2841),
.Y(n_2855)
);

AOI21xp5_ASAP7_75t_L g2856 ( 
.A1(n_2834),
.A2(n_2814),
.B(n_2815),
.Y(n_2856)
);

AOI22xp5_ASAP7_75t_L g2857 ( 
.A1(n_2842),
.A2(n_2835),
.B1(n_2839),
.B2(n_2845),
.Y(n_2857)
);

BUFx2_ASAP7_75t_L g2858 ( 
.A(n_2836),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2843),
.B(n_2825),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2848),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2850),
.Y(n_2861)
);

AND2x2_ASAP7_75t_L g2862 ( 
.A(n_2844),
.B(n_2847),
.Y(n_2862)
);

OAI21xp5_ASAP7_75t_L g2863 ( 
.A1(n_2846),
.A2(n_2820),
.B(n_2659),
.Y(n_2863)
);

INVx2_ASAP7_75t_SL g2864 ( 
.A(n_2849),
.Y(n_2864)
);

AOI21xp5_ASAP7_75t_SL g2865 ( 
.A1(n_2833),
.A2(n_2450),
.B(n_2504),
.Y(n_2865)
);

AOI22xp5_ASAP7_75t_L g2866 ( 
.A1(n_2840),
.A2(n_2820),
.B1(n_2450),
.B2(n_2504),
.Y(n_2866)
);

AOI222xp33_ASAP7_75t_L g2867 ( 
.A1(n_2851),
.A2(n_2621),
.B1(n_2623),
.B2(n_2613),
.C1(n_2607),
.C2(n_2606),
.Y(n_2867)
);

AOI221xp5_ASAP7_75t_L g2868 ( 
.A1(n_2860),
.A2(n_2473),
.B1(n_2611),
.B2(n_2629),
.C(n_2630),
.Y(n_2868)
);

AOI222xp33_ASAP7_75t_L g2869 ( 
.A1(n_2861),
.A2(n_2562),
.B1(n_2569),
.B2(n_2641),
.C1(n_2639),
.C2(n_2645),
.Y(n_2869)
);

OAI21xp5_ASAP7_75t_SL g2870 ( 
.A1(n_2858),
.A2(n_2550),
.B(n_2649),
.Y(n_2870)
);

OAI211xp5_ASAP7_75t_SL g2871 ( 
.A1(n_2857),
.A2(n_2588),
.B(n_2497),
.C(n_2372),
.Y(n_2871)
);

AO21x1_ASAP7_75t_L g2872 ( 
.A1(n_2856),
.A2(n_2586),
.B(n_2426),
.Y(n_2872)
);

NAND3xp33_ASAP7_75t_SL g2873 ( 
.A(n_2866),
.B(n_2539),
.C(n_2582),
.Y(n_2873)
);

NAND3xp33_ASAP7_75t_SL g2874 ( 
.A(n_2866),
.B(n_2853),
.C(n_2862),
.Y(n_2874)
);

NAND3xp33_ASAP7_75t_L g2875 ( 
.A(n_2859),
.B(n_2587),
.C(n_2397),
.Y(n_2875)
);

OAI211xp5_ASAP7_75t_L g2876 ( 
.A1(n_2865),
.A2(n_2662),
.B(n_2562),
.C(n_2372),
.Y(n_2876)
);

AOI22xp33_ASAP7_75t_L g2877 ( 
.A1(n_2864),
.A2(n_2687),
.B1(n_2696),
.B2(n_2662),
.Y(n_2877)
);

OAI211xp5_ASAP7_75t_SL g2878 ( 
.A1(n_2852),
.A2(n_2649),
.B(n_2395),
.C(n_2430),
.Y(n_2878)
);

OAI211xp5_ASAP7_75t_SL g2879 ( 
.A1(n_2855),
.A2(n_2649),
.B(n_2431),
.C(n_2428),
.Y(n_2879)
);

NOR2x1p5_ASAP7_75t_L g2880 ( 
.A(n_2874),
.B(n_2854),
.Y(n_2880)
);

AO22x2_ASAP7_75t_L g2881 ( 
.A1(n_2870),
.A2(n_2863),
.B1(n_2433),
.B2(n_2424),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2872),
.Y(n_2882)
);

AOI22xp5_ASAP7_75t_L g2883 ( 
.A1(n_2878),
.A2(n_2548),
.B1(n_2549),
.B2(n_2575),
.Y(n_2883)
);

AOI22xp33_ASAP7_75t_L g2884 ( 
.A1(n_2871),
.A2(n_2687),
.B1(n_2696),
.B2(n_2652),
.Y(n_2884)
);

NOR2x1p5_ASAP7_75t_L g2885 ( 
.A(n_2873),
.B(n_2293),
.Y(n_2885)
);

NOR2x1_ASAP7_75t_L g2886 ( 
.A(n_2875),
.B(n_2876),
.Y(n_2886)
);

INVxp33_ASAP7_75t_L g2887 ( 
.A(n_2868),
.Y(n_2887)
);

NOR2xp33_ASAP7_75t_L g2888 ( 
.A(n_2879),
.B(n_2642),
.Y(n_2888)
);

NOR2xp33_ASAP7_75t_L g2889 ( 
.A(n_2877),
.B(n_2632),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2867),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2880),
.B(n_2869),
.Y(n_2891)
);

AND2x4_ASAP7_75t_L g2892 ( 
.A(n_2885),
.B(n_2737),
.Y(n_2892)
);

OAI221xp5_ASAP7_75t_L g2893 ( 
.A1(n_2886),
.A2(n_2567),
.B1(n_2426),
.B2(n_2570),
.C(n_2573),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2882),
.Y(n_2894)
);

AND3x4_ASAP7_75t_L g2895 ( 
.A(n_2887),
.B(n_2571),
.C(n_2535),
.Y(n_2895)
);

AND2x2_ASAP7_75t_L g2896 ( 
.A(n_2881),
.B(n_2780),
.Y(n_2896)
);

AND2x2_ASAP7_75t_L g2897 ( 
.A(n_2889),
.B(n_2727),
.Y(n_2897)
);

AND2x2_ASAP7_75t_L g2898 ( 
.A(n_2890),
.B(n_2727),
.Y(n_2898)
);

NAND3xp33_ASAP7_75t_L g2899 ( 
.A(n_2888),
.B(n_2306),
.C(n_2293),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2883),
.Y(n_2900)
);

OAI22xp33_ASAP7_75t_L g2901 ( 
.A1(n_2884),
.A2(n_2567),
.B1(n_2573),
.B2(n_2570),
.Y(n_2901)
);

BUFx12f_ASAP7_75t_L g2902 ( 
.A(n_2892),
.Y(n_2902)
);

INVx1_ASAP7_75t_SL g2903 ( 
.A(n_2894),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2898),
.Y(n_2904)
);

INVx1_ASAP7_75t_SL g2905 ( 
.A(n_2891),
.Y(n_2905)
);

BUFx3_ASAP7_75t_L g2906 ( 
.A(n_2900),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2896),
.B(n_2633),
.Y(n_2907)
);

XNOR2xp5_ASAP7_75t_SL g2908 ( 
.A(n_2904),
.B(n_2895),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_2906),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2902),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2903),
.Y(n_2911)
);

XNOR2x1_ASAP7_75t_L g2912 ( 
.A(n_2905),
.B(n_2899),
.Y(n_2912)
);

AOI22xp5_ASAP7_75t_L g2913 ( 
.A1(n_2903),
.A2(n_2893),
.B1(n_2901),
.B2(n_2892),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2909),
.Y(n_2914)
);

AOI31xp33_ASAP7_75t_L g2915 ( 
.A1(n_2910),
.A2(n_2907),
.A3(n_2897),
.B(n_2386),
.Y(n_2915)
);

AOI211xp5_ASAP7_75t_L g2916 ( 
.A1(n_2911),
.A2(n_2293),
.B(n_2362),
.C(n_2306),
.Y(n_2916)
);

HB1xp67_ASAP7_75t_L g2917 ( 
.A(n_2914),
.Y(n_2917)
);

OAI21xp5_ASAP7_75t_L g2918 ( 
.A1(n_2915),
.A2(n_2908),
.B(n_2912),
.Y(n_2918)
);

OAI22xp5_ASAP7_75t_L g2919 ( 
.A1(n_2917),
.A2(n_2913),
.B1(n_2916),
.B2(n_2603),
.Y(n_2919)
);

OAI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2919),
.A2(n_2918),
.B(n_2441),
.Y(n_2920)
);

AOI22xp5_ASAP7_75t_L g2921 ( 
.A1(n_2920),
.A2(n_2306),
.B1(n_2362),
.B2(n_2571),
.Y(n_2921)
);

OR2x2_ASAP7_75t_L g2922 ( 
.A(n_2921),
.B(n_2584),
.Y(n_2922)
);

OAI22xp5_ASAP7_75t_L g2923 ( 
.A1(n_2922),
.A2(n_2362),
.B1(n_2584),
.B2(n_2603),
.Y(n_2923)
);


endmodule