module fake_ariane_2249_n_791 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_791);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_791;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_754;
wire n_336;
wire n_731;
wire n_779;
wire n_665;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_531;
wire n_783;
wire n_675;

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_41),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_88),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_56),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_110),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_8),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_4),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_150),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_106),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_25),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_11),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_49),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_121),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_122),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_118),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_46),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_156),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_60),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_125),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_57),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_95),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_44),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_130),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_86),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_76),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_141),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_43),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_34),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_152),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_63),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_148),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_27),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_37),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_97),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_51),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_133),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_73),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_52),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_102),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_45),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_11),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_128),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_89),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_155),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_74),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_26),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_31),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_80),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_19),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_42),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_66),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_17),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_82),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_109),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_77),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_87),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_220),
.Y(n_223)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_164),
.Y(n_230)
);

OAI21x1_ASAP7_75t_L g231 ( 
.A1(n_202),
.A2(n_221),
.B(n_213),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_163),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_163),
.A2(n_169),
.B1(n_217),
.B2(n_172),
.Y(n_234)
);

BUFx8_ASAP7_75t_SL g235 ( 
.A(n_169),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

BUFx8_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_166),
.Y(n_238)
);

CKINVDCx11_ASAP7_75t_R g239 ( 
.A(n_210),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_168),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_186),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_218),
.Y(n_245)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_165),
.B(n_0),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_192),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_195),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_198),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_200),
.B(n_0),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_201),
.B(n_1),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_205),
.Y(n_257)
);

OAI22x1_ASAP7_75t_SL g258 ( 
.A1(n_208),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_258)
);

AND2x4_ASAP7_75t_L g259 ( 
.A(n_212),
.B(n_215),
.Y(n_259)
);

AND2x4_ASAP7_75t_L g260 ( 
.A(n_170),
.B(n_2),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_171),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_173),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_174),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_175),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_176),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_177),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_225),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_235),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_222),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_235),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_239),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_239),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_232),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_245),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_R g275 ( 
.A(n_223),
.B(n_178),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_232),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_245),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_179),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_238),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_223),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_R g281 ( 
.A(n_244),
.B(n_180),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_236),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_R g283 ( 
.A(n_244),
.B(n_181),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_247),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_234),
.B(n_3),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_263),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_266),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_222),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_R g289 ( 
.A(n_246),
.B(n_182),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_227),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_247),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_266),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_225),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_247),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_260),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_222),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_253),
.B(n_184),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g298 ( 
.A1(n_231),
.A2(n_216),
.B(n_214),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_R g299 ( 
.A(n_246),
.B(n_185),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_226),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_266),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_266),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_222),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_246),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_247),
.Y(n_305)
);

INVx4_ASAP7_75t_SL g306 ( 
.A(n_248),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_248),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_R g308 ( 
.A(n_248),
.B(n_187),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_226),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_261),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_237),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_225),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_257),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_229),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_237),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_257),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_237),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_261),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_304),
.B(n_260),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_264),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_267),
.B(n_264),
.Y(n_321)
);

NOR3xp33_ASAP7_75t_L g322 ( 
.A(n_274),
.B(n_254),
.C(n_255),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_293),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_267),
.B(n_265),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_297),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_312),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_307),
.B(n_260),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_300),
.Y(n_328)
);

NAND3xp33_ASAP7_75t_L g329 ( 
.A(n_278),
.B(n_249),
.C(n_240),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_284),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_278),
.B(n_265),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_282),
.B(n_250),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_268),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_242),
.Y(n_335)
);

NOR2xp67_ASAP7_75t_SL g336 ( 
.A(n_286),
.B(n_254),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_309),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_279),
.Y(n_338)
);

NOR3xp33_ASAP7_75t_L g339 ( 
.A(n_277),
.B(n_256),
.C(n_252),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_229),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_287),
.B(n_259),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_292),
.B(n_259),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_295),
.B(n_259),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_294),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_290),
.B(n_251),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_301),
.B(n_302),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_295),
.B(n_257),
.Y(n_347)
);

NAND3xp33_ASAP7_75t_L g348 ( 
.A(n_305),
.B(n_257),
.C(n_230),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_313),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_275),
.B(n_252),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_273),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_L g352 ( 
.A(n_289),
.B(n_191),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_316),
.Y(n_353)
);

BUFx6f_ASAP7_75t_SL g354 ( 
.A(n_270),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_269),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_311),
.B(n_256),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_289),
.B(n_256),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_269),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_275),
.B(n_230),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_288),
.Y(n_360)
);

NOR3xp33_ASAP7_75t_L g361 ( 
.A(n_276),
.B(n_272),
.C(n_271),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_299),
.B(n_233),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_288),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_299),
.B(n_308),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_296),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_296),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_308),
.B(n_233),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_303),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_303),
.B(n_224),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_281),
.B(n_283),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_315),
.B(n_233),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_306),
.B(n_233),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_317),
.B(n_241),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_281),
.Y(n_374)
);

NOR2x1_ASAP7_75t_L g375 ( 
.A(n_280),
.B(n_241),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_298),
.Y(n_376)
);

BUFx5_ASAP7_75t_L g377 ( 
.A(n_306),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_306),
.B(n_241),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_283),
.B(n_241),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_285),
.A2(n_258),
.B1(n_243),
.B2(n_207),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_300),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_310),
.B(n_243),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_290),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_300),
.B(n_231),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_310),
.B(n_243),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_383),
.B(n_243),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_345),
.B(n_332),
.Y(n_387)
);

NAND3xp33_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_199),
.C(n_194),
.Y(n_388)
);

AND3x1_ASAP7_75t_L g389 ( 
.A(n_380),
.B(n_4),
.C(n_5),
.Y(n_389)
);

OR2x6_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_5),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_326),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_322),
.A2(n_203),
.B1(n_196),
.B2(n_211),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_338),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_344),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_350),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_334),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_335),
.B(n_193),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_323),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_364),
.B(n_197),
.Y(n_399)
);

NAND2x1p5_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_224),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_320),
.B(n_209),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_326),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_346),
.B(n_6),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_351),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_342),
.B(n_224),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_382),
.B(n_224),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_344),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_228),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_341),
.B(n_228),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_340),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_326),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_325),
.B(n_343),
.Y(n_412)
);

OAI22x1_ASAP7_75t_R g413 ( 
.A1(n_354),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_349),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_357),
.B(n_228),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_333),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_356),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_384),
.B(n_228),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_384),
.Y(n_420)
);

OR2x6_ASAP7_75t_L g421 ( 
.A(n_370),
.B(n_7),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_362),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_321),
.B(n_9),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_329),
.B(n_9),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_339),
.B(n_10),
.Y(n_425)
);

OR2x2_ASAP7_75t_SL g426 ( 
.A(n_380),
.B(n_10),
.Y(n_426)
);

OAI22x1_ASAP7_75t_L g427 ( 
.A1(n_328),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_324),
.B(n_12),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_353),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_359),
.B(n_319),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_355),
.Y(n_432)
);

INVx5_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_337),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_365),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_376),
.A2(n_91),
.B(n_160),
.Y(n_436)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_377),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_327),
.B(n_381),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_371),
.B(n_13),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_379),
.B(n_14),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_347),
.A2(n_92),
.B(n_159),
.Y(n_441)
);

OR2x6_ASAP7_75t_L g442 ( 
.A(n_373),
.B(n_15),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_358),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_336),
.B(n_15),
.Y(n_444)
);

A2O1A1Ixp33_ASAP7_75t_L g445 ( 
.A1(n_352),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_360),
.B(n_16),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_361),
.B(n_20),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_367),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_366),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_377),
.B(n_24),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_363),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_348),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_SL g453 ( 
.A(n_354),
.B(n_372),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_420),
.B(n_377),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_393),
.Y(n_455)
);

AOI33xp33_ASAP7_75t_L g456 ( 
.A1(n_387),
.A2(n_348),
.A3(n_368),
.B1(n_363),
.B2(n_369),
.B3(n_378),
.Y(n_456)
);

AOI21xp33_ASAP7_75t_L g457 ( 
.A1(n_418),
.A2(n_368),
.B(n_369),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_410),
.B(n_368),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_433),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_396),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_414),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_415),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_397),
.B(n_377),
.Y(n_463)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_404),
.Y(n_464)
);

AOI21x1_ASAP7_75t_L g465 ( 
.A1(n_419),
.A2(n_377),
.B(n_29),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_430),
.Y(n_466)
);

AOI21x1_ASAP7_75t_L g467 ( 
.A1(n_419),
.A2(n_28),
.B(n_30),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_432),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_434),
.B(n_32),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_433),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_403),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_471)
);

AOI221xp5_ASAP7_75t_L g472 ( 
.A1(n_389),
.A2(n_427),
.B1(n_438),
.B2(n_392),
.C(n_412),
.Y(n_472)
);

O2A1O1Ixp33_ASAP7_75t_L g473 ( 
.A1(n_424),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_473)
);

INVx6_ASAP7_75t_L g474 ( 
.A(n_386),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_395),
.B(n_412),
.Y(n_475)
);

OAI22x1_ASAP7_75t_L g476 ( 
.A1(n_447),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_476)
);

O2A1O1Ixp33_ASAP7_75t_L g477 ( 
.A1(n_425),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_423),
.A2(n_58),
.B(n_59),
.Y(n_478)
);

AOI31xp33_ASAP7_75t_L g479 ( 
.A1(n_389),
.A2(n_61),
.A3(n_62),
.B(n_64),
.Y(n_479)
);

O2A1O1Ixp33_ASAP7_75t_L g480 ( 
.A1(n_444),
.A2(n_429),
.B(n_445),
.C(n_399),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_433),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_449),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_439),
.B(n_65),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_409),
.A2(n_67),
.B(n_68),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_439),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_406),
.A2(n_69),
.B(n_70),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_401),
.B(n_71),
.Y(n_487)
);

O2A1O1Ixp33_ASAP7_75t_L g488 ( 
.A1(n_390),
.A2(n_72),
.B(n_75),
.C(n_78),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_431),
.B(n_442),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_422),
.B(n_79),
.Y(n_490)
);

NOR3xp33_ASAP7_75t_SL g491 ( 
.A(n_388),
.B(n_81),
.C(n_83),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_408),
.A2(n_84),
.B(n_85),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_442),
.B(n_90),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_417),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_405),
.A2(n_93),
.B(n_94),
.Y(n_495)
);

NAND2x1p5_ASAP7_75t_L g496 ( 
.A(n_394),
.B(n_96),
.Y(n_496)
);

AO31x2_ASAP7_75t_L g497 ( 
.A1(n_446),
.A2(n_98),
.A3(n_99),
.B(n_101),
.Y(n_497)
);

OR2x6_ASAP7_75t_L g498 ( 
.A(n_421),
.B(n_103),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_442),
.B(n_105),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_398),
.B(n_107),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_443),
.Y(n_501)
);

BUFx8_ASAP7_75t_SL g502 ( 
.A(n_421),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_421),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_394),
.B(n_108),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_435),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_447),
.B(n_111),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_426),
.B(n_112),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_437),
.A2(n_113),
.B(n_114),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_407),
.B(n_115),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_388),
.B(n_116),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_464),
.B(n_390),
.Y(n_511)
);

BUFx12f_ASAP7_75t_L g512 ( 
.A(n_498),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_455),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_481),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_472),
.B(n_390),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_480),
.A2(n_446),
.B(n_440),
.Y(n_516)
);

BUFx6f_ASAP7_75t_SL g517 ( 
.A(n_498),
.Y(n_517)
);

BUFx12f_ASAP7_75t_L g518 ( 
.A(n_503),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_481),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_461),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_459),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_474),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_463),
.A2(n_437),
.B(n_416),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_466),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_465),
.A2(n_436),
.B(n_448),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_478),
.A2(n_448),
.B(n_441),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_502),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_468),
.A2(n_391),
.B(n_411),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_507),
.Y(n_529)
);

INVx6_ASAP7_75t_L g530 ( 
.A(n_459),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_474),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_482),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_467),
.A2(n_450),
.B(n_402),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_459),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_504),
.A2(n_509),
.B(n_490),
.Y(n_535)
);

AO21x2_ASAP7_75t_L g536 ( 
.A1(n_500),
.A2(n_452),
.B(n_451),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_485),
.B(n_453),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_489),
.B(n_407),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_475),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_460),
.B(n_400),
.Y(n_540)
);

INVx8_ASAP7_75t_L g541 ( 
.A(n_470),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_501),
.Y(n_542)
);

AO21x2_ASAP7_75t_L g543 ( 
.A1(n_487),
.A2(n_428),
.B(n_400),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_475),
.B(n_428),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_493),
.B(n_413),
.Y(n_545)
);

AO21x2_ASAP7_75t_L g546 ( 
.A1(n_458),
.A2(n_117),
.B(n_119),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_470),
.Y(n_547)
);

BUFx2_ASAP7_75t_SL g548 ( 
.A(n_470),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_510),
.A2(n_454),
.B(n_483),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_496),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_462),
.Y(n_551)
);

BUFx8_ASAP7_75t_L g552 ( 
.A(n_506),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_505),
.Y(n_553)
);

BUFx2_ASAP7_75t_R g554 ( 
.A(n_479),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_506),
.Y(n_555)
);

OR2x6_ASAP7_75t_L g556 ( 
.A(n_499),
.B(n_161),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_513),
.Y(n_557)
);

BUFx2_ASAP7_75t_R g558 ( 
.A(n_527),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_551),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_520),
.Y(n_560)
);

BUFx4f_ASAP7_75t_SL g561 ( 
.A(n_512),
.Y(n_561)
);

OAI21x1_ASAP7_75t_L g562 ( 
.A1(n_525),
.A2(n_495),
.B(n_486),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_549),
.B(n_476),
.Y(n_563)
);

INVx6_ASAP7_75t_L g564 ( 
.A(n_552),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_551),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_547),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_539),
.Y(n_567)
);

NAND2x1p5_ASAP7_75t_L g568 ( 
.A(n_555),
.B(n_469),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_524),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_553),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_555),
.Y(n_571)
);

AOI21xp33_ASAP7_75t_L g572 ( 
.A1(n_515),
.A2(n_457),
.B(n_494),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_532),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_542),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_SL g575 ( 
.A1(n_529),
.A2(n_471),
.B1(n_491),
.B2(n_488),
.Y(n_575)
);

INVx4_ASAP7_75t_SL g576 ( 
.A(n_517),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_539),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_536),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_544),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_555),
.A2(n_477),
.B1(n_473),
.B2(n_508),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_547),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_530),
.Y(n_582)
);

AOI21x1_ASAP7_75t_L g583 ( 
.A1(n_535),
.A2(n_526),
.B(n_525),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_530),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_536),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_530),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_554),
.B(n_456),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_533),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_517),
.A2(n_484),
.B1(n_492),
.B2(n_497),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_533),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_547),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_531),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_527),
.Y(n_593)
);

CKINVDCx11_ASAP7_75t_R g594 ( 
.A(n_512),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_547),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_537),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_516),
.A2(n_497),
.B(n_124),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_546),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_531),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_R g600 ( 
.A(n_587),
.B(n_556),
.Y(n_600)
);

O2A1O1Ixp33_ASAP7_75t_SL g601 ( 
.A1(n_563),
.A2(n_519),
.B(n_514),
.C(n_550),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_557),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_575),
.A2(n_556),
.B1(n_538),
.B2(n_511),
.Y(n_603)
);

OAI21x1_ASAP7_75t_L g604 ( 
.A1(n_562),
.A2(n_535),
.B(n_526),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_R g605 ( 
.A(n_593),
.B(n_552),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_567),
.B(n_538),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_564),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_SL g608 ( 
.A1(n_587),
.A2(n_552),
.B1(n_545),
.B2(n_556),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_563),
.A2(n_518),
.B1(n_522),
.B2(n_528),
.Y(n_609)
);

AO31x2_ASAP7_75t_L g610 ( 
.A1(n_578),
.A2(n_523),
.A3(n_546),
.B(n_543),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_560),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_566),
.B(n_550),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_572),
.A2(n_518),
.B1(n_550),
.B2(n_543),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_569),
.Y(n_614)
);

NAND2x1_ASAP7_75t_L g615 ( 
.A(n_571),
.B(n_566),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_568),
.A2(n_514),
.B1(n_519),
.B2(n_521),
.Y(n_616)
);

OR2x6_ASAP7_75t_L g617 ( 
.A(n_564),
.B(n_548),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_SL g618 ( 
.A1(n_597),
.A2(n_540),
.B1(n_534),
.B2(n_521),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_576),
.B(n_534),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_573),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_570),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_592),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_592),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_568),
.A2(n_519),
.B1(n_514),
.B2(n_521),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_570),
.Y(n_625)
);

CKINVDCx16_ASAP7_75t_R g626 ( 
.A(n_593),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_577),
.B(n_534),
.Y(n_627)
);

CKINVDCx16_ASAP7_75t_R g628 ( 
.A(n_599),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_R g629 ( 
.A(n_596),
.B(n_123),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_R g630 ( 
.A(n_594),
.B(n_541),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_574),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_576),
.B(n_497),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_599),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_R g634 ( 
.A(n_594),
.B(n_561),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_582),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_R g636 ( 
.A(n_564),
.B(n_541),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_579),
.B(n_541),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_559),
.A2(n_565),
.B1(n_576),
.B2(n_571),
.Y(n_638)
);

OR2x2_ASAP7_75t_SL g639 ( 
.A(n_576),
.B(n_541),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_584),
.B(n_126),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_586),
.B(n_127),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_565),
.Y(n_642)
);

CKINVDCx16_ASAP7_75t_R g643 ( 
.A(n_558),
.Y(n_643)
);

NAND2xp33_ASAP7_75t_R g644 ( 
.A(n_591),
.B(n_129),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_R g645 ( 
.A(n_595),
.B(n_131),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_566),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_566),
.B(n_132),
.Y(n_647)
);

O2A1O1Ixp33_ASAP7_75t_SL g648 ( 
.A1(n_580),
.A2(n_135),
.B(n_136),
.C(n_137),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_602),
.B(n_590),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_611),
.B(n_590),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_606),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_614),
.B(n_581),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_621),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_627),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_615),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_620),
.B(n_588),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_631),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_642),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_625),
.B(n_588),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_632),
.B(n_628),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_632),
.B(n_583),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_635),
.B(n_581),
.Y(n_662)
);

OAI33xp33_ASAP7_75t_L g663 ( 
.A1(n_603),
.A2(n_585),
.A3(n_598),
.B1(n_589),
.B2(n_142),
.B3(n_143),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_622),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_610),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_623),
.B(n_581),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_633),
.B(n_581),
.Y(n_667)
);

INVx5_ASAP7_75t_L g668 ( 
.A(n_647),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_604),
.B(n_589),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_601),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_647),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_638),
.B(n_607),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_648),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_618),
.B(n_598),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_637),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_608),
.B(n_562),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_646),
.B(n_138),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_609),
.B(n_139),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_640),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_639),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_616),
.A2(n_140),
.B(n_144),
.Y(n_681)
);

NOR4xp25_ASAP7_75t_SL g682 ( 
.A(n_644),
.B(n_145),
.C(n_146),
.D(n_147),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_619),
.B(n_149),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_612),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_613),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_605),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_624),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_612),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_617),
.B(n_151),
.Y(n_689)
);

NOR2x1_ASAP7_75t_L g690 ( 
.A(n_670),
.B(n_617),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_651),
.B(n_654),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_657),
.B(n_626),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_653),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_675),
.B(n_612),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_660),
.B(n_641),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_661),
.B(n_676),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_661),
.B(n_643),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_662),
.B(n_630),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_662),
.B(n_634),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_660),
.B(n_600),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_676),
.B(n_636),
.Y(n_701)
);

INVxp67_ASAP7_75t_SL g702 ( 
.A(n_687),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_666),
.B(n_629),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_666),
.B(n_154),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_649),
.B(n_157),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_667),
.B(n_158),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_652),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_653),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_667),
.B(n_645),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_649),
.B(n_650),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_650),
.B(n_656),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_656),
.B(n_669),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_669),
.B(n_659),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_658),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_659),
.B(n_658),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_674),
.B(n_655),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_679),
.B(n_664),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_702),
.B(n_668),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_708),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_708),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_696),
.B(n_674),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_696),
.B(n_655),
.Y(n_722)
);

BUFx2_ASAP7_75t_SL g723 ( 
.A(n_697),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_712),
.B(n_670),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_714),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_712),
.B(n_672),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_697),
.B(n_686),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_714),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_710),
.B(n_680),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_710),
.B(n_685),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_716),
.B(n_680),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_711),
.B(n_685),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_720),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_719),
.Y(n_734)
);

NOR2x1p5_ASAP7_75t_L g735 ( 
.A(n_727),
.B(n_692),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_721),
.A2(n_716),
.B1(n_671),
.B2(n_672),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_723),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_728),
.Y(n_738)
);

OAI21xp33_ASAP7_75t_SL g739 ( 
.A1(n_724),
.A2(n_692),
.B(n_699),
.Y(n_739)
);

AOI32xp33_ASAP7_75t_L g740 ( 
.A1(n_721),
.A2(n_678),
.A3(n_673),
.B1(n_695),
.B2(n_677),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_722),
.B(n_711),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_739),
.A2(n_703),
.B1(n_709),
.B2(n_671),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_733),
.Y(n_743)
);

NOR3xp33_ASAP7_75t_L g744 ( 
.A(n_739),
.B(n_718),
.C(n_663),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_735),
.A2(n_678),
.B1(n_700),
.B2(n_679),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_734),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_737),
.A2(n_724),
.B1(n_718),
.B2(n_722),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_746),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_744),
.B(n_742),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_743),
.Y(n_750)
);

AOI21xp33_ASAP7_75t_SL g751 ( 
.A1(n_747),
.A2(n_740),
.B(n_691),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_745),
.B(n_726),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_749),
.A2(n_717),
.B(n_738),
.Y(n_753)
);

OAI21xp33_ASAP7_75t_L g754 ( 
.A1(n_751),
.A2(n_736),
.B(n_741),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_748),
.B(n_726),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_752),
.B(n_698),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_750),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_757),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_755),
.B(n_729),
.Y(n_759)
);

AOI221xp5_ASAP7_75t_SL g760 ( 
.A1(n_758),
.A2(n_754),
.B1(n_753),
.B2(n_756),
.C(n_673),
.Y(n_760)
);

AOI221xp5_ASAP7_75t_L g761 ( 
.A1(n_759),
.A2(n_693),
.B1(n_681),
.B2(n_695),
.C(n_707),
.Y(n_761)
);

OAI21xp33_ASAP7_75t_L g762 ( 
.A1(n_759),
.A2(n_694),
.B(n_690),
.Y(n_762)
);

AOI31xp33_ASAP7_75t_L g763 ( 
.A1(n_760),
.A2(n_677),
.A3(n_689),
.B(n_683),
.Y(n_763)
);

NOR3xp33_ASAP7_75t_L g764 ( 
.A(n_762),
.B(n_706),
.C(n_704),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_761),
.B(n_732),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_760),
.A2(n_695),
.B1(n_700),
.B2(n_701),
.Y(n_766)
);

INVxp33_ASAP7_75t_SL g767 ( 
.A(n_760),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_767),
.B(n_730),
.Y(n_768)
);

OAI221xp5_ASAP7_75t_SL g769 ( 
.A1(n_766),
.A2(n_701),
.B1(n_705),
.B2(n_688),
.C(n_684),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_765),
.Y(n_770)
);

NAND5xp2_ASAP7_75t_L g771 ( 
.A(n_763),
.B(n_764),
.C(n_705),
.D(n_689),
.E(n_713),
.Y(n_771)
);

AND2x2_ASAP7_75t_SL g772 ( 
.A(n_767),
.B(n_689),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_768),
.B(n_731),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_772),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_770),
.Y(n_775)
);

XOR2xp5_ASAP7_75t_L g776 ( 
.A(n_775),
.B(n_700),
.Y(n_776)
);

XOR2x2_ASAP7_75t_L g777 ( 
.A(n_774),
.B(n_769),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_773),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_778),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_L g780 ( 
.A1(n_777),
.A2(n_771),
.B1(n_668),
.B2(n_689),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_776),
.Y(n_781)
);

AO22x2_ASAP7_75t_L g782 ( 
.A1(n_779),
.A2(n_683),
.B1(n_731),
.B2(n_720),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_780),
.A2(n_668),
.B1(n_683),
.B2(n_682),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_781),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_779),
.A2(n_683),
.B1(n_668),
.B2(n_731),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_779),
.A2(n_668),
.B1(n_688),
.B2(n_684),
.Y(n_786)
);

XNOR2xp5_ASAP7_75t_L g787 ( 
.A(n_784),
.B(n_715),
.Y(n_787)
);

XNOR2xp5_ASAP7_75t_L g788 ( 
.A(n_787),
.B(n_783),
.Y(n_788)
);

AOI222xp33_ASAP7_75t_L g789 ( 
.A1(n_788),
.A2(n_782),
.B1(n_786),
.B2(n_785),
.C1(n_668),
.C2(n_725),
.Y(n_789)
);

OR2x6_ASAP7_75t_L g790 ( 
.A(n_789),
.B(n_725),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_790),
.A2(n_713),
.B1(n_715),
.B2(n_665),
.Y(n_791)
);


endmodule