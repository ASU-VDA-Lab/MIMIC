module fake_netlist_6_1653_n_1173 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_303, n_256, n_298, n_18, n_21, n_193, n_147, n_269, n_258, n_281, n_154, n_191, n_88, n_3, n_209, n_98, n_277, n_260, n_265, n_283, n_113, n_39, n_63, n_223, n_278, n_270, n_73, n_279, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_296, n_166, n_28, n_184, n_212, n_268, n_271, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_299, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_297, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_285, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_292, n_129, n_13, n_121, n_294, n_302, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_286, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_291, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_284, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_301, n_214, n_274, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_289, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_267, n_282, n_58, n_116, n_280, n_211, n_287, n_64, n_220, n_288, n_290, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_273, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_300, n_107, n_10, n_295, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_272, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_275, n_43, n_194, n_171, n_293, n_31, n_192, n_57, n_169, n_53, n_276, n_51, n_44, n_56, n_221, n_1173);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_303;
input n_256;
input n_298;
input n_18;
input n_21;
input n_193;
input n_147;
input n_269;
input n_258;
input n_281;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_277;
input n_260;
input n_265;
input n_283;
input n_113;
input n_39;
input n_63;
input n_223;
input n_278;
input n_270;
input n_73;
input n_279;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_296;
input n_166;
input n_28;
input n_184;
input n_212;
input n_268;
input n_271;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_299;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_297;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_285;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_292;
input n_129;
input n_13;
input n_121;
input n_294;
input n_302;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_286;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_291;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_284;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_301;
input n_214;
input n_274;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_289;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_267;
input n_282;
input n_58;
input n_116;
input n_280;
input n_211;
input n_287;
input n_64;
input n_220;
input n_288;
input n_290;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_273;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_300;
input n_107;
input n_10;
input n_295;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_272;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_275;
input n_43;
input n_194;
input n_171;
input n_293;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_276;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1173;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_760;
wire n_680;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_1079;
wire n_341;
wire n_362;
wire n_828;
wire n_462;
wire n_671;
wire n_607;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_1164;
wire n_310;
wire n_509;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1160;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_898;
wire n_617;
wire n_698;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_865;
wire n_1138;
wire n_893;
wire n_925;
wire n_485;
wire n_1101;
wire n_1026;
wire n_443;
wire n_1099;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_1139;
wire n_718;
wire n_517;
wire n_1018;
wire n_1172;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_742;
wire n_532;
wire n_535;
wire n_691;
wire n_901;
wire n_544;
wire n_372;
wire n_468;
wire n_1078;
wire n_504;
wire n_923;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_601;
wire n_375;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_1163;
wire n_1116;
wire n_611;
wire n_943;
wire n_1168;
wire n_491;
wire n_656;
wire n_843;
wire n_772;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_838;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_343;
wire n_886;
wire n_448;
wire n_953;
wire n_844;
wire n_1004;
wire n_1017;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_986;
wire n_839;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_870;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1148;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_1152;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_492;
wire n_972;
wire n_551;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_719;
wire n_565;
wire n_594;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_984;
wire n_818;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_981;
wire n_476;
wire n_880;
wire n_714;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_1110;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_409;
wire n_345;
wire n_689;
wire n_354;
wire n_799;
wire n_505;
wire n_1155;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_1051;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_1125;
wire n_970;
wire n_553;
wire n_652;
wire n_849;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_882;
wire n_811;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_1167;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_651;
wire n_404;
wire n_1153;
wire n_439;
wire n_518;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_1169;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_515;
wire n_983;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_1082;
wire n_1154;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_398;
wire n_410;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;

BUFx3_ASAP7_75t_L g304 ( 
.A(n_56),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_114),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_81),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_167),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_60),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_228),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_252),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_159),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_100),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_260),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_37),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_69),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_36),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_68),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_63),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_115),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_151),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_248),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_194),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_95),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_153),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_245),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_266),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_132),
.Y(n_327)
);

INVx4_ASAP7_75t_R g328 ( 
.A(n_21),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_164),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_102),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_123),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_273),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_30),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_82),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_196),
.Y(n_335)
);

BUFx8_ASAP7_75t_SL g336 ( 
.A(n_202),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_298),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_241),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_99),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_191),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_122),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_227),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_32),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_190),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_176),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_180),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_296),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_303),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_128),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_133),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_295),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_188),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_112),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_110),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_225),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_217),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_208),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_212),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_161),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_172),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_256),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_222),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_79),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_12),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_6),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_90),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_223),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_285),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_126),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_170),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_288),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_272),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_74),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_183),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_111),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_130),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_270),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_179),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_200),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_118),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_57),
.Y(n_381)
);

BUFx10_ASAP7_75t_L g382 ( 
.A(n_293),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_84),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_25),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_65),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_175),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_87),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_291),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_64),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_286),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_91),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_174),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_83),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_249),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_92),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_155),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_277),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_187),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_108),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_216),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_23),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_35),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_71),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_229),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_142),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_3),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_278),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_58),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_77),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_157),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_70),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_166),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_9),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_156),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_10),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_220),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_129),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_215),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_287),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_232),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_254),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_80),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_300),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_255),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_72),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_163),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_106),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_218),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_62),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_105),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_134),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_290),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_203),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_40),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_137),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_61),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_59),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_274),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_85),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_50),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_143),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_192),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_136),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_243),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_28),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_158),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_276),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_46),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_15),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_271),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_18),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_51),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_24),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_141),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_15),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_18),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_120),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_116),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_147),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_117),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_284),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_135),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_264),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_193),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_263),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_124),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_73),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_31),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_2),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_301),
.Y(n_470)
);

BUFx10_ASAP7_75t_L g471 ( 
.A(n_261),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_302),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_97),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_149),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_262),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_0),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_26),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_13),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_299),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_162),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_259),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_54),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_204),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_279),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_76),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_42),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_21),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_39),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_283),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_205),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_370),
.Y(n_491)
);

INVx5_ASAP7_75t_L g492 ( 
.A(n_370),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_309),
.B(n_0),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_393),
.B(n_1),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_382),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_370),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_413),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_398),
.B(n_1),
.Y(n_498)
);

BUFx8_ASAP7_75t_L g499 ( 
.A(n_445),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_382),
.B(n_471),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_455),
.Y(n_501)
);

BUFx12f_ASAP7_75t_L g502 ( 
.A(n_382),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_370),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_409),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_456),
.Y(n_505)
);

AND2x6_ASAP7_75t_L g506 ( 
.A(n_409),
.B(n_33),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_409),
.B(n_34),
.Y(n_507)
);

BUFx12f_ASAP7_75t_L g508 ( 
.A(n_471),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_409),
.Y(n_509)
);

BUFx8_ASAP7_75t_SL g510 ( 
.A(n_336),
.Y(n_510)
);

BUFx8_ASAP7_75t_L g511 ( 
.A(n_478),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_304),
.B(n_2),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_397),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_340),
.B(n_3),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_326),
.B(n_4),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_379),
.B(n_4),
.Y(n_516)
);

INVx5_ASAP7_75t_L g517 ( 
.A(n_471),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_304),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_327),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_397),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_434),
.B(n_5),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_428),
.B(n_5),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_327),
.B(n_6),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_340),
.B(n_7),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_352),
.B(n_7),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_352),
.Y(n_526)
);

INVx4_ASAP7_75t_L g527 ( 
.A(n_472),
.Y(n_527)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_472),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_428),
.B(n_8),
.Y(n_529)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_436),
.Y(n_530)
);

INVx5_ASAP7_75t_L g531 ( 
.A(n_436),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_438),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_438),
.Y(n_533)
);

CKINVDCx14_ASAP7_75t_R g534 ( 
.A(n_311),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_486),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_486),
.B(n_8),
.Y(n_536)
);

BUFx8_ASAP7_75t_SL g537 ( 
.A(n_451),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_333),
.B(n_9),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_364),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_365),
.B(n_10),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_316),
.B(n_11),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_308),
.Y(n_542)
);

BUFx8_ASAP7_75t_L g543 ( 
.A(n_312),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_313),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_344),
.B(n_11),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_384),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_330),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_401),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_406),
.B(n_12),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_415),
.B(n_13),
.Y(n_550)
);

INVx5_ASAP7_75t_L g551 ( 
.A(n_328),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_334),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_354),
.B(n_14),
.Y(n_553)
);

NOR2x1_ASAP7_75t_L g554 ( 
.A(n_337),
.B(n_14),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_342),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_347),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_305),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_348),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_349),
.B(n_16),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_372),
.B(n_16),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_350),
.Y(n_561)
);

BUFx12f_ASAP7_75t_L g562 ( 
.A(n_449),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_331),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_355),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_357),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_361),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_373),
.B(n_17),
.Y(n_567)
);

BUFx12f_ASAP7_75t_L g568 ( 
.A(n_453),
.Y(n_568)
);

AND2x6_ASAP7_75t_L g569 ( 
.A(n_403),
.B(n_38),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_468),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_469),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_306),
.Y(n_572)
);

BUFx8_ASAP7_75t_SL g573 ( 
.A(n_356),
.Y(n_573)
);

INVx5_ASAP7_75t_L g574 ( 
.A(n_476),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_477),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_307),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_487),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_366),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_368),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_377),
.B(n_17),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_310),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_466),
.B(n_19),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_483),
.B(n_380),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_383),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_385),
.B(n_391),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_394),
.Y(n_586)
);

INVx5_ASAP7_75t_L g587 ( 
.A(n_314),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_395),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_396),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_402),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_360),
.B(n_19),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_404),
.B(n_20),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_407),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_411),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_493),
.Y(n_595)
);

OR2x6_ASAP7_75t_L g596 ( 
.A(n_562),
.B(n_414),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_514),
.A2(n_399),
.B1(n_422),
.B2(n_378),
.Y(n_597)
);

OR2x6_ASAP7_75t_L g598 ( 
.A(n_568),
.B(n_418),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_503),
.Y(n_599)
);

AO22x2_ASAP7_75t_L g600 ( 
.A1(n_512),
.A2(n_423),
.B1(n_429),
.B2(n_421),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_500),
.A2(n_437),
.B1(n_424),
.B2(n_317),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_551),
.B(n_315),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_524),
.A2(n_319),
.B1(n_320),
.B2(n_318),
.Y(n_603)
);

OAI22xp33_ASAP7_75t_SL g604 ( 
.A1(n_494),
.A2(n_591),
.B1(n_521),
.B2(n_495),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_517),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_503),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_504),
.Y(n_607)
);

OA22x2_ASAP7_75t_L g608 ( 
.A1(n_590),
.A2(n_431),
.B1(n_442),
.B2(n_430),
.Y(n_608)
);

AO22x2_ASAP7_75t_L g609 ( 
.A1(n_512),
.A2(n_450),
.B1(n_462),
.B2(n_444),
.Y(n_609)
);

CKINVDCx6p67_ASAP7_75t_R g610 ( 
.A(n_502),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_557),
.B(n_467),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_504),
.Y(n_612)
);

AO22x2_ASAP7_75t_L g613 ( 
.A1(n_523),
.A2(n_481),
.B1(n_488),
.B2(n_479),
.Y(n_613)
);

OAI22xp33_ASAP7_75t_SL g614 ( 
.A1(n_495),
.A2(n_322),
.B1(n_323),
.B2(n_321),
.Y(n_614)
);

NAND3x1_ASAP7_75t_L g615 ( 
.A(n_554),
.B(n_20),
.C(n_22),
.Y(n_615)
);

OAI22xp33_ASAP7_75t_R g616 ( 
.A1(n_498),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_541),
.A2(n_490),
.B1(n_489),
.B2(n_485),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_551),
.B(n_324),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_509),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_509),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_496),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_582),
.A2(n_412),
.B1(n_482),
.B2(n_480),
.Y(n_622)
);

NAND2xp33_ASAP7_75t_SL g623 ( 
.A(n_525),
.B(n_325),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_572),
.B(n_329),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_496),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_519),
.B(n_332),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_553),
.A2(n_416),
.B1(n_475),
.B2(n_474),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_551),
.B(n_335),
.Y(n_628)
);

AOI22x1_ASAP7_75t_L g629 ( 
.A1(n_590),
.A2(n_585),
.B1(n_523),
.B2(n_588),
.Y(n_629)
);

OAI22xp33_ASAP7_75t_SL g630 ( 
.A1(n_550),
.A2(n_484),
.B1(n_473),
.B2(n_470),
.Y(n_630)
);

AND2x4_ASAP7_75t_SL g631 ( 
.A(n_563),
.B(n_338),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_519),
.B(n_465),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_560),
.A2(n_464),
.B1(n_463),
.B2(n_461),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_576),
.B(n_581),
.Y(n_634)
);

OAI22xp33_ASAP7_75t_L g635 ( 
.A1(n_545),
.A2(n_460),
.B1(n_459),
.B2(n_458),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_533),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_533),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_567),
.A2(n_457),
.B1(n_454),
.B2(n_452),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_535),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_535),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_497),
.Y(n_641)
);

OAI22xp33_ASAP7_75t_L g642 ( 
.A1(n_517),
.A2(n_516),
.B1(n_515),
.B2(n_522),
.Y(n_642)
);

OAI22xp33_ASAP7_75t_L g643 ( 
.A1(n_517),
.A2(n_448),
.B1(n_447),
.B2(n_446),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_542),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_571),
.B(n_339),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_548),
.B(n_341),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_519),
.B(n_343),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_574),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_583),
.B(n_539),
.Y(n_649)
);

AO22x2_ASAP7_75t_L g650 ( 
.A1(n_529),
.A2(n_536),
.B1(n_540),
.B2(n_538),
.Y(n_650)
);

NOR2x1p5_ASAP7_75t_L g651 ( 
.A(n_508),
.B(n_345),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_559),
.A2(n_443),
.B1(n_441),
.B2(n_440),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_539),
.B(n_346),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_580),
.A2(n_439),
.B1(n_435),
.B2(n_433),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_501),
.Y(n_655)
);

NAND2xp33_ASAP7_75t_SL g656 ( 
.A(n_549),
.B(n_351),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_526),
.Y(n_657)
);

AO22x2_ASAP7_75t_L g658 ( 
.A1(n_592),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_574),
.B(n_353),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_534),
.A2(n_388),
.B1(n_427),
.B2(n_426),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_572),
.B(n_358),
.Y(n_661)
);

OAI22xp33_ASAP7_75t_L g662 ( 
.A1(n_527),
.A2(n_432),
.B1(n_425),
.B2(n_420),
.Y(n_662)
);

OAI22xp33_ASAP7_75t_L g663 ( 
.A1(n_527),
.A2(n_419),
.B1(n_417),
.B2(n_410),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_573),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_546),
.B(n_27),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_546),
.B(n_570),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_558),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_561),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_570),
.A2(n_408),
.B1(n_405),
.B2(n_400),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_575),
.B(n_359),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_575),
.B(n_362),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_569),
.A2(n_376),
.B1(n_390),
.B2(n_389),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_564),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_578),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_544),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_636),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_637),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_640),
.Y(n_678)
);

XNOR2x2_ASAP7_75t_L g679 ( 
.A(n_658),
.B(n_554),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_666),
.B(n_587),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_631),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_657),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_649),
.A2(n_666),
.B(n_629),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_621),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_R g685 ( 
.A(n_646),
.B(n_363),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_606),
.Y(n_686)
);

CKINVDCx14_ASAP7_75t_R g687 ( 
.A(n_610),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_629),
.A2(n_589),
.B(n_566),
.Y(n_688)
);

INVxp67_ASAP7_75t_SL g689 ( 
.A(n_639),
.Y(n_689)
);

XOR2xp5_ASAP7_75t_L g690 ( 
.A(n_601),
.B(n_367),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_653),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_670),
.B(n_587),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_625),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_626),
.A2(n_566),
.B(n_520),
.Y(n_694)
);

NAND2xp33_ASAP7_75t_R g695 ( 
.A(n_634),
.B(n_369),
.Y(n_695)
);

XOR2xp5_ASAP7_75t_L g696 ( 
.A(n_660),
.B(n_371),
.Y(n_696)
);

AOI21x1_ASAP7_75t_L g697 ( 
.A1(n_671),
.A2(n_520),
.B(n_513),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_639),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_639),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_607),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_612),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_620),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_620),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_645),
.B(n_574),
.Y(n_704)
);

OAI21xp5_ASAP7_75t_L g705 ( 
.A1(n_608),
.A2(n_507),
.B(n_506),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_641),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_599),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_619),
.Y(n_708)
);

XOR2xp5_ASAP7_75t_L g709 ( 
.A(n_664),
.B(n_374),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_605),
.B(n_577),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_597),
.B(n_577),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_675),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_667),
.Y(n_713)
);

INVxp67_ASAP7_75t_SL g714 ( 
.A(n_655),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_669),
.B(n_587),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_668),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_673),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_644),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_634),
.B(n_577),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_627),
.B(n_518),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_656),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_602),
.B(n_528),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_674),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_623),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_611),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_611),
.Y(n_726)
);

INVxp33_ASAP7_75t_L g727 ( 
.A(n_665),
.Y(n_727)
);

NOR2xp67_ASAP7_75t_L g728 ( 
.A(n_633),
.B(n_528),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_600),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_595),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_600),
.Y(n_731)
);

XOR2xp5_ASAP7_75t_L g732 ( 
.A(n_672),
.B(n_375),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_609),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_618),
.B(n_628),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_595),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_638),
.B(n_518),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_609),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_613),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_648),
.B(n_528),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_613),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_632),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_622),
.B(n_544),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_647),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_624),
.B(n_661),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_650),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_603),
.B(n_547),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_650),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_642),
.B(n_530),
.Y(n_748)
);

NOR2xp67_ASAP7_75t_L g749 ( 
.A(n_652),
.B(n_491),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_615),
.Y(n_750)
);

OAI21xp33_ASAP7_75t_L g751 ( 
.A1(n_604),
.A2(n_505),
.B(n_513),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_659),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_658),
.Y(n_753)
);

INVx4_ASAP7_75t_SL g754 ( 
.A(n_596),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_654),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_630),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_614),
.Y(n_757)
);

NOR2xp67_ASAP7_75t_L g758 ( 
.A(n_662),
.B(n_491),
.Y(n_758)
);

INVxp67_ASAP7_75t_SL g759 ( 
.A(n_616),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_663),
.B(n_547),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_617),
.Y(n_761)
);

AND2x6_ASAP7_75t_L g762 ( 
.A(n_745),
.B(n_505),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_744),
.B(n_635),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_697),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_727),
.B(n_596),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_706),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_734),
.B(n_569),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_684),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_693),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_712),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_691),
.B(n_569),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_747),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_712),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_691),
.B(n_643),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_725),
.B(n_651),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_714),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_743),
.B(n_741),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_720),
.B(n_598),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_739),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_746),
.B(n_598),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_712),
.Y(n_781)
);

NAND2x1p5_ASAP7_75t_L g782 ( 
.A(n_724),
.B(n_491),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_714),
.B(n_506),
.Y(n_783)
);

AND2x2_ASAP7_75t_SL g784 ( 
.A(n_750),
.B(n_616),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_713),
.Y(n_785)
);

NAND2x1p5_ASAP7_75t_L g786 ( 
.A(n_752),
.B(n_492),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_719),
.Y(n_787)
);

AND2x2_ASAP7_75t_SL g788 ( 
.A(n_761),
.B(n_506),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_736),
.B(n_692),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_711),
.B(n_552),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_716),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_730),
.B(n_552),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_683),
.B(n_507),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_737),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_735),
.B(n_555),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_726),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_695),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_686),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_688),
.B(n_555),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_742),
.Y(n_800)
);

AND3x1_ASAP7_75t_SL g801 ( 
.A(n_729),
.B(n_733),
.C(n_731),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_683),
.B(n_507),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_755),
.B(n_530),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_688),
.B(n_556),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_682),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_738),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_717),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_718),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_723),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_704),
.B(n_556),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_740),
.B(n_565),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_760),
.B(n_381),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_756),
.B(n_386),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_680),
.B(n_676),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_722),
.B(n_530),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_705),
.A2(n_387),
.B(n_392),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_687),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_702),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_709),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_689),
.B(n_531),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_689),
.B(n_531),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_677),
.Y(n_822)
);

BUFx8_ASAP7_75t_L g823 ( 
.A(n_757),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_678),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_700),
.B(n_565),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_753),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_701),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_707),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_698),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_699),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_710),
.B(n_579),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_705),
.A2(n_492),
.B(n_531),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_751),
.B(n_579),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_753),
.Y(n_834)
);

INVx4_ASAP7_75t_L g835 ( 
.A(n_708),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_728),
.B(n_584),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_679),
.Y(n_837)
);

NOR2xp67_ASAP7_75t_R g838 ( 
.A(n_703),
.B(n_510),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_748),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_748),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_715),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_766),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_766),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_785),
.Y(n_844)
);

OR2x6_ASAP7_75t_L g845 ( 
.A(n_800),
.B(n_694),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_785),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_817),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_768),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_796),
.Y(n_849)
);

NAND2x1p5_ASAP7_75t_L g850 ( 
.A(n_770),
.B(n_758),
.Y(n_850)
);

NAND2x1p5_ASAP7_75t_L g851 ( 
.A(n_770),
.B(n_749),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_789),
.B(n_694),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_796),
.B(n_754),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_797),
.B(n_759),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_812),
.B(n_732),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_797),
.B(n_759),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_792),
.B(n_795),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_812),
.B(n_690),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_791),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_826),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_826),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_790),
.Y(n_862)
);

BUFx4f_ASAP7_75t_L g863 ( 
.A(n_839),
.Y(n_863)
);

INVx5_ASAP7_75t_L g864 ( 
.A(n_762),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_763),
.B(n_696),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_839),
.B(n_537),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_SL g867 ( 
.A(n_778),
.B(n_721),
.Y(n_867)
);

OR2x6_ASAP7_75t_L g868 ( 
.A(n_775),
.B(n_754),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_777),
.B(n_754),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_810),
.B(n_681),
.Y(n_870)
);

OR2x6_ASAP7_75t_L g871 ( 
.A(n_775),
.B(n_584),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_776),
.B(n_586),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_830),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_834),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_833),
.B(n_685),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_840),
.B(n_532),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_840),
.B(n_586),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_780),
.B(n_593),
.Y(n_878)
);

INVxp67_ASAP7_75t_L g879 ( 
.A(n_794),
.Y(n_879)
);

NAND2x1p5_ASAP7_75t_L g880 ( 
.A(n_773),
.B(n_492),
.Y(n_880)
);

OR2x6_ASAP7_75t_L g881 ( 
.A(n_839),
.B(n_593),
.Y(n_881)
);

AND2x2_ASAP7_75t_SL g882 ( 
.A(n_784),
.B(n_594),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_836),
.B(n_594),
.Y(n_883)
);

BUFx5_ASAP7_75t_L g884 ( 
.A(n_762),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_794),
.B(n_532),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_773),
.Y(n_886)
);

AND2x6_ASAP7_75t_L g887 ( 
.A(n_793),
.B(n_41),
.Y(n_887)
);

NAND2x1p5_ASAP7_75t_L g888 ( 
.A(n_781),
.B(n_532),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_768),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_769),
.Y(n_890)
);

BUFx4f_ASAP7_75t_L g891 ( 
.A(n_839),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_834),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_841),
.B(n_543),
.Y(n_893)
);

BUFx4_ASAP7_75t_SL g894 ( 
.A(n_868),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_848),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_886),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_861),
.Y(n_897)
);

BUFx12f_ASAP7_75t_L g898 ( 
.A(n_868),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_848),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_857),
.B(n_784),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_873),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_842),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_860),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_889),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_864),
.B(n_781),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_889),
.Y(n_906)
);

NAND2x1p5_ASAP7_75t_L g907 ( 
.A(n_864),
.B(n_828),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_849),
.B(n_853),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_892),
.Y(n_909)
);

BUFx4_ASAP7_75t_SL g910 ( 
.A(n_871),
.Y(n_910)
);

INVx1_ASAP7_75t_SL g911 ( 
.A(n_870),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_890),
.Y(n_912)
);

INVx5_ASAP7_75t_L g913 ( 
.A(n_864),
.Y(n_913)
);

INVx8_ASAP7_75t_L g914 ( 
.A(n_853),
.Y(n_914)
);

NAND2x1p5_ASAP7_75t_L g915 ( 
.A(n_863),
.B(n_828),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_863),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_847),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_842),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_886),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_890),
.Y(n_920)
);

NAND2x1p5_ASAP7_75t_L g921 ( 
.A(n_891),
.B(n_830),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_874),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_843),
.Y(n_923)
);

BUFx12f_ASAP7_75t_L g924 ( 
.A(n_871),
.Y(n_924)
);

BUFx4f_ASAP7_75t_L g925 ( 
.A(n_849),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_886),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_849),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_895),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_900),
.A2(n_855),
.B1(n_865),
.B2(n_858),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_920),
.A2(n_882),
.B1(n_837),
.B2(n_813),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_SL g931 ( 
.A1(n_911),
.A2(n_778),
.B(n_819),
.Y(n_931)
);

BUFx2_ASAP7_75t_SL g932 ( 
.A(n_903),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_899),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_SL g934 ( 
.A1(n_924),
.A2(n_837),
.B1(n_867),
.B2(n_823),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_917),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_920),
.Y(n_936)
);

BUFx10_ASAP7_75t_L g937 ( 
.A(n_917),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_923),
.A2(n_875),
.B1(n_854),
.B2(n_856),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_903),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_908),
.B(n_841),
.Y(n_940)
);

BUFx12f_ASAP7_75t_L g941 ( 
.A(n_924),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_904),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_916),
.A2(n_841),
.B1(n_891),
.B2(n_771),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_906),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_902),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_SL g946 ( 
.A1(n_909),
.A2(n_867),
.B1(n_823),
.B2(n_841),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_916),
.A2(n_850),
.B1(n_881),
.B2(n_767),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_912),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_925),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_902),
.Y(n_950)
);

INVxp67_ASAP7_75t_SL g951 ( 
.A(n_918),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_918),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_901),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_901),
.Y(n_954)
);

CKINVDCx11_ASAP7_75t_R g955 ( 
.A(n_898),
.Y(n_955)
);

BUFx8_ASAP7_75t_L g956 ( 
.A(n_898),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_915),
.A2(n_813),
.B1(n_816),
.B2(n_799),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_929),
.A2(n_866),
.B1(n_845),
.B2(n_878),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_928),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_929),
.A2(n_881),
.B1(n_909),
.B2(n_925),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_930),
.A2(n_804),
.B1(n_893),
.B2(n_845),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_930),
.A2(n_922),
.B1(n_774),
.B2(n_897),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_949),
.B(n_908),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_938),
.B(n_877),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_931),
.A2(n_915),
.B1(n_879),
.B2(n_862),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_936),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_935),
.Y(n_967)
);

INVx4_ASAP7_75t_L g968 ( 
.A(n_949),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_946),
.B(n_908),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_933),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_942),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_932),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_953),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_934),
.A2(n_946),
.B1(n_957),
.B2(n_762),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_944),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_948),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_SL g977 ( 
.A1(n_939),
.A2(n_765),
.B1(n_887),
.B2(n_788),
.Y(n_977)
);

OAI22xp33_ASAP7_75t_L g978 ( 
.A1(n_951),
.A2(n_940),
.B1(n_852),
.B2(n_950),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_934),
.B(n_885),
.Y(n_979)
);

HB1xp67_ASAP7_75t_SL g980 ( 
.A(n_956),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_957),
.A2(n_762),
.B1(n_835),
.B2(n_788),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_947),
.A2(n_762),
.B1(n_835),
.B2(n_809),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_937),
.B(n_927),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_937),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_951),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_943),
.A2(n_809),
.B1(n_887),
.B2(n_814),
.Y(n_986)
);

OAI22x1_ASAP7_75t_SL g987 ( 
.A1(n_955),
.A2(n_894),
.B1(n_910),
.B2(n_896),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_952),
.A2(n_887),
.B1(n_846),
.B2(n_844),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_956),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_945),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_954),
.B(n_806),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_941),
.A2(n_887),
.B1(n_769),
.B2(n_808),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_974),
.A2(n_543),
.B1(n_869),
.B2(n_791),
.Y(n_993)
);

NAND3xp33_ASAP7_75t_L g994 ( 
.A(n_958),
.B(n_511),
.C(n_499),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_979),
.A2(n_883),
.B1(n_831),
.B2(n_787),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_969),
.B(n_927),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_SL g997 ( 
.A1(n_960),
.A2(n_499),
.B1(n_511),
.B2(n_802),
.Y(n_997)
);

NAND3xp33_ASAP7_75t_SL g998 ( 
.A(n_974),
.B(n_851),
.C(n_803),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_961),
.A2(n_807),
.B1(n_827),
.B2(n_824),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_990),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_961),
.A2(n_807),
.B1(n_827),
.B2(n_824),
.Y(n_1001)
);

OAI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_964),
.A2(n_962),
.B1(n_985),
.B2(n_965),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_SL g1003 ( 
.A(n_967),
.B(n_896),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_SL g1004 ( 
.A1(n_984),
.A2(n_913),
.B1(n_884),
.B2(n_782),
.Y(n_1004)
);

OAI211xp5_ASAP7_75t_L g1005 ( 
.A1(n_977),
.A2(n_772),
.B(n_811),
.C(n_805),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_985),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_981),
.A2(n_822),
.B1(n_859),
.B2(n_872),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_963),
.A2(n_825),
.B1(n_818),
.B2(n_914),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_959),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_990),
.B(n_772),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_966),
.B(n_919),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_970),
.B(n_919),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_SL g1013 ( 
.A1(n_984),
.A2(n_972),
.B1(n_968),
.B2(n_983),
.Y(n_1013)
);

OAI221xp5_ASAP7_75t_L g1014 ( 
.A1(n_982),
.A2(n_782),
.B1(n_786),
.B2(n_779),
.C(n_822),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_SL g1015 ( 
.A1(n_992),
.A2(n_910),
.B(n_832),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_986),
.A2(n_798),
.B1(n_830),
.B2(n_884),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_SL g1017 ( 
.A1(n_984),
.A2(n_913),
.B1(n_884),
.B2(n_914),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_984),
.A2(n_798),
.B1(n_830),
.B2(n_884),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_963),
.A2(n_798),
.B1(n_884),
.B2(n_829),
.Y(n_1019)
);

OAI222xp33_ASAP7_75t_L g1020 ( 
.A1(n_980),
.A2(n_921),
.B1(n_876),
.B2(n_907),
.C1(n_905),
.C2(n_786),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_991),
.Y(n_1021)
);

INVxp67_ASAP7_75t_SL g1022 ( 
.A(n_978),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_968),
.A2(n_798),
.B1(n_926),
.B2(n_876),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_971),
.Y(n_1024)
);

AOI221xp5_ASAP7_75t_L g1025 ( 
.A1(n_978),
.A2(n_806),
.B1(n_914),
.B2(n_783),
.C(n_815),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_973),
.A2(n_926),
.B1(n_873),
.B2(n_921),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_988),
.A2(n_907),
.B1(n_913),
.B2(n_905),
.Y(n_1027)
);

OAI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_975),
.A2(n_913),
.B1(n_926),
.B2(n_894),
.Y(n_1028)
);

NAND3xp33_ASAP7_75t_L g1029 ( 
.A(n_988),
.B(n_926),
.C(n_821),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_976),
.A2(n_764),
.B1(n_888),
.B2(n_30),
.Y(n_1030)
);

NAND4xp25_ASAP7_75t_L g1031 ( 
.A(n_994),
.B(n_973),
.C(n_838),
.D(n_801),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_996),
.B(n_28),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_1021),
.B(n_29),
.Y(n_1033)
);

NAND3xp33_ASAP7_75t_L g1034 ( 
.A(n_997),
.B(n_989),
.C(n_820),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_SL g1035 ( 
.A1(n_1005),
.A2(n_987),
.B(n_880),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1000),
.B(n_29),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1009),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1002),
.B(n_1022),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1002),
.B(n_31),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_SL g1040 ( 
.A(n_1003),
.B(n_764),
.Y(n_1040)
);

NAND3xp33_ASAP7_75t_L g1041 ( 
.A(n_1030),
.B(n_801),
.C(n_44),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1024),
.B(n_43),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1006),
.B(n_45),
.Y(n_1043)
);

OAI221xp5_ASAP7_75t_SL g1044 ( 
.A1(n_1015),
.A2(n_1030),
.B1(n_993),
.B2(n_995),
.C(n_1025),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1013),
.B(n_47),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1012),
.B(n_48),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1011),
.B(n_49),
.Y(n_1047)
);

OA211x2_ASAP7_75t_L g1048 ( 
.A1(n_998),
.A2(n_52),
.B(n_53),
.C(n_55),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1010),
.B(n_66),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1028),
.B(n_67),
.Y(n_1050)
);

OAI221xp5_ASAP7_75t_L g1051 ( 
.A1(n_1008),
.A2(n_75),
.B1(n_78),
.B2(n_86),
.C(n_88),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_1028),
.A2(n_89),
.B1(n_93),
.B2(n_94),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_999),
.B(n_96),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_SL g1054 ( 
.A1(n_1020),
.A2(n_98),
.B(n_101),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_1001),
.A2(n_103),
.B1(n_104),
.B2(n_107),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_SL g1056 ( 
.A1(n_1004),
.A2(n_109),
.B(n_113),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_SL g1057 ( 
.A(n_1014),
.B(n_119),
.Y(n_1057)
);

AOI221xp5_ASAP7_75t_L g1058 ( 
.A1(n_1029),
.A2(n_121),
.B1(n_125),
.B2(n_127),
.C(n_131),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1026),
.B(n_1007),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_1017),
.B(n_138),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1027),
.A2(n_139),
.B(n_140),
.Y(n_1061)
);

AOI221xp5_ASAP7_75t_L g1062 ( 
.A1(n_1039),
.A2(n_1023),
.B1(n_1016),
.B2(n_1019),
.C(n_1018),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1037),
.B(n_144),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_1038),
.B(n_145),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1032),
.B(n_146),
.Y(n_1065)
);

AO21x2_ASAP7_75t_L g1066 ( 
.A1(n_1035),
.A2(n_148),
.B(n_150),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1036),
.B(n_152),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1043),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_SL g1069 ( 
.A1(n_1034),
.A2(n_154),
.B1(n_160),
.B2(n_165),
.Y(n_1069)
);

NAND3xp33_ASAP7_75t_L g1070 ( 
.A(n_1044),
.B(n_168),
.C(n_169),
.Y(n_1070)
);

NOR3xp33_ASAP7_75t_L g1071 ( 
.A(n_1054),
.B(n_171),
.C(n_173),
.Y(n_1071)
);

OAI211xp5_ASAP7_75t_L g1072 ( 
.A1(n_1035),
.A2(n_177),
.B(n_178),
.C(n_181),
.Y(n_1072)
);

AO21x2_ASAP7_75t_L g1073 ( 
.A1(n_1060),
.A2(n_182),
.B(n_184),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1033),
.B(n_185),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1042),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1049),
.B(n_186),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_1059),
.B(n_189),
.Y(n_1077)
);

OAI211xp5_ASAP7_75t_SL g1078 ( 
.A1(n_1058),
.A2(n_1046),
.B(n_1050),
.C(n_1051),
.Y(n_1078)
);

NAND3xp33_ASAP7_75t_L g1079 ( 
.A(n_1041),
.B(n_195),
.C(n_197),
.Y(n_1079)
);

OAI211xp5_ASAP7_75t_SL g1080 ( 
.A1(n_1056),
.A2(n_198),
.B(n_199),
.C(n_201),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1057),
.A2(n_206),
.B(n_207),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_1047),
.Y(n_1082)
);

NOR3xp33_ASAP7_75t_SL g1083 ( 
.A(n_1031),
.B(n_297),
.C(n_210),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1075),
.B(n_1045),
.Y(n_1084)
);

NAND4xp75_ASAP7_75t_L g1085 ( 
.A(n_1081),
.B(n_1048),
.C(n_1060),
.D(n_1061),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1082),
.B(n_1040),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_1068),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_1067),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_SL g1089 ( 
.A(n_1070),
.B(n_1078),
.C(n_1072),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1063),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_1063),
.B(n_1052),
.Y(n_1091)
);

NOR3xp33_ASAP7_75t_SL g1092 ( 
.A(n_1080),
.B(n_1081),
.C(n_1064),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1067),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1074),
.B(n_1053),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1077),
.B(n_1055),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1073),
.B(n_1055),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_1065),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1066),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_1076),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_1066),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1073),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1071),
.A2(n_209),
.B1(n_211),
.B2(n_213),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1083),
.B(n_214),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_1087),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1093),
.B(n_1062),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1087),
.Y(n_1106)
);

INVxp67_ASAP7_75t_SL g1107 ( 
.A(n_1100),
.Y(n_1107)
);

INVxp67_ASAP7_75t_L g1108 ( 
.A(n_1100),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1088),
.B(n_1069),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1090),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1101),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1101),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1098),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1089),
.A2(n_1085),
.B1(n_1092),
.B2(n_1102),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1097),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1084),
.B(n_1079),
.Y(n_1116)
);

XOR2x2_ASAP7_75t_L g1117 ( 
.A(n_1099),
.B(n_219),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1086),
.B(n_221),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_1096),
.B(n_224),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1091),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1094),
.Y(n_1121)
);

XNOR2x1_ASAP7_75t_L g1122 ( 
.A(n_1095),
.B(n_226),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1113),
.Y(n_1123)
);

OA22x2_ASAP7_75t_L g1124 ( 
.A1(n_1114),
.A2(n_1103),
.B1(n_1089),
.B2(n_1092),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1106),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1110),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1111),
.Y(n_1127)
);

OA22x2_ASAP7_75t_L g1128 ( 
.A1(n_1105),
.A2(n_230),
.B1(n_231),
.B2(n_233),
.Y(n_1128)
);

XNOR2xp5_ASAP7_75t_L g1129 ( 
.A(n_1122),
.B(n_234),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_SL g1130 ( 
.A(n_1120),
.B(n_235),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1105),
.B(n_236),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1115),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1104),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_1117),
.Y(n_1134)
);

OA22x2_ASAP7_75t_L g1135 ( 
.A1(n_1109),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_1121),
.Y(n_1136)
);

OA22x2_ASAP7_75t_L g1137 ( 
.A1(n_1116),
.A2(n_240),
.B1(n_242),
.B2(n_244),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1107),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1112),
.Y(n_1139)
);

INVx6_ASAP7_75t_L g1140 ( 
.A(n_1118),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1126),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1123),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1123),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1138),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1133),
.Y(n_1145)
);

OAI22x1_ASAP7_75t_SL g1146 ( 
.A1(n_1145),
.A2(n_1134),
.B1(n_1133),
.B2(n_1124),
.Y(n_1146)
);

OAI22x1_ASAP7_75t_L g1147 ( 
.A1(n_1144),
.A2(n_1129),
.B1(n_1107),
.B2(n_1132),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1144),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1141),
.A2(n_1128),
.B1(n_1135),
.B2(n_1137),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_1142),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1149),
.A2(n_1131),
.B(n_1108),
.C(n_1116),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1146),
.A2(n_1147),
.B1(n_1129),
.B2(n_1150),
.Y(n_1152)
);

OAI22x1_ASAP7_75t_L g1153 ( 
.A1(n_1148),
.A2(n_1143),
.B1(n_1108),
.B2(n_1138),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1149),
.A2(n_1140),
.B1(n_1136),
.B2(n_1119),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1153),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1152),
.A2(n_1140),
.B1(n_1125),
.B2(n_1139),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1154),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1151),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_1155),
.Y(n_1159)
);

NOR2x1_ASAP7_75t_L g1160 ( 
.A(n_1158),
.B(n_1127),
.Y(n_1160)
);

AND4x1_ASAP7_75t_L g1161 ( 
.A(n_1160),
.B(n_1157),
.C(n_1130),
.D(n_1159),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1161),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1162),
.A2(n_1156),
.B1(n_247),
.B2(n_250),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1162),
.A2(n_246),
.B1(n_251),
.B2(n_253),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1163),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1165),
.A2(n_1164),
.B1(n_258),
.B2(n_265),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1166),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1166),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1167),
.A2(n_257),
.B1(n_267),
.B2(n_268),
.Y(n_1169)
);

OAI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1168),
.A2(n_269),
.B1(n_275),
.B2(n_280),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1169),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1171),
.A2(n_1170),
.B1(n_282),
.B2(n_289),
.Y(n_1172)
);

AOI211xp5_ASAP7_75t_L g1173 ( 
.A1(n_1172),
.A2(n_281),
.B(n_292),
.C(n_294),
.Y(n_1173)
);


endmodule