module fake_jpeg_8595_n_285 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_285);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx4f_ASAP7_75t_SL g14 ( 
.A(n_8),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_1),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_48),
.Y(n_64)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

OR2x2_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_14),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_66),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_55),
.A2(n_26),
.B1(n_24),
.B2(n_17),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_20),
.B(n_19),
.Y(n_94)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_65),
.Y(n_82)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_18),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_15),
.B1(n_26),
.B2(n_17),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_16),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_71),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_39),
.A2(n_24),
.B(n_15),
.C(n_23),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_15),
.B1(n_23),
.B2(n_21),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_74),
.B1(n_20),
.B2(n_41),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_75),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_41),
.A2(n_22),
.B1(n_29),
.B2(n_21),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g77 ( 
.A(n_45),
.Y(n_77)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_63),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_80),
.A2(n_89),
.B1(n_59),
.B2(n_73),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_64),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_87),
.B(n_90),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_68),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_92),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_43),
.Y(n_92)
);

AO21x1_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_19),
.B(n_25),
.Y(n_121)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_22),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_51),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_74),
.C(n_77),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_105),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_71),
.B(n_60),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_103),
.A2(n_43),
.B(n_46),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_59),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_77),
.C(n_35),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_108),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_88),
.C(n_98),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_49),
.C(n_48),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_112),
.B(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_118),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_92),
.B(n_83),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_81),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_119),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_121),
.A2(n_90),
.B(n_91),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_83),
.B(n_92),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_134),
.B(n_136),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_120),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_129),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_120),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_130),
.A2(n_135),
.B1(n_140),
.B2(n_143),
.Y(n_168)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_132),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_104),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_19),
.B(n_13),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_61),
.B1(n_65),
.B2(n_95),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_137),
.A2(n_73),
.B1(n_109),
.B2(n_86),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_115),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_141),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_121),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_16),
.Y(n_160)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_100),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_81),
.B1(n_117),
.B2(n_107),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_122),
.B1(n_101),
.B2(n_103),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_147),
.A2(n_50),
.B1(n_51),
.B2(n_76),
.Y(n_192)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_110),
.C(n_117),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_159),
.Y(n_180)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_155),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_162),
.B(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_113),
.C(n_107),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_146),
.B(n_134),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_130),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_163),
.A2(n_145),
.B1(n_140),
.B2(n_109),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_131),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_164),
.B(n_170),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_16),
.Y(n_165)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_78),
.Y(n_169)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_141),
.B(n_97),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_1),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_171),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_187),
.B1(n_190),
.B2(n_150),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_173),
.A2(n_19),
.B(n_13),
.Y(n_205)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_133),
.C(n_142),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_172),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_177),
.A2(n_126),
.B1(n_47),
.B2(n_62),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_152),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_183),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_153),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_161),
.Y(n_184)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_151),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_133),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_40),
.Y(n_206)
);

NOR2x1_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_139),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_160),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_171),
.B(n_167),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_193),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_148),
.A2(n_97),
.B1(n_126),
.B2(n_102),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_194),
.A2(n_156),
.B1(n_159),
.B2(n_165),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_187),
.B(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_188),
.B(n_147),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_205),
.Y(n_218)
);

AOI21xp33_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_178),
.B(n_176),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_201),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_162),
.B1(n_163),
.B2(n_155),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_202),
.A2(n_207),
.B1(n_177),
.B2(n_62),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_203),
.A2(n_212),
.B1(n_193),
.B2(n_185),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_208),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_126),
.B1(n_99),
.B2(n_47),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_173),
.B(n_13),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_179),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_179),
.Y(n_213)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_180),
.C(n_191),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_220),
.C(n_224),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_215),
.A2(n_221),
.B(n_9),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_228),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_180),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_182),
.B1(n_191),
.B2(n_178),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_190),
.C(n_194),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_199),
.C(n_209),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_7),
.C(n_12),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_207),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_1),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_222),
.A2(n_196),
.B1(n_210),
.B2(n_195),
.Y(n_231)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_226),
.A2(n_196),
.B(n_201),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_232),
.A2(n_239),
.B(n_240),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_208),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_243),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_219),
.B(n_8),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_235),
.B(n_236),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_214),
.B(n_9),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_237),
.B(n_11),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_229),
.A2(n_70),
.B(n_7),
.Y(n_239)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_230),
.A2(n_1),
.B(n_2),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_223),
.C(n_217),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_221),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_216),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_6),
.B(n_11),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_241),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_247),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_225),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_244),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_254),
.Y(n_261)
);

INVx11_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_256),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_238),
.C(n_220),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_258),
.C(n_262),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_218),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_225),
.Y(n_259)
);

OAI211xp5_ASAP7_75t_SL g272 ( 
.A1(n_259),
.A2(n_4),
.B(n_5),
.C(n_10),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_249),
.A2(n_56),
.B(n_53),
.Y(n_265)
);

AO21x1_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_266),
.B(n_4),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_4),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_260),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_269),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_263),
.A2(n_255),
.B1(n_253),
.B2(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_268),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_253),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_246),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_271),
.B(n_272),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_258),
.Y(n_274)
);

NAND4xp25_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_267),
.C(n_259),
.D(n_270),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);

AOI322xp5_ASAP7_75t_L g280 ( 
.A1(n_278),
.A2(n_279),
.A3(n_276),
.B1(n_264),
.B2(n_275),
.C1(n_10),
.C2(n_5),
.Y(n_280)
);

OAI21x1_ASAP7_75t_L g281 ( 
.A1(n_280),
.A2(n_10),
.B(n_2),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_281),
.A2(n_2),
.B(n_3),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_282),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_3),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_3),
.B(n_246),
.Y(n_285)
);


endmodule