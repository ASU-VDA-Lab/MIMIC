module fake_jpeg_19092_n_215 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_215);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_15),
.B1(n_14),
.B2(n_30),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_49),
.B1(n_54),
.B2(n_16),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_15),
.B1(n_14),
.B2(n_30),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_31),
.A2(n_15),
.B1(n_30),
.B2(n_17),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_69),
.B1(n_70),
.B2(n_86),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_39),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_56),
.A2(n_57),
.B(n_74),
.Y(n_92)
);

OR2x6_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_58),
.B(n_71),
.Y(n_104)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_24),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_61),
.B(n_66),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_46),
.B(n_20),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_74),
.C(n_55),
.Y(n_99)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_19),
.C(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_24),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_75),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_34),
.B1(n_23),
.B2(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_26),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_22),
.B1(n_17),
.B2(n_21),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_79),
.B1(n_20),
.B2(n_3),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_34),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_84),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_27),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_77),
.B(n_80),
.Y(n_110)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_40),
.A2(n_22),
.B1(n_17),
.B2(n_21),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_85),
.Y(n_91)
);

NOR2xp67_ASAP7_75t_R g83 ( 
.A(n_49),
.B(n_29),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_87),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_29),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_54),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_28),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_28),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_88),
.B(n_94),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_59),
.Y(n_94)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_27),
.C(n_20),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_99),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_26),
.B1(n_22),
.B2(n_21),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_100),
.A2(n_101),
.B1(n_103),
.B2(n_106),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_16),
.B1(n_28),
.B2(n_18),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_69),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_28),
.B1(n_2),
.B2(n_3),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_109),
.B1(n_62),
.B2(n_56),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_106),
.A2(n_108),
.B(n_100),
.Y(n_122)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_81),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_109)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_89),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_62),
.C(n_82),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_127),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_129),
.B1(n_132),
.B2(n_134),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_58),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_94),
.B(n_93),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_92),
.A2(n_56),
.B(n_74),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_101),
.B(n_109),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_71),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_128),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_76),
.B(n_64),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_126),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_92),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_78),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_65),
.B1(n_73),
.B2(n_68),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_98),
.A2(n_65),
.B1(n_73),
.B2(n_68),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_91),
.A2(n_60),
.B1(n_5),
.B2(n_6),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_60),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_SL g157 ( 
.A(n_135),
.B(n_97),
.C(n_112),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_88),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_137),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_63),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_132),
.B1(n_120),
.B2(n_126),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_144),
.B1(n_107),
.B2(n_113),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_105),
.B1(n_102),
.B2(n_103),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_91),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_147),
.Y(n_174)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_111),
.C(n_108),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_152),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_119),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_150),
.B(n_133),
.Y(n_166)
);

NAND2xp33_ASAP7_75t_SL g160 ( 
.A(n_151),
.B(n_157),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_97),
.B(n_60),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_118),
.Y(n_158)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

OAI321xp33_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_125),
.A3(n_128),
.B1(n_127),
.B2(n_117),
.C(n_131),
.Y(n_159)
);

OAI321xp33_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_148),
.A3(n_145),
.B1(n_140),
.B2(n_9),
.C(n_10),
.Y(n_186)
);

INVxp33_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_173),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_115),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_164),
.B(n_170),
.Y(n_176)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_167),
.Y(n_179)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_125),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_171),
.Y(n_182)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_172),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_141),
.B(n_130),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_116),
.C(n_113),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_139),
.B1(n_143),
.B2(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_160),
.A2(n_144),
.B1(n_139),
.B2(n_138),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_163),
.B1(n_169),
.B2(n_167),
.Y(n_194)
);

A2O1A1O1Ixp25_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_151),
.B(n_152),
.C(n_158),
.D(n_157),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_171),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_162),
.A2(n_142),
.B(n_158),
.Y(n_180)
);

OA21x2_ASAP7_75t_L g184 ( 
.A1(n_162),
.A2(n_150),
.B(n_154),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_140),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_187),
.Y(n_190)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_185),
.Y(n_189)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_179),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_193),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_163),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_195),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_161),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_197),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_172),
.B(n_7),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_200),
.B(n_202),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_184),
.C(n_180),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_204),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_201),
.A2(n_188),
.B1(n_194),
.B2(n_181),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_198),
.C(n_203),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_205),
.A2(n_199),
.B(n_178),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_210),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_206),
.A2(n_198),
.B1(n_192),
.B2(n_183),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_193),
.C(n_207),
.Y(n_212)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_63),
.A3(n_112),
.B1(n_8),
.B2(n_9),
.C1(n_11),
.C2(n_1),
.Y(n_213)
);

AOI31xp67_ASAP7_75t_L g214 ( 
.A1(n_213),
.A2(n_7),
.A3(n_11),
.B(n_12),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_211),
.Y(n_215)
);


endmodule