module fake_jpeg_21053_n_324 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_33),
.B1(n_19),
.B2(n_27),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_28),
.B1(n_25),
.B2(n_32),
.Y(n_60)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

AOI22x1_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_28),
.B1(n_37),
.B2(n_43),
.Y(n_48)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_32),
.B1(n_36),
.B2(n_35),
.Y(n_74)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_33),
.B1(n_30),
.B2(n_27),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_37),
.B1(n_36),
.B2(n_44),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_19),
.B1(n_13),
.B2(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_60),
.B1(n_37),
.B2(n_25),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_58),
.Y(n_77)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_59),
.Y(n_80)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

OR2x4_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_39),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_63),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_54),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_69),
.B1(n_78),
.B2(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_82),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_25),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_72),
.B(n_81),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVxp33_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_38),
.B1(n_44),
.B2(n_41),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_32),
.B1(n_35),
.B2(n_19),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_45),
.B1(n_49),
.B2(n_35),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_84),
.A2(n_92),
.B1(n_74),
.B2(n_70),
.Y(n_115)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_103),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_70),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_35),
.B1(n_38),
.B2(n_29),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_13),
.B1(n_19),
.B2(n_38),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_96),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_100),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_40),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_102),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_81),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_26),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_72),
.C(n_81),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_110),
.C(n_119),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_72),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_121),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_82),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_99),
.B(n_100),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_112),
.A2(n_116),
.B(n_129),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_115),
.B1(n_128),
.B2(n_66),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_67),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_89),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_128),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_64),
.C(n_80),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_64),
.C(n_80),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_130),
.C(n_31),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_74),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_74),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_74),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_75),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_74),
.Y(n_127)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_66),
.B1(n_65),
.B2(n_70),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_97),
.B(n_86),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_103),
.B(n_78),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_71),
.C(n_29),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_136),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_116),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_137),
.B(n_155),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_103),
.B1(n_101),
.B2(n_38),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_138),
.B(n_146),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_13),
.B1(n_101),
.B2(n_11),
.Y(n_139)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_61),
.B1(n_56),
.B2(n_58),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_147),
.B1(n_150),
.B2(n_118),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_105),
.B(n_22),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_142),
.B(n_22),
.Y(n_176)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_41),
.B1(n_52),
.B2(n_44),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_121),
.B1(n_127),
.B2(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_129),
.A2(n_104),
.B1(n_109),
.B2(n_119),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_13),
.C(n_20),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_152),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_107),
.B(n_123),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_9),
.B(n_8),
.Y(n_188)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_163),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_8),
.B(n_10),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_157),
.A2(n_161),
.B(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_159),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_105),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_55),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_118),
.A2(n_111),
.B1(n_108),
.B2(n_106),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_162),
.A2(n_22),
.B1(n_17),
.B2(n_14),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_34),
.C(n_26),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_47),
.C(n_46),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_118),
.B(n_9),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_14),
.B(n_12),
.Y(n_183)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_167),
.A2(n_171),
.B1(n_177),
.B2(n_180),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_170),
.C(n_187),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_150),
.B1(n_145),
.B2(n_166),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_176),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_154),
.A2(n_11),
.B1(n_12),
.B2(n_17),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_178),
.A2(n_183),
.B(n_12),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_20),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_188),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_46),
.B1(n_47),
.B2(n_26),
.Y(n_180)
);

BUFx24_ASAP7_75t_SL g185 ( 
.A(n_151),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_165),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_132),
.A2(n_14),
.B(n_17),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_186),
.A2(n_190),
.B1(n_196),
.B2(n_157),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_34),
.C(n_31),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_31),
.B1(n_1),
.B2(n_2),
.Y(n_190)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_156),
.B(n_20),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_140),
.C(n_148),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_144),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_199),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_211),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_144),
.B1(n_135),
.B2(n_164),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_210),
.B1(n_212),
.B2(n_216),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_141),
.Y(n_203)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_141),
.Y(n_204)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_147),
.Y(n_206)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_208),
.Y(n_234)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_195),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_138),
.Y(n_213)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_168),
.A2(n_148),
.B(n_195),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_218),
.A2(n_55),
.B(n_34),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_178),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_174),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_136),
.B1(n_146),
.B2(n_133),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_182),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_228),
.Y(n_260)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_226),
.B(n_238),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_215),
.B(n_171),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_170),
.C(n_187),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_233),
.C(n_213),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_209),
.A2(n_167),
.B1(n_188),
.B2(n_194),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_232),
.A2(n_217),
.B1(n_210),
.B2(n_213),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_179),
.C(n_169),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_192),
.C(n_177),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_183),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_239),
.B(n_243),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_206),
.Y(n_240)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_241),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_20),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_202),
.B(n_18),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_217),
.C(n_214),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_250),
.C(n_261),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_246),
.A2(n_262),
.B1(n_237),
.B2(n_227),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_259),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_221),
.C(n_208),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_252),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_223),
.B(n_199),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_253),
.B(n_258),
.Y(n_266)
);

FAx1_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_239),
.CI(n_243),
.CON(n_254),
.SN(n_254)
);

XNOR2x1_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_23),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_207),
.Y(n_257)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_34),
.C(n_23),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_34),
.C(n_23),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_21),
.C(n_15),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_226),
.A2(n_6),
.B1(n_7),
.B2(n_2),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_257),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_245),
.C(n_251),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_15),
.C(n_1),
.Y(n_285)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_224),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_274),
.Y(n_283)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

OAI321xp33_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_230),
.A3(n_235),
.B1(n_222),
.B2(n_244),
.C(n_241),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_248),
.A2(n_6),
.B1(n_7),
.B2(n_2),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_276),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_254),
.A2(n_23),
.B1(n_16),
.B2(n_21),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_277),
.B(n_0),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_256),
.C(n_260),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_279),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_254),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_256),
.C(n_21),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_282),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_15),
.C(n_1),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_285),
.B(n_0),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_15),
.C(n_1),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_289),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_0),
.C(n_2),
.Y(n_289)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_269),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_299),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_290),
.A2(n_264),
.B1(n_271),
.B2(n_266),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_288),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_294),
.B(n_301),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_285),
.A2(n_0),
.B(n_3),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_4),
.B(n_5),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_3),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_3),
.Y(n_299)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_287),
.A2(n_3),
.B(n_4),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_287),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_3),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_305),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_295),
.B(n_280),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_310),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_4),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_303),
.B(n_4),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_296),
.B(n_302),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_298),
.B(n_300),
.Y(n_314)
);

AOI21x1_ASAP7_75t_SL g318 ( 
.A1(n_314),
.A2(n_306),
.B(n_312),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_315),
.B(n_307),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_318),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_316),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_313),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_322),
.A2(n_306),
.B(n_5),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_323),
.B(n_5),
.Y(n_324)
);


endmodule