module fake_netlist_5_205_n_1834 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1834);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1834;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_604;
wire n_314;
wire n_433;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_111),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_77),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_125),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_168),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_2),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_34),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_101),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_25),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_87),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_95),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_89),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_131),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_102),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_119),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_71),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

BUFx8_ASAP7_75t_SL g193 ( 
.A(n_169),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_59),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_69),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_45),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_74),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_54),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_60),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_34),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_22),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_30),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_29),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_144),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_85),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_127),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_135),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_165),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_8),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_8),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_149),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_109),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_10),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_67),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_160),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_18),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_3),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_72),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_33),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_83),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_4),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_146),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_54),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_46),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_79),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_22),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_33),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_14),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_92),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_116),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_44),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_26),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_90),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_59),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_42),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_132),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_35),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_100),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_81),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_110),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_65),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_42),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_91),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_27),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_21),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_17),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_82),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_18),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_28),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_20),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_157),
.Y(n_252)
);

INVxp67_ASAP7_75t_SL g253 ( 
.A(n_17),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_73),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_128),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_41),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_124),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_63),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_3),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_51),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_88),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_45),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_35),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_103),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_136),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_80),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_108),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_164),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_152),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_64),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_107),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_23),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_58),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_130),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_1),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_99),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_84),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_167),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_40),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_2),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_70),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_53),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_147),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_143),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_155),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_161),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_20),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_43),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_44),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_137),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_38),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_53),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_57),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_76),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_58),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_25),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_37),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_13),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_86),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_121),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_55),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_19),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_162),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_29),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_117),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_66),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_115),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_24),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_10),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_24),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_51),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_48),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_148),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_134),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_141),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_57),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_154),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_61),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_30),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_96),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_41),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_142),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_23),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_120),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_139),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_68),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_113),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_31),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_64),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_5),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_21),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_78),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_26),
.Y(n_333)
);

BUFx10_ASAP7_75t_L g334 ( 
.A(n_1),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_14),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_122),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_163),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_145),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_159),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_11),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g341 ( 
.A(n_36),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_93),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_98),
.Y(n_343)
);

INVxp33_ASAP7_75t_SL g344 ( 
.A(n_200),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_0),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_211),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_186),
.Y(n_347)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_279),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_193),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_171),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_189),
.B(n_0),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_205),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_211),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_211),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_171),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_221),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_211),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_170),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_198),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_211),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_172),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_173),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_180),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_234),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_211),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_182),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_188),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_191),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_308),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_195),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_308),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_206),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_308),
.Y(n_373)
);

INVxp33_ASAP7_75t_SL g374 ( 
.A(n_287),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_210),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_208),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_283),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_189),
.B(n_4),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_308),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_308),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_171),
.B(n_5),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_284),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_326),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_257),
.B(n_6),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_210),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_209),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_328),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_213),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_328),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_270),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_216),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_328),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_328),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_338),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_219),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_178),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_328),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_202),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_223),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_226),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_174),
.B(n_6),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_202),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_323),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_230),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_221),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_270),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_310),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_298),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_298),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_311),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_221),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_310),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_343),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_311),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_333),
.Y(n_417)
);

BUFx6f_ASAP7_75t_SL g418 ( 
.A(n_215),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_184),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_333),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_178),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_184),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_239),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_178),
.B(n_7),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_323),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_190),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_241),
.Y(n_427)
);

INVxp33_ASAP7_75t_L g428 ( 
.A(n_203),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_259),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_252),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_346),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_350),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_407),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_421),
.B(n_255),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_407),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_346),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_407),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_344),
.A2(n_194),
.B1(n_296),
.B2(n_309),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_408),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_408),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_429),
.B(n_313),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_175),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_413),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_353),
.B(n_313),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_413),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_356),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_350),
.B(n_264),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_350),
.B(n_342),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_356),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_353),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_354),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g452 ( 
.A(n_378),
.B(n_321),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_354),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_357),
.B(n_313),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_357),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_355),
.B(n_265),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_360),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_355),
.B(n_266),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_355),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_360),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_365),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_365),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_345),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_369),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_369),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_371),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_356),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_398),
.B(n_267),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_371),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_356),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_373),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_398),
.B(n_274),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_373),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_419),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_379),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_379),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_398),
.B(n_278),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_380),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_380),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_429),
.B(n_327),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_384),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_384),
.B(n_388),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_388),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_390),
.B(n_327),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_390),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_358),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_393),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_393),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_394),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_394),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_395),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_395),
.B(n_286),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_399),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_399),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_400),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_400),
.Y(n_496)
);

XOR2x2_ASAP7_75t_SL g497 ( 
.A(n_381),
.B(n_203),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_351),
.B(n_190),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_422),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_404),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_404),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_410),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_386),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_410),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_411),
.Y(n_505)
);

OA21x2_ASAP7_75t_L g506 ( 
.A1(n_411),
.A2(n_217),
.B(n_214),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_412),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_450),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_450),
.Y(n_509)
);

INVxp33_ASAP7_75t_L g510 ( 
.A(n_439),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_450),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_450),
.Y(n_512)
);

OR2x6_ASAP7_75t_L g513 ( 
.A(n_498),
.B(n_424),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_361),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_452),
.A2(n_403),
.B1(n_409),
.B2(n_359),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_506),
.Y(n_516)
);

CKINVDCx6p67_ASAP7_75t_R g517 ( 
.A(n_439),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_452),
.A2(n_409),
.B1(n_374),
.B2(n_348),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_451),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_449),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_506),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_497),
.B(n_362),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_432),
.A2(n_385),
.B1(n_391),
.B2(n_375),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_506),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_440),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_440),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_463),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_506),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_451),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_459),
.B(n_363),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_449),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_449),
.Y(n_532)
);

NOR2x1p5_ASAP7_75t_L g533 ( 
.A(n_486),
.B(n_349),
.Y(n_533)
);

AND2x6_ASAP7_75t_L g534 ( 
.A(n_484),
.B(n_175),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_506),
.Y(n_535)
);

OR2x6_ASAP7_75t_L g536 ( 
.A(n_447),
.B(n_448),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_506),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_459),
.B(n_432),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_434),
.B(n_366),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_432),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_486),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_473),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_432),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_L g544 ( 
.A1(n_463),
.A2(n_405),
.B1(n_425),
.B2(n_212),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_449),
.Y(n_545)
);

INVxp33_ASAP7_75t_L g546 ( 
.A(n_438),
.Y(n_546)
);

BUFx4f_ASAP7_75t_L g547 ( 
.A(n_444),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_451),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_434),
.B(n_367),
.Y(n_549)
);

INVx5_ASAP7_75t_L g550 ( 
.A(n_442),
.Y(n_550)
);

BUFx6f_ASAP7_75t_SL g551 ( 
.A(n_444),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_451),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_447),
.B(n_368),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_474),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_449),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_449),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_503),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_449),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_461),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_SL g560 ( 
.A(n_448),
.B(n_426),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_444),
.A2(n_414),
.B1(n_345),
.B2(n_259),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_461),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_461),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_461),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_473),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_465),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_459),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_444),
.B(n_327),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_475),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_465),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_475),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_431),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_456),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_449),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_444),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_497),
.B(n_370),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_465),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_497),
.B(n_372),
.Y(n_578)
);

NOR2x1p5_ASAP7_75t_L g579 ( 
.A(n_456),
.B(n_259),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_431),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_503),
.B(n_405),
.Y(n_581)
);

OR2x6_ASAP7_75t_L g582 ( 
.A(n_458),
.B(n_229),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_458),
.B(n_376),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_468),
.B(n_387),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_468),
.B(n_389),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_472),
.B(n_425),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_467),
.Y(n_587)
);

AND2x6_ASAP7_75t_L g588 ( 
.A(n_484),
.B(n_187),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_472),
.B(n_392),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_431),
.Y(n_590)
);

INVx5_ASAP7_75t_L g591 ( 
.A(n_442),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_444),
.A2(n_418),
.B1(n_335),
.B2(n_297),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_474),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_465),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_467),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_454),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_477),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_467),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_474),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_436),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_436),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_492),
.B(n_397),
.Y(n_602)
);

INVxp33_ASAP7_75t_SL g603 ( 
.A(n_438),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_436),
.Y(n_604)
);

BUFx4f_ASAP7_75t_L g605 ( 
.A(n_454),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_467),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_485),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_485),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_453),
.Y(n_609)
);

BUFx4f_ASAP7_75t_L g610 ( 
.A(n_454),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_485),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_492),
.B(n_401),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_485),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_467),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_467),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_487),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_454),
.A2(n_212),
.B1(n_427),
.B2(n_423),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_484),
.B(n_402),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_499),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_454),
.A2(n_418),
.B1(n_297),
.B2(n_217),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_454),
.B(n_406),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_453),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_487),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_487),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_441),
.B(n_430),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_441),
.B(n_418),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_441),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_L g628 ( 
.A(n_442),
.B(n_187),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_499),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_480),
.Y(n_630)
);

CKINVDCx16_ASAP7_75t_R g631 ( 
.A(n_499),
.Y(n_631)
);

OR2x6_ASAP7_75t_L g632 ( 
.A(n_480),
.B(n_238),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_480),
.B(n_412),
.Y(n_633)
);

INVx4_ASAP7_75t_SL g634 ( 
.A(n_442),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_500),
.A2(n_253),
.B1(n_260),
.B2(n_258),
.Y(n_635)
);

INVx6_ASAP7_75t_L g636 ( 
.A(n_467),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_453),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_500),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_455),
.B(n_281),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_455),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_455),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_500),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_457),
.B(n_324),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_442),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_495),
.B(n_215),
.Y(n_645)
);

CKINVDCx6p67_ASAP7_75t_R g646 ( 
.A(n_442),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_487),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_495),
.B(n_215),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_501),
.A2(n_291),
.B1(n_232),
.B2(n_235),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_493),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_457),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_501),
.B(n_416),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_457),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_493),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_495),
.B(n_215),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_501),
.B(n_418),
.Y(n_656)
);

OAI22xp33_ASAP7_75t_L g657 ( 
.A1(n_505),
.A2(n_428),
.B1(n_340),
.B2(n_176),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_482),
.A2(n_272),
.B1(n_218),
.B2(n_220),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_L g659 ( 
.A1(n_513),
.A2(n_271),
.B1(n_174),
.B2(n_277),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_528),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_528),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_543),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_528),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_513),
.A2(n_597),
.B1(n_573),
.B2(n_588),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_575),
.Y(n_665)
);

BUFx12f_ASAP7_75t_SL g666 ( 
.A(n_582),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_528),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_528),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_573),
.B(n_460),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_543),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_575),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_514),
.B(n_347),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_539),
.B(n_352),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_525),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_597),
.B(n_460),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_625),
.B(n_627),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_549),
.B(n_364),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_627),
.B(n_377),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_630),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_612),
.B(n_462),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_553),
.B(n_382),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_572),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_583),
.B(n_383),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_630),
.B(n_396),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_589),
.B(n_462),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_567),
.B(n_462),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_572),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_567),
.B(n_464),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_638),
.B(n_464),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_638),
.B(n_464),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_510),
.B(n_415),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_580),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_618),
.B(n_303),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_557),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_642),
.B(n_466),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_642),
.B(n_466),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_602),
.B(n_177),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_584),
.B(n_466),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_585),
.B(n_469),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_580),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_536),
.B(n_469),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_536),
.B(n_478),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_590),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_586),
.B(n_307),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_536),
.B(n_478),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_586),
.B(n_315),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_526),
.B(n_181),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_513),
.A2(n_254),
.B1(n_276),
.B2(n_317),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_536),
.B(n_478),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_590),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_617),
.B(n_320),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_540),
.B(n_481),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_522),
.B(n_197),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_540),
.B(n_481),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_516),
.B(n_481),
.Y(n_715)
);

NAND2x1p5_ASAP7_75t_L g716 ( 
.A(n_547),
.B(n_179),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_576),
.B(n_199),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_521),
.B(n_483),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_600),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_538),
.A2(n_482),
.B(n_446),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_600),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_527),
.B(n_322),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_578),
.B(n_201),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_601),
.Y(n_724)
);

A2O1A1Ixp33_ASAP7_75t_L g725 ( 
.A1(n_521),
.A2(n_254),
.B(n_276),
.C(n_317),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_513),
.A2(n_560),
.B1(n_579),
.B2(n_582),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_524),
.B(n_483),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_527),
.B(n_204),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_601),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_581),
.B(n_222),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_604),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_604),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_609),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_609),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_622),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_581),
.B(n_214),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_547),
.A2(n_446),
.B(n_443),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_544),
.B(n_325),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_524),
.B(n_488),
.Y(n_739)
);

A2O1A1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_535),
.A2(n_314),
.B(n_237),
.C(n_207),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_622),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_535),
.B(n_488),
.Y(n_742)
);

BUFx2_ASAP7_75t_SL g743 ( 
.A(n_551),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_592),
.B(n_336),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_637),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_537),
.B(n_488),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_537),
.B(n_489),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_530),
.B(n_224),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_620),
.B(n_337),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_579),
.Y(n_750)
);

INVx8_ASAP7_75t_L g751 ( 
.A(n_551),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_542),
.B(n_489),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_637),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_542),
.B(n_489),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_621),
.B(n_306),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_565),
.B(n_490),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_640),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_640),
.Y(n_758)
);

AO22x2_ASAP7_75t_L g759 ( 
.A1(n_568),
.A2(n_299),
.B1(n_183),
.B2(n_185),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_565),
.B(n_490),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_641),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_596),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_569),
.B(n_490),
.Y(n_763)
);

NOR3xp33_ASAP7_75t_L g764 ( 
.A(n_631),
.B(n_227),
.C(n_225),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_641),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_569),
.B(n_491),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_541),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_571),
.B(n_491),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_651),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_633),
.B(n_507),
.Y(n_770)
);

NAND2xp33_ASAP7_75t_L g771 ( 
.A(n_534),
.B(n_442),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_582),
.B(n_228),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_651),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_571),
.B(n_491),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_626),
.B(n_476),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_653),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_653),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_568),
.B(n_476),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_582),
.B(n_233),
.Y(n_779)
);

NAND2x1_ASAP7_75t_L g780 ( 
.A(n_636),
.B(n_555),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_517),
.B(n_546),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_633),
.B(n_505),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_561),
.B(n_306),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_517),
.B(n_236),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_649),
.B(n_306),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_652),
.B(n_507),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_652),
.B(n_507),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_656),
.B(n_476),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_508),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_639),
.B(n_479),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_508),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_509),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_632),
.B(n_505),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_649),
.B(n_306),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_509),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_643),
.B(n_479),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_534),
.B(n_479),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_534),
.B(n_479),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_599),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_632),
.B(n_243),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_632),
.B(n_245),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_511),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_632),
.B(n_496),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_534),
.B(n_479),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_603),
.B(n_246),
.Y(n_805)
);

BUFx6f_ASAP7_75t_SL g806 ( 
.A(n_534),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_511),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_523),
.B(n_496),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_657),
.B(n_179),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_512),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_L g811 ( 
.A(n_534),
.B(n_442),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_547),
.B(n_183),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_605),
.B(n_185),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_603),
.B(n_249),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_541),
.B(n_250),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_534),
.B(n_446),
.Y(n_816)
);

INVxp67_ASAP7_75t_SL g817 ( 
.A(n_558),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_605),
.B(n_192),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_512),
.Y(n_819)
);

NAND2x1_ASAP7_75t_L g820 ( 
.A(n_636),
.B(n_442),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_596),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_554),
.B(n_256),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_519),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_588),
.B(n_446),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_588),
.A2(n_192),
.B1(n_196),
.B2(n_207),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_605),
.Y(n_826)
);

AOI21x1_ASAP7_75t_L g827 ( 
.A1(n_715),
.A2(n_648),
.B(n_645),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_680),
.B(n_588),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_780),
.A2(n_610),
.B(n_574),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_780),
.A2(n_610),
.B(n_574),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_685),
.B(n_588),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_817),
.A2(n_610),
.B(n_574),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_698),
.B(n_588),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_720),
.A2(n_588),
.B(n_531),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_778),
.A2(n_615),
.B(n_555),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_692),
.Y(n_836)
);

INVx1_ASAP7_75t_SL g837 ( 
.A(n_674),
.Y(n_837)
);

BUFx8_ASAP7_75t_L g838 ( 
.A(n_736),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_682),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_699),
.B(n_515),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_692),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_679),
.Y(n_842)
);

AOI21xp33_ASAP7_75t_L g843 ( 
.A1(n_713),
.A2(n_518),
.B(n_593),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_679),
.B(n_533),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_697),
.B(n_520),
.Y(n_845)
);

O2A1O1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_659),
.A2(n_658),
.B(n_655),
.C(n_628),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_700),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_751),
.Y(n_848)
);

CKINVDCx10_ASAP7_75t_R g849 ( 
.A(n_767),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_682),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_718),
.A2(n_531),
.B(n_520),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_786),
.B(n_787),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_717),
.A2(n_551),
.B1(n_596),
.B2(n_533),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_786),
.B(n_531),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_787),
.B(n_532),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_700),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_816),
.A2(n_558),
.B(n_545),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_727),
.A2(n_545),
.B(n_532),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_770),
.B(n_532),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_824),
.A2(n_558),
.B(n_556),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_728),
.B(n_619),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_770),
.B(n_545),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_790),
.A2(n_558),
.B(n_556),
.Y(n_863)
);

AO21x1_ASAP7_75t_L g864 ( 
.A1(n_716),
.A2(n_723),
.B(n_809),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_751),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_751),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_796),
.A2(n_558),
.B(n_556),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_662),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_805),
.B(n_814),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_673),
.B(n_599),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_SL g871 ( 
.A1(n_740),
.A2(n_294),
.B(n_290),
.C(n_299),
.Y(n_871)
);

OAI321xp33_ASAP7_75t_L g872 ( 
.A1(n_785),
.A2(n_635),
.A3(n_247),
.B1(n_251),
.B2(n_301),
.C(n_304),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_703),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_662),
.B(n_670),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_762),
.A2(n_595),
.B(n_587),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_762),
.A2(n_821),
.B(n_742),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_782),
.B(n_587),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_782),
.B(n_587),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_676),
.A2(n_294),
.B(n_339),
.C(n_332),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_739),
.A2(n_598),
.B(n_595),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_669),
.B(n_595),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_675),
.B(n_598),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_664),
.A2(n_635),
.B1(n_646),
.B2(n_629),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_762),
.A2(n_606),
.B(n_598),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_748),
.B(n_606),
.Y(n_885)
);

AOI21x1_ASAP7_75t_L g886 ( 
.A1(n_746),
.A2(n_548),
.B(n_529),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_821),
.A2(n_614),
.B(n_606),
.Y(n_887)
);

NOR3xp33_ASAP7_75t_L g888 ( 
.A(n_678),
.B(n_631),
.C(n_629),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_808),
.B(n_614),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_703),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_808),
.B(n_614),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_821),
.A2(n_591),
.B(n_550),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_826),
.B(n_550),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_747),
.A2(n_591),
.B(n_550),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_799),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_701),
.A2(n_552),
.B(n_548),
.Y(n_896)
);

O2A1O1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_794),
.A2(n_285),
.B(n_277),
.C(n_290),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_767),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_751),
.Y(n_899)
);

NAND2xp33_ASAP7_75t_L g900 ( 
.A(n_826),
.B(n_196),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_793),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_687),
.B(n_654),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_710),
.B(n_654),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_737),
.A2(n_591),
.B(n_550),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_797),
.A2(n_591),
.B(n_550),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_710),
.B(n_650),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_677),
.B(n_681),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_719),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_793),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_803),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_719),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_666),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_683),
.B(n_262),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_798),
.A2(n_644),
.B(n_591),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_721),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_702),
.A2(n_559),
.B(n_552),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_729),
.B(n_733),
.Y(n_917)
);

NAND3xp33_ASAP7_75t_L g918 ( 
.A(n_815),
.B(n_275),
.C(n_273),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_705),
.A2(n_650),
.B(n_647),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_735),
.B(n_647),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_804),
.A2(n_644),
.B(n_470),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_735),
.B(n_559),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_753),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_775),
.A2(n_644),
.B(n_470),
.Y(n_924)
);

A2O1A1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_708),
.A2(n_726),
.B(n_757),
.C(n_753),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_826),
.A2(n_644),
.B(n_470),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_826),
.A2(n_644),
.B(n_470),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_826),
.A2(n_470),
.B(n_467),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_812),
.A2(n_470),
.B(n_435),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_757),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_694),
.B(n_280),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_758),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_660),
.B(n_634),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_813),
.A2(n_470),
.B(n_435),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_758),
.B(n_562),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_818),
.A2(n_470),
.B(n_435),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_765),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_765),
.Y(n_938)
);

AOI21x1_ASAP7_75t_L g939 ( 
.A1(n_788),
.A2(n_577),
.B(n_562),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_712),
.A2(n_435),
.B(n_443),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_672),
.B(n_282),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_714),
.A2(n_443),
.B(n_437),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_660),
.A2(n_443),
.B(n_437),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_665),
.A2(n_646),
.B1(n_636),
.B2(n_268),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_661),
.B(n_634),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_709),
.A2(n_563),
.B(n_624),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_773),
.B(n_563),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_661),
.A2(n_445),
.B(n_433),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_663),
.A2(n_332),
.B1(n_314),
.B2(n_305),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_SL g950 ( 
.A(n_691),
.B(n_263),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_776),
.A2(n_777),
.B(n_772),
.C(n_779),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_663),
.A2(n_668),
.B(n_667),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_776),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_721),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_724),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_666),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_724),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_731),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_736),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_777),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_667),
.B(n_564),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_668),
.B(n_564),
.Y(n_962)
);

NOR3xp33_ASAP7_75t_L g963 ( 
.A(n_684),
.B(n_261),
.C(n_269),
.Y(n_963)
);

OAI21x1_ASAP7_75t_L g964 ( 
.A1(n_791),
.A2(n_607),
.B(n_624),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_731),
.B(n_566),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_665),
.B(n_634),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_732),
.A2(n_566),
.B(n_623),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_732),
.A2(n_570),
.B(n_623),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_771),
.A2(n_445),
.B(n_437),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_734),
.B(n_570),
.Y(n_970)
);

INVx4_ASAP7_75t_L g971 ( 
.A(n_670),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_771),
.A2(n_445),
.B(n_437),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_820),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_811),
.A2(n_445),
.B(n_437),
.Y(n_974)
);

CKINVDCx11_ASAP7_75t_R g975 ( 
.A(n_764),
.Y(n_975)
);

AOI21xp33_ASAP7_75t_L g976 ( 
.A1(n_730),
.A2(n_231),
.B(n_339),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_822),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_671),
.B(n_634),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_820),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_734),
.B(n_577),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_811),
.A2(n_688),
.B(n_686),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_800),
.A2(n_247),
.B(n_251),
.C(n_301),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_689),
.A2(n_445),
.B(n_433),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_741),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_671),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_707),
.B(n_288),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_750),
.A2(n_237),
.B(n_240),
.C(n_242),
.Y(n_987)
);

AOI21x1_ASAP7_75t_L g988 ( 
.A1(n_752),
.A2(n_607),
.B(n_616),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_690),
.A2(n_433),
.B(n_446),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_695),
.A2(n_433),
.B(n_616),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_741),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_745),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_745),
.B(n_761),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_750),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_761),
.A2(n_242),
.B(n_231),
.C(n_240),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_769),
.B(n_594),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_781),
.B(n_263),
.Y(n_997)
);

INVxp67_ASAP7_75t_L g998 ( 
.A(n_803),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_759),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_806),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_716),
.A2(n_769),
.B1(n_806),
.B2(n_743),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_696),
.B(n_594),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_716),
.A2(n_433),
.B(n_613),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_693),
.A2(n_636),
.B1(n_244),
.B2(n_305),
.Y(n_1004)
);

AOI21x1_ASAP7_75t_L g1005 ( 
.A1(n_754),
.A2(n_613),
.B(n_611),
.Y(n_1005)
);

AO21x1_ASAP7_75t_L g1006 ( 
.A1(n_711),
.A2(n_244),
.B(n_248),
.Y(n_1006)
);

AOI33xp33_ASAP7_75t_L g1007 ( 
.A1(n_825),
.A2(n_318),
.A3(n_304),
.B1(n_335),
.B2(n_331),
.B3(n_330),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_756),
.B(n_608),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_760),
.A2(n_611),
.B(n_608),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_784),
.B(n_263),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_763),
.B(n_248),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_743),
.Y(n_1012)
);

NOR2xp67_ASAP7_75t_SL g1013 ( 
.A(n_848),
.B(n_783),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_839),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_876),
.A2(n_806),
.B(n_766),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_874),
.B(n_704),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_845),
.A2(n_774),
.B(n_768),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_869),
.B(n_801),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_850),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_973),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_833),
.A2(n_755),
.B(n_819),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_848),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_861),
.B(n_722),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_964),
.A2(n_823),
.B(n_819),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_973),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_869),
.A2(n_738),
.B(n_706),
.C(n_744),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_910),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_907),
.A2(n_749),
.B(n_725),
.C(n_823),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_907),
.B(n_789),
.Y(n_1029)
);

NAND3xp33_ASAP7_75t_SL g1030 ( 
.A(n_913),
.B(n_292),
.C(n_312),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_843),
.A2(n_261),
.B(n_268),
.C(n_300),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_986),
.A2(n_789),
.B(n_792),
.C(n_795),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_832),
.A2(n_795),
.B(n_792),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_841),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_847),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_874),
.B(n_791),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_829),
.A2(n_810),
.B(n_807),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_848),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_868),
.B(n_807),
.Y(n_1039)
);

NOR2x1_ASAP7_75t_L g1040 ( 
.A(n_971),
.B(n_802),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_830),
.A2(n_810),
.B(n_759),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_868),
.B(n_269),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_828),
.A2(n_759),
.B(n_271),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_SL g1044 ( 
.A1(n_913),
.A2(n_285),
.B(n_300),
.C(n_502),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_977),
.B(n_289),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_898),
.Y(n_1046)
);

NAND2xp33_ASAP7_75t_SL g1047 ( 
.A(n_848),
.B(n_316),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_986),
.A2(n_329),
.B(n_316),
.C(n_318),
.Y(n_1048)
);

OAI22x1_ASAP7_75t_L g1049 ( 
.A1(n_870),
.A2(n_293),
.B1(n_295),
.B2(n_302),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_831),
.A2(n_759),
.B(n_493),
.Y(n_1050)
);

CKINVDCx6p67_ASAP7_75t_R g1051 ( 
.A(n_849),
.Y(n_1051)
);

INVx1_ASAP7_75t_SL g1052 ( 
.A(n_837),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_SL g1053 ( 
.A(n_872),
.B(n_319),
.C(n_329),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_885),
.A2(n_493),
.B(n_494),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_976),
.A2(n_330),
.B(n_331),
.C(n_417),
.Y(n_1055)
);

BUFx12f_ASAP7_75t_L g1056 ( 
.A(n_838),
.Y(n_1056)
);

NAND2x1p5_ASAP7_75t_L g1057 ( 
.A(n_865),
.B(n_504),
.Y(n_1057)
);

NOR3xp33_ASAP7_75t_L g1058 ( 
.A(n_870),
.B(n_977),
.C(n_888),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_951),
.A2(n_420),
.B(n_416),
.C(n_417),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_840),
.B(n_504),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_852),
.B(n_341),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_842),
.B(n_504),
.Y(n_1062)
);

NAND3xp33_ASAP7_75t_SL g1063 ( 
.A(n_950),
.B(n_420),
.C(n_502),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_959),
.B(n_504),
.Y(n_1064)
);

NAND2xp33_ASAP7_75t_SL g1065 ( 
.A(n_865),
.B(n_495),
.Y(n_1065)
);

BUFx10_ASAP7_75t_L g1066 ( 
.A(n_941),
.Y(n_1066)
);

AOI33xp33_ASAP7_75t_L g1067 ( 
.A1(n_997),
.A2(n_341),
.A3(n_334),
.B1(n_263),
.B2(n_502),
.B3(n_496),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_842),
.B(n_502),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_R g1069 ( 
.A(n_1012),
.B(n_123),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_998),
.B(n_496),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_951),
.A2(n_494),
.B(n_495),
.C(n_471),
.Y(n_1071)
);

NAND2x1p5_ASAP7_75t_L g1072 ( 
.A(n_865),
.B(n_495),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_941),
.A2(n_846),
.B(n_925),
.C(n_981),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_999),
.A2(n_341),
.B1(n_334),
.B2(n_495),
.Y(n_1074)
);

OA21x2_ASAP7_75t_L g1075 ( 
.A1(n_851),
.A2(n_494),
.B(n_442),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_883),
.B(n_341),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_864),
.A2(n_334),
.B1(n_495),
.B2(n_442),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_925),
.A2(n_471),
.B1(n_118),
.B2(n_166),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_998),
.B(n_471),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_923),
.A2(n_334),
.B1(n_471),
.B2(n_11),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_901),
.B(n_7),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_838),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_901),
.B(n_9),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_834),
.A2(n_471),
.B(n_158),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_917),
.A2(n_910),
.B1(n_953),
.B2(n_930),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_R g1086 ( 
.A(n_956),
.B(n_865),
.Y(n_1086)
);

NOR3xp33_ASAP7_75t_SL g1087 ( 
.A(n_982),
.B(n_918),
.C(n_931),
.Y(n_1087)
);

OR2x2_ASAP7_75t_L g1088 ( 
.A(n_909),
.B(n_9),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_835),
.A2(n_471),
.B(n_153),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_R g1090 ( 
.A(n_866),
.B(n_140),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_909),
.B(n_12),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1010),
.B(n_12),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_982),
.A2(n_13),
.B(n_15),
.C(n_16),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_932),
.B(n_15),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_937),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_985),
.B(n_138),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_938),
.B(n_16),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_960),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_931),
.B(n_19),
.Y(n_1099)
);

AO22x1_ASAP7_75t_L g1100 ( 
.A1(n_888),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_973),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_985),
.B(n_106),
.Y(n_1102)
);

O2A1O1Ixp5_ASAP7_75t_L g1103 ( 
.A1(n_1006),
.A2(n_104),
.B(n_97),
.C(n_94),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_847),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_897),
.A2(n_32),
.B(n_36),
.C(n_37),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_912),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_963),
.A2(n_32),
.B(n_38),
.C(n_39),
.Y(n_1107)
);

INVxp67_ASAP7_75t_L g1108 ( 
.A(n_895),
.Y(n_1108)
);

NOR3xp33_ASAP7_75t_SL g1109 ( 
.A(n_949),
.B(n_39),
.C(n_40),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_L g1110 ( 
.A(n_963),
.B(n_43),
.C(n_46),
.Y(n_1110)
);

OAI22x1_ASAP7_75t_L g1111 ( 
.A1(n_895),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_858),
.A2(n_75),
.B(n_49),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_994),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_908),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_975),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_908),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_844),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_889),
.B(n_47),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_975),
.Y(n_1119)
);

BUFx8_ASAP7_75t_SL g1120 ( 
.A(n_844),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_891),
.B(n_50),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_971),
.B(n_50),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_859),
.B(n_52),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_853),
.A2(n_52),
.B(n_55),
.C(n_56),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_879),
.A2(n_1004),
.B(n_991),
.C(n_992),
.Y(n_1125)
);

BUFx8_ASAP7_75t_L g1126 ( 
.A(n_866),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_987),
.A2(n_56),
.B(n_60),
.C(n_61),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_900),
.A2(n_62),
.B(n_63),
.C(n_1011),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_SL g1129 ( 
.A1(n_880),
.A2(n_62),
.B(n_896),
.C(n_919),
.Y(n_1129)
);

OAI22x1_ASAP7_75t_L g1130 ( 
.A1(n_966),
.A2(n_978),
.B1(n_1000),
.B2(n_933),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_857),
.A2(n_860),
.B(n_854),
.Y(n_1131)
);

AO21x1_ASAP7_75t_L g1132 ( 
.A1(n_1001),
.A2(n_993),
.B(n_978),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_862),
.B(n_877),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_985),
.A2(n_955),
.B1(n_991),
.B2(n_992),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_866),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_952),
.A2(n_878),
.B(n_855),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_SL g1137 ( 
.A1(n_966),
.A2(n_933),
.B(n_945),
.C(n_893),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_955),
.B(n_836),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_856),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_961),
.A2(n_962),
.B(n_882),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_985),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_944),
.A2(n_1000),
.B1(n_911),
.B2(n_915),
.Y(n_1142)
);

INVx1_ASAP7_75t_SL g1143 ( 
.A(n_866),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_873),
.B(n_890),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_899),
.B(n_973),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_881),
.A2(n_863),
.B(n_867),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_954),
.A2(n_958),
.B(n_957),
.C(n_984),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_979),
.A2(n_1008),
.B1(n_935),
.B2(n_920),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_902),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_965),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_970),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_899),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1002),
.A2(n_922),
.B1(n_903),
.B2(n_906),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_899),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_871),
.A2(n_995),
.B(n_947),
.C(n_945),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_893),
.A2(n_887),
.B(n_875),
.Y(n_1156)
);

CKINVDCx14_ASAP7_75t_R g1157 ( 
.A(n_899),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_884),
.A2(n_924),
.B(n_980),
.Y(n_1158)
);

NOR3xp33_ASAP7_75t_L g1159 ( 
.A(n_1007),
.B(n_827),
.C(n_946),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1007),
.B(n_916),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_979),
.B(n_996),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_921),
.A2(n_892),
.B(n_894),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_905),
.A2(n_914),
.B(n_927),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_979),
.B(n_989),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_988),
.Y(n_1165)
);

INVx4_ASAP7_75t_L g1166 ( 
.A(n_979),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_967),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1018),
.B(n_983),
.Y(n_1168)
);

NOR2xp67_ASAP7_75t_SL g1169 ( 
.A(n_1056),
.B(n_969),
.Y(n_1169)
);

NAND3x1_ASAP7_75t_L g1170 ( 
.A(n_1058),
.B(n_972),
.C(n_974),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1014),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1019),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1073),
.A2(n_1009),
.B(n_968),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1026),
.A2(n_1003),
.B(n_990),
.C(n_942),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1030),
.A2(n_928),
.B1(n_926),
.B2(n_934),
.Y(n_1175)
);

OA22x2_ASAP7_75t_L g1176 ( 
.A1(n_1111),
.A2(n_1052),
.B1(n_1049),
.B2(n_1108),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1030),
.A2(n_929),
.B1(n_936),
.B2(n_948),
.Y(n_1177)
);

BUFx2_ASAP7_75t_R g1178 ( 
.A(n_1120),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_1071),
.A2(n_940),
.A3(n_943),
.B(n_904),
.Y(n_1179)
);

BUFx10_ASAP7_75t_L g1180 ( 
.A(n_1083),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1087),
.A2(n_871),
.B(n_1005),
.C(n_886),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_1051),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_1113),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1017),
.A2(n_1015),
.B(n_1146),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_1106),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1058),
.A2(n_1124),
.B(n_1076),
.C(n_1031),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_1046),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1016),
.B(n_1117),
.Y(n_1188)
);

INVx4_ASAP7_75t_L g1189 ( 
.A(n_1022),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1016),
.B(n_1036),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1023),
.A2(n_1099),
.B1(n_1061),
.B2(n_1066),
.Y(n_1191)
);

BUFx2_ASAP7_75t_SL g1192 ( 
.A(n_1152),
.Y(n_1192)
);

AOI221x1_ASAP7_75t_L g1193 ( 
.A1(n_1112),
.A2(n_1078),
.B1(n_1084),
.B2(n_1159),
.C(n_1043),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1131),
.A2(n_1148),
.B(n_1158),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1163),
.A2(n_1156),
.B(n_1033),
.Y(n_1195)
);

NAND3x1_ASAP7_75t_L g1196 ( 
.A(n_1083),
.B(n_1091),
.C(n_1067),
.Y(n_1196)
);

AO31x2_ASAP7_75t_L g1197 ( 
.A1(n_1132),
.A2(n_1059),
.A3(n_1032),
.B(n_1165),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1061),
.B(n_1027),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1095),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1027),
.B(n_1108),
.Y(n_1200)
);

INVx5_ASAP7_75t_L g1201 ( 
.A(n_1022),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1140),
.A2(n_1136),
.B(n_1133),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1060),
.A2(n_1021),
.B(n_1028),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1029),
.B(n_1149),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_SL g1205 ( 
.A1(n_1041),
.A2(n_1155),
.B(n_1093),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1081),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1166),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1118),
.A2(n_1121),
.B(n_1123),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1050),
.A2(n_1087),
.B(n_1160),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1022),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1129),
.A2(n_1153),
.B(n_1161),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1150),
.B(n_1151),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_1086),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1098),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1153),
.A2(n_1167),
.B(n_1037),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1089),
.A2(n_1164),
.B(n_1065),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1139),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1130),
.A2(n_1085),
.A3(n_1125),
.B(n_1048),
.Y(n_1218)
);

AOI21xp33_ASAP7_75t_SL g1219 ( 
.A1(n_1045),
.A2(n_1119),
.B(n_1100),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1070),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_1147),
.A2(n_1142),
.A3(n_1054),
.B(n_1105),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1134),
.A2(n_1107),
.A3(n_1144),
.B(n_1094),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_SL g1223 ( 
.A1(n_1166),
.A2(n_1096),
.B(n_1102),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1064),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1159),
.A2(n_1077),
.B(n_1144),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1092),
.B(n_1091),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1079),
.A2(n_1072),
.B(n_1057),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1066),
.B(n_1036),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1053),
.B(n_1074),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1138),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1062),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1053),
.A2(n_1063),
.B(n_1128),
.C(n_1097),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1086),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1145),
.A2(n_1137),
.B(n_1020),
.Y(n_1234)
);

OA21x2_ASAP7_75t_L g1235 ( 
.A1(n_1077),
.A2(n_1103),
.B(n_1102),
.Y(n_1235)
);

OAI22x1_ASAP7_75t_L g1236 ( 
.A1(n_1110),
.A2(n_1042),
.B1(n_1122),
.B2(n_1088),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1075),
.A2(n_1068),
.B(n_1040),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1115),
.Y(n_1238)
);

INVxp67_ASAP7_75t_L g1239 ( 
.A(n_1042),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1063),
.A2(n_1080),
.B1(n_1074),
.B2(n_1039),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1039),
.B(n_1114),
.Y(n_1241)
);

AO32x2_ASAP7_75t_L g1242 ( 
.A1(n_1109),
.A2(n_1044),
.A3(n_1080),
.B1(n_1127),
.B2(n_1103),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1154),
.B(n_1143),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_SL g1244 ( 
.A1(n_1096),
.A2(n_1044),
.B(n_1055),
.C(n_1141),
.Y(n_1244)
);

AOI221x1_ASAP7_75t_L g1245 ( 
.A1(n_1047),
.A2(n_1109),
.B1(n_1034),
.B2(n_1104),
.C(n_1035),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1013),
.A2(n_1020),
.B(n_1025),
.C(n_1101),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_SL g1247 ( 
.A(n_1082),
.B(n_1126),
.Y(n_1247)
);

AOI221xp5_ASAP7_75t_L g1248 ( 
.A1(n_1069),
.A2(n_1116),
.B1(n_1090),
.B2(n_1157),
.C(n_1101),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1025),
.B(n_1069),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1022),
.B(n_1038),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1126),
.A2(n_1038),
.B(n_1135),
.Y(n_1251)
);

NOR4xp25_ASAP7_75t_L g1252 ( 
.A(n_1038),
.B(n_869),
.C(n_498),
.D(n_907),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1038),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1135),
.A2(n_869),
.B(n_907),
.C(n_1026),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1135),
.Y(n_1255)
);

NAND3xp33_ASAP7_75t_L g1256 ( 
.A(n_1018),
.B(n_869),
.C(n_907),
.Y(n_1256)
);

AOI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1041),
.A2(n_939),
.B(n_1131),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1024),
.A2(n_1162),
.B(n_1163),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1026),
.A2(n_869),
.B(n_907),
.C(n_986),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1014),
.Y(n_1260)
);

AOI221xp5_ASAP7_75t_L g1261 ( 
.A1(n_1018),
.A2(n_869),
.B1(n_843),
.B2(n_907),
.C(n_814),
.Y(n_1261)
);

AOI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1041),
.A2(n_939),
.B(n_1131),
.Y(n_1262)
);

BUFx2_ASAP7_75t_SL g1263 ( 
.A(n_1046),
.Y(n_1263)
);

AO31x2_ASAP7_75t_L g1264 ( 
.A1(n_1071),
.A2(n_1132),
.A3(n_1073),
.B(n_1059),
.Y(n_1264)
);

O2A1O1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1018),
.A2(n_869),
.B(n_907),
.C(n_843),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1073),
.A2(n_826),
.B(n_1017),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1052),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1073),
.A2(n_826),
.B(n_1017),
.Y(n_1268)
);

AOI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1041),
.A2(n_939),
.B(n_1131),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1014),
.Y(n_1270)
);

NOR2x1_ASAP7_75t_L g1271 ( 
.A(n_1029),
.B(n_1166),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1018),
.B(n_869),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1014),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1018),
.B(n_869),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1018),
.B(n_869),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1073),
.A2(n_826),
.B(n_1017),
.Y(n_1276)
);

INVxp67_ASAP7_75t_SL g1277 ( 
.A(n_1027),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1023),
.B(n_861),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1018),
.A2(n_869),
.B1(n_907),
.B2(n_673),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1024),
.A2(n_1162),
.B(n_1163),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1024),
.A2(n_1162),
.B(n_1163),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1073),
.A2(n_869),
.B(n_1018),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1073),
.A2(n_869),
.B(n_1018),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1014),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1018),
.B(n_869),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1024),
.A2(n_1162),
.B(n_1163),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1018),
.B(n_869),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1051),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1018),
.B(n_869),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1018),
.B(n_525),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1024),
.A2(n_1162),
.B(n_1163),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1071),
.A2(n_1132),
.A3(n_1073),
.B(n_1059),
.Y(n_1292)
);

OR2x6_ASAP7_75t_L g1293 ( 
.A(n_1046),
.B(n_899),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1022),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1018),
.A2(n_869),
.B1(n_907),
.B2(n_673),
.Y(n_1295)
);

OA21x2_ASAP7_75t_L g1296 ( 
.A1(n_1071),
.A2(n_1073),
.B(n_1041),
.Y(n_1296)
);

BUFx10_ASAP7_75t_L g1297 ( 
.A(n_1083),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1018),
.B(n_869),
.Y(n_1298)
);

AOI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1041),
.A2(n_939),
.B(n_1131),
.Y(n_1299)
);

NAND3xp33_ASAP7_75t_SL g1300 ( 
.A(n_1018),
.B(n_869),
.C(n_907),
.Y(n_1300)
);

AO32x2_ASAP7_75t_L g1301 ( 
.A1(n_1085),
.A2(n_1078),
.A3(n_949),
.B1(n_1148),
.B2(n_883),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1014),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1071),
.A2(n_1132),
.A3(n_1073),
.B(n_1059),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1016),
.B(n_874),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1024),
.A2(n_1162),
.B(n_1163),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1024),
.A2(n_1162),
.B(n_1163),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1022),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_SL g1308 ( 
.A(n_1051),
.B(n_767),
.Y(n_1308)
);

CKINVDCx11_ASAP7_75t_R g1309 ( 
.A(n_1051),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1018),
.B(n_869),
.Y(n_1310)
);

BUFx12f_ASAP7_75t_L g1311 ( 
.A(n_1056),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_1051),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1024),
.A2(n_1162),
.B(n_1163),
.Y(n_1313)
);

AO31x2_ASAP7_75t_L g1314 ( 
.A1(n_1071),
.A2(n_1132),
.A3(n_1073),
.B(n_1059),
.Y(n_1314)
);

OAI22x1_ASAP7_75t_L g1315 ( 
.A1(n_1018),
.A2(n_869),
.B1(n_907),
.B2(n_870),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1024),
.A2(n_1162),
.B(n_1163),
.Y(n_1316)
);

AO32x2_ASAP7_75t_L g1317 ( 
.A1(n_1085),
.A2(n_1078),
.A3(n_949),
.B1(n_1148),
.B2(n_883),
.Y(n_1317)
);

CKINVDCx11_ASAP7_75t_R g1318 ( 
.A(n_1309),
.Y(n_1318)
);

OAI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1279),
.A2(n_1295),
.B1(n_1256),
.B2(n_1261),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1285),
.A2(n_1289),
.B1(n_1176),
.B2(n_1272),
.Y(n_1320)
);

INVx5_ASAP7_75t_L g1321 ( 
.A(n_1201),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1204),
.A2(n_1275),
.B1(n_1274),
.B2(n_1310),
.Y(n_1322)
);

INVx6_ASAP7_75t_L g1323 ( 
.A(n_1293),
.Y(n_1323)
);

INVx6_ASAP7_75t_L g1324 ( 
.A(n_1185),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1267),
.Y(n_1325)
);

INVx8_ASAP7_75t_L g1326 ( 
.A(n_1293),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1298),
.A2(n_1283),
.B1(n_1282),
.B2(n_1229),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1171),
.Y(n_1328)
);

BUFx10_ASAP7_75t_L g1329 ( 
.A(n_1288),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1300),
.A2(n_1265),
.B(n_1259),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1188),
.Y(n_1331)
);

OAI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1191),
.A2(n_1315),
.B1(n_1290),
.B2(n_1219),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1287),
.A2(n_1236),
.B1(n_1278),
.B2(n_1226),
.Y(n_1333)
);

INVx2_ASAP7_75t_SL g1334 ( 
.A(n_1187),
.Y(n_1334)
);

INVx8_ASAP7_75t_L g1335 ( 
.A(n_1250),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1180),
.A2(n_1297),
.B1(n_1198),
.B2(n_1240),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1180),
.A2(n_1297),
.B1(n_1247),
.B2(n_1233),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1209),
.A2(n_1190),
.B1(n_1188),
.B2(n_1206),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1183),
.Y(n_1339)
);

BUFx12f_ASAP7_75t_L g1340 ( 
.A(n_1311),
.Y(n_1340)
);

INVx6_ASAP7_75t_L g1341 ( 
.A(n_1189),
.Y(n_1341)
);

BUFx10_ASAP7_75t_L g1342 ( 
.A(n_1238),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1190),
.A2(n_1168),
.B1(n_1304),
.B2(n_1208),
.Y(n_1343)
);

BUFx12f_ASAP7_75t_L g1344 ( 
.A(n_1304),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1199),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1225),
.A2(n_1239),
.B1(n_1271),
.B2(n_1205),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1248),
.A2(n_1169),
.B1(n_1224),
.B2(n_1235),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1199),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1308),
.A2(n_1263),
.B1(n_1235),
.B2(n_1228),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1200),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1189),
.Y(n_1351)
);

OAI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1249),
.A2(n_1245),
.B1(n_1212),
.B2(n_1193),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1241),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1231),
.A2(n_1220),
.B1(n_1230),
.B2(n_1217),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1270),
.A2(n_1273),
.B1(n_1243),
.B2(n_1211),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1254),
.A2(n_1196),
.B1(n_1214),
.B2(n_1302),
.Y(n_1356)
);

BUFx4f_ASAP7_75t_SL g1357 ( 
.A(n_1182),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1178),
.Y(n_1358)
);

CKINVDCx11_ASAP7_75t_R g1359 ( 
.A(n_1312),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1214),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1192),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1296),
.A2(n_1277),
.B1(n_1276),
.B2(n_1268),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1260),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1260),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_1255),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1284),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1232),
.A2(n_1302),
.B1(n_1170),
.B2(n_1252),
.Y(n_1367)
);

INVx6_ASAP7_75t_L g1368 ( 
.A(n_1210),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1266),
.A2(n_1296),
.B1(n_1202),
.B2(n_1215),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1234),
.A2(n_1216),
.B1(n_1253),
.B2(n_1203),
.Y(n_1370)
);

NAND2x1p5_ASAP7_75t_L g1371 ( 
.A(n_1251),
.B(n_1207),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1253),
.B(n_1307),
.Y(n_1372)
);

CKINVDCx11_ASAP7_75t_R g1373 ( 
.A(n_1294),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1207),
.B(n_1294),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1175),
.A2(n_1177),
.B1(n_1173),
.B2(n_1307),
.Y(n_1375)
);

CKINVDCx6p67_ASAP7_75t_R g1376 ( 
.A(n_1294),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1194),
.A2(n_1184),
.B1(n_1307),
.B2(n_1237),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1246),
.Y(n_1378)
);

BUFx8_ASAP7_75t_L g1379 ( 
.A(n_1242),
.Y(n_1379)
);

INVx6_ASAP7_75t_L g1380 ( 
.A(n_1223),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1218),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1218),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1227),
.Y(n_1383)
);

OAI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1186),
.A2(n_1242),
.B1(n_1317),
.B2(n_1301),
.Y(n_1384)
);

INVx2_ASAP7_75t_SL g1385 ( 
.A(n_1222),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1222),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1195),
.A2(n_1305),
.B(n_1316),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1181),
.A2(n_1174),
.B(n_1244),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_SL g1389 ( 
.A1(n_1242),
.A2(n_1317),
.B(n_1301),
.Y(n_1389)
);

OAI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1301),
.A2(n_1317),
.B1(n_1257),
.B2(n_1299),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1262),
.A2(n_1269),
.B1(n_1222),
.B2(n_1314),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1264),
.A2(n_1314),
.B1(n_1303),
.B2(n_1292),
.Y(n_1392)
);

CKINVDCx11_ASAP7_75t_R g1393 ( 
.A(n_1221),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1197),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1258),
.A2(n_1281),
.B(n_1280),
.Y(n_1395)
);

AOI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1286),
.A2(n_1313),
.B1(n_1306),
.B2(n_1291),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1221),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1197),
.Y(n_1398)
);

BUFx4f_ASAP7_75t_SL g1399 ( 
.A(n_1221),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1292),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1303),
.A2(n_869),
.B1(n_907),
.B2(n_1261),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1179),
.Y(n_1402)
);

INVx6_ASAP7_75t_L g1403 ( 
.A(n_1179),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1201),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1171),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1279),
.A2(n_869),
.B1(n_1295),
.B2(n_1289),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1261),
.A2(n_869),
.B1(n_907),
.B2(n_913),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1261),
.A2(n_869),
.B1(n_907),
.B2(n_913),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1261),
.A2(n_869),
.B1(n_907),
.B2(n_913),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1185),
.Y(n_1410)
);

INVx3_ASAP7_75t_SL g1411 ( 
.A(n_1213),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_SL g1412 ( 
.A1(n_1285),
.A2(n_869),
.B1(n_907),
.B2(n_950),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1267),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1279),
.A2(n_869),
.B1(n_1295),
.B2(n_1289),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1285),
.A2(n_869),
.B1(n_907),
.B2(n_950),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_SL g1416 ( 
.A1(n_1279),
.A2(n_869),
.B(n_907),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1261),
.A2(n_869),
.B1(n_907),
.B2(n_677),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1279),
.A2(n_869),
.B1(n_1295),
.B2(n_950),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1261),
.A2(n_869),
.B1(n_907),
.B2(n_677),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1261),
.A2(n_869),
.B1(n_907),
.B2(n_913),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1279),
.A2(n_869),
.B1(n_1295),
.B2(n_1289),
.Y(n_1421)
);

INVx6_ASAP7_75t_L g1422 ( 
.A(n_1201),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1279),
.A2(n_869),
.B1(n_1295),
.B2(n_950),
.Y(n_1423)
);

OAI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1279),
.A2(n_869),
.B1(n_1295),
.B2(n_950),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1261),
.A2(n_869),
.B1(n_907),
.B2(n_913),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1285),
.A2(n_869),
.B1(n_907),
.B2(n_950),
.Y(n_1426)
);

AOI21xp33_ASAP7_75t_L g1427 ( 
.A1(n_1265),
.A2(n_869),
.B(n_907),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1204),
.B(n_1282),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1261),
.A2(n_869),
.B1(n_907),
.B2(n_677),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1261),
.A2(n_869),
.B1(n_907),
.B2(n_913),
.Y(n_1430)
);

CKINVDCx11_ASAP7_75t_R g1431 ( 
.A(n_1309),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1279),
.A2(n_869),
.B1(n_1295),
.B2(n_1289),
.Y(n_1432)
);

BUFx10_ASAP7_75t_L g1433 ( 
.A(n_1288),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1278),
.B(n_1226),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1172),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_SL g1436 ( 
.A1(n_1285),
.A2(n_869),
.B1(n_907),
.B2(n_950),
.Y(n_1436)
);

CKINVDCx20_ASAP7_75t_R g1437 ( 
.A(n_1309),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1171),
.Y(n_1438)
);

OAI22x1_ASAP7_75t_SL g1439 ( 
.A1(n_1288),
.A2(n_1119),
.B1(n_1182),
.B2(n_1312),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1204),
.B(n_1282),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1386),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1402),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1350),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1380),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1395),
.A2(n_1387),
.B(n_1377),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1380),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1383),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1350),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1353),
.Y(n_1449)
);

AO31x2_ASAP7_75t_L g1450 ( 
.A1(n_1392),
.A2(n_1398),
.A3(n_1394),
.B(n_1382),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1328),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1434),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1322),
.B(n_1327),
.Y(n_1453)
);

OR2x6_ASAP7_75t_L g1454 ( 
.A(n_1380),
.B(n_1388),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1400),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1383),
.B(n_1367),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1381),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1412),
.A2(n_1426),
.B1(n_1436),
.B2(n_1415),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1407),
.A2(n_1430),
.B1(n_1425),
.B2(n_1409),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1397),
.B(n_1392),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1345),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1417),
.A2(n_1419),
.B(n_1429),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1348),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1406),
.A2(n_1421),
.B(n_1432),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1360),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1403),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1405),
.Y(n_1467)
);

AO21x2_ASAP7_75t_L g1468 ( 
.A1(n_1387),
.A2(n_1395),
.B(n_1388),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1385),
.B(n_1428),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1369),
.A2(n_1396),
.B(n_1370),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1408),
.A2(n_1420),
.B(n_1427),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1438),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1363),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1323),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1364),
.Y(n_1475)
);

INVx8_ASAP7_75t_L g1476 ( 
.A(n_1321),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1366),
.B(n_1393),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1399),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1389),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1389),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1378),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1371),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1325),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1413),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1321),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1379),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1371),
.Y(n_1487)
);

AOI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1406),
.A2(n_1414),
.B1(n_1432),
.B2(n_1421),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1391),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1330),
.B(n_1440),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1322),
.B(n_1319),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1428),
.B(n_1440),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1435),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1330),
.B(n_1372),
.Y(n_1494)
);

AO21x2_ASAP7_75t_L g1495 ( 
.A1(n_1390),
.A2(n_1375),
.B(n_1384),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1333),
.B(n_1346),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1356),
.B(n_1336),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1362),
.Y(n_1498)
);

OA21x2_ASAP7_75t_L g1499 ( 
.A1(n_1427),
.A2(n_1401),
.B(n_1347),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1352),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1355),
.A2(n_1354),
.B(n_1343),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1349),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1323),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1365),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1416),
.B(n_1331),
.Y(n_1505)
);

INVx4_ASAP7_75t_L g1506 ( 
.A(n_1404),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1338),
.A2(n_1351),
.B(n_1416),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1374),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1332),
.Y(n_1509)
);

INVx6_ASAP7_75t_L g1510 ( 
.A(n_1344),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1422),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1422),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1404),
.Y(n_1513)
);

AO21x1_ASAP7_75t_L g1514 ( 
.A1(n_1418),
.A2(n_1424),
.B(n_1423),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1320),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1376),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1326),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1326),
.A2(n_1335),
.B(n_1341),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_1341),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1337),
.B(n_1368),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_SL g1521 ( 
.A(n_1358),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1368),
.B(n_1373),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1334),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1490),
.B(n_1361),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1462),
.A2(n_1339),
.B(n_1410),
.C(n_1437),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1491),
.B(n_1411),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1494),
.B(n_1477),
.Y(n_1527)
);

O2A1O1Ixp33_ASAP7_75t_SL g1528 ( 
.A1(n_1458),
.A2(n_1439),
.B(n_1342),
.C(n_1318),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1494),
.B(n_1342),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1477),
.B(n_1324),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1505),
.B(n_1324),
.Y(n_1531)
);

INVxp67_ASAP7_75t_L g1532 ( 
.A(n_1483),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1482),
.B(n_1329),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1490),
.B(n_1329),
.Y(n_1534)
);

AO32x2_ASAP7_75t_L g1535 ( 
.A1(n_1479),
.A2(n_1480),
.A3(n_1474),
.B1(n_1503),
.B2(n_1460),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1459),
.A2(n_1357),
.B1(n_1340),
.B2(n_1433),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1521),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1452),
.B(n_1433),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1449),
.B(n_1359),
.Y(n_1539)
);

A2O1A1Ixp33_ASAP7_75t_L g1540 ( 
.A1(n_1488),
.A2(n_1431),
.B(n_1471),
.C(n_1453),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1514),
.B(n_1488),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1443),
.B(n_1448),
.Y(n_1542)
);

AOI211xp5_ASAP7_75t_L g1543 ( 
.A1(n_1514),
.A2(n_1464),
.B(n_1515),
.C(n_1509),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1469),
.B(n_1480),
.Y(n_1544)
);

A2O1A1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1515),
.A2(n_1509),
.B(n_1497),
.C(n_1501),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1469),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1464),
.A2(n_1454),
.B(n_1476),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1492),
.B(n_1472),
.Y(n_1548)
);

OR3x1_ASAP7_75t_L g1549 ( 
.A(n_1500),
.B(n_1502),
.C(n_1478),
.Y(n_1549)
);

O2A1O1Ixp33_ASAP7_75t_SL g1550 ( 
.A1(n_1497),
.A2(n_1478),
.B(n_1500),
.C(n_1516),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1482),
.B(n_1487),
.Y(n_1551)
);

AO32x2_ASAP7_75t_L g1552 ( 
.A1(n_1474),
.A2(n_1503),
.A3(n_1460),
.B1(n_1519),
.B2(n_1506),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1492),
.B(n_1472),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1472),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1502),
.B(n_1520),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1451),
.Y(n_1556)
);

OAI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1504),
.A2(n_1499),
.B1(n_1498),
.B2(n_1446),
.C(n_1484),
.Y(n_1557)
);

INVxp33_ASAP7_75t_L g1558 ( 
.A(n_1517),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_1523),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1501),
.A2(n_1507),
.B(n_1499),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1508),
.B(n_1496),
.Y(n_1561)
);

NAND4xp25_ASAP7_75t_L g1562 ( 
.A(n_1523),
.B(n_1496),
.C(n_1498),
.D(n_1473),
.Y(n_1562)
);

A2O1A1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1507),
.A2(n_1486),
.B(n_1456),
.C(n_1446),
.Y(n_1563)
);

A2O1A1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1456),
.A2(n_1470),
.B(n_1489),
.C(n_1476),
.Y(n_1564)
);

OAI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1499),
.A2(n_1512),
.B(n_1511),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1465),
.B(n_1467),
.Y(n_1566)
);

OA21x2_ASAP7_75t_L g1567 ( 
.A1(n_1445),
.A2(n_1441),
.B(n_1457),
.Y(n_1567)
);

A2O1A1Ixp33_ASAP7_75t_L g1568 ( 
.A1(n_1476),
.A2(n_1481),
.B(n_1444),
.C(n_1518),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1475),
.B(n_1493),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1461),
.B(n_1463),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1554),
.Y(n_1571)
);

INVxp67_ASAP7_75t_SL g1572 ( 
.A(n_1567),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1543),
.B(n_1444),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1552),
.B(n_1442),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1554),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1566),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1546),
.B(n_1544),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1537),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1552),
.B(n_1442),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1548),
.B(n_1495),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1567),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1553),
.B(n_1495),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1570),
.B(n_1495),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1552),
.B(n_1455),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1535),
.B(n_1455),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1556),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1565),
.Y(n_1587)
);

OR2x6_ASAP7_75t_SL g1588 ( 
.A(n_1542),
.B(n_1466),
.Y(n_1588)
);

INVxp67_ASAP7_75t_SL g1589 ( 
.A(n_1559),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1541),
.A2(n_1499),
.B1(n_1444),
.B2(n_1510),
.Y(n_1590)
);

INVxp67_ASAP7_75t_SL g1591 ( 
.A(n_1569),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1535),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1541),
.A2(n_1540),
.B1(n_1549),
.B2(n_1525),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1535),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1560),
.B(n_1468),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1551),
.B(n_1447),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1532),
.B(n_1450),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1574),
.B(n_1563),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1574),
.B(n_1568),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1596),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1596),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1583),
.B(n_1563),
.Y(n_1602)
);

NOR2x1_ASAP7_75t_L g1603 ( 
.A(n_1597),
.B(n_1549),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1581),
.Y(n_1604)
);

NAND4xp25_ASAP7_75t_L g1605 ( 
.A(n_1593),
.B(n_1540),
.C(n_1528),
.D(n_1545),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_1588),
.Y(n_1606)
);

NAND4xp25_ASAP7_75t_L g1607 ( 
.A(n_1593),
.B(n_1528),
.C(n_1545),
.D(n_1525),
.Y(n_1607)
);

OAI211xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1590),
.A2(n_1557),
.B(n_1524),
.C(n_1536),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1573),
.B(n_1533),
.Y(n_1609)
);

AOI21xp33_ASAP7_75t_L g1610 ( 
.A1(n_1587),
.A2(n_1558),
.B(n_1526),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1579),
.B(n_1564),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1571),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1579),
.B(n_1564),
.Y(n_1613)
);

NOR3xp33_ASAP7_75t_SL g1614 ( 
.A(n_1580),
.B(n_1537),
.C(n_1526),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1571),
.Y(n_1615)
);

AOI31xp33_ASAP7_75t_L g1616 ( 
.A1(n_1587),
.A2(n_1550),
.A3(n_1529),
.B(n_1534),
.Y(n_1616)
);

INVxp67_ASAP7_75t_L g1617 ( 
.A(n_1588),
.Y(n_1617)
);

INVxp67_ASAP7_75t_SL g1618 ( 
.A(n_1572),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1577),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1591),
.B(n_1580),
.Y(n_1620)
);

AOI31xp33_ASAP7_75t_L g1621 ( 
.A1(n_1595),
.A2(n_1550),
.A3(n_1547),
.B(n_1527),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1575),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1583),
.B(n_1562),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1577),
.B(n_1561),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1588),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1586),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1592),
.B(n_1594),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1584),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1626),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1626),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1625),
.B(n_1584),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1600),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1605),
.B(n_1558),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1625),
.B(n_1585),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1623),
.B(n_1591),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1619),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1627),
.B(n_1582),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1612),
.Y(n_1638)
);

NAND2xp33_ASAP7_75t_R g1639 ( 
.A(n_1614),
.B(n_1533),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1612),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1615),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1627),
.B(n_1620),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1628),
.B(n_1599),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1599),
.B(n_1576),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1615),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1620),
.B(n_1602),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1604),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1599),
.B(n_1576),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1622),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1600),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1623),
.B(n_1589),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1599),
.B(n_1576),
.Y(n_1652)
);

NOR2x1_ASAP7_75t_L g1653 ( 
.A(n_1607),
.B(n_1578),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1604),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1646),
.B(n_1602),
.Y(n_1655)
);

NAND2x1p5_ASAP7_75t_L g1656 ( 
.A(n_1653),
.B(n_1603),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1644),
.B(n_1606),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1641),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1646),
.B(n_1619),
.Y(n_1659)
);

NOR2xp67_ASAP7_75t_L g1660 ( 
.A(n_1632),
.B(n_1606),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1646),
.B(n_1617),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1644),
.B(n_1617),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1651),
.B(n_1598),
.Y(n_1663)
);

OAI21xp33_ASAP7_75t_L g1664 ( 
.A1(n_1653),
.A2(n_1605),
.B(n_1607),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1644),
.B(n_1598),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1641),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1647),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1648),
.B(n_1598),
.Y(n_1668)
);

NAND2x1_ASAP7_75t_L g1669 ( 
.A(n_1648),
.B(n_1599),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1641),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1648),
.B(n_1611),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1647),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1629),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1651),
.B(n_1624),
.Y(n_1674)
);

INVx1_ASAP7_75t_SL g1675 ( 
.A(n_1636),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1629),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1630),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1647),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1652),
.B(n_1611),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1633),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1635),
.B(n_1611),
.Y(n_1681)
);

INVxp67_ASAP7_75t_SL g1682 ( 
.A(n_1647),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1630),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1638),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1654),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1654),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1635),
.B(n_1642),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1654),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1638),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1636),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1640),
.B(n_1613),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1652),
.B(n_1613),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1652),
.B(n_1613),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1640),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1645),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1634),
.B(n_1600),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1634),
.B(n_1601),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1658),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1680),
.B(n_1633),
.Y(n_1699)
);

NAND3xp33_ASAP7_75t_L g1700 ( 
.A(n_1664),
.B(n_1608),
.C(n_1614),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1696),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1656),
.B(n_1634),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1656),
.B(n_1631),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1658),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1675),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1656),
.B(n_1671),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1680),
.B(n_1610),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1664),
.B(n_1610),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1696),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1697),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1666),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1675),
.B(n_1539),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1690),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1655),
.B(n_1642),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1690),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1655),
.B(n_1642),
.Y(n_1716)
);

OR2x6_ASAP7_75t_L g1717 ( 
.A(n_1656),
.B(n_1518),
.Y(n_1717)
);

OAI21xp33_ASAP7_75t_L g1718 ( 
.A1(n_1661),
.A2(n_1621),
.B(n_1608),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1697),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1661),
.B(n_1637),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1663),
.B(n_1681),
.Y(n_1721)
);

OAI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1660),
.A2(n_1621),
.B(n_1663),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1671),
.B(n_1631),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1666),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1670),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1670),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1659),
.B(n_1637),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1695),
.Y(n_1728)
);

NAND4xp75_ASAP7_75t_L g1729 ( 
.A(n_1660),
.B(n_1603),
.C(n_1522),
.D(n_1609),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1659),
.B(n_1637),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1657),
.B(n_1631),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1681),
.B(n_1555),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1657),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1674),
.B(n_1530),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1705),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1715),
.B(n_1674),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1713),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1698),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1708),
.B(n_1662),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1706),
.B(n_1662),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1699),
.Y(n_1741)
);

NAND3xp33_ASAP7_75t_L g1742 ( 
.A(n_1700),
.B(n_1687),
.C(n_1691),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1718),
.A2(n_1639),
.B1(n_1669),
.B2(n_1691),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1722),
.B(n_1687),
.Y(n_1744)
);

NOR3xp33_ASAP7_75t_SL g1745 ( 
.A(n_1707),
.B(n_1639),
.C(n_1516),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1698),
.Y(n_1746)
);

AOI211x1_ASAP7_75t_L g1747 ( 
.A1(n_1702),
.A2(n_1679),
.B(n_1693),
.C(n_1692),
.Y(n_1747)
);

INVxp67_ASAP7_75t_L g1748 ( 
.A(n_1712),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1704),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1734),
.B(n_1665),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1706),
.B(n_1733),
.Y(n_1751)
);

OAI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1721),
.A2(n_1669),
.B1(n_1616),
.B2(n_1668),
.C(n_1665),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1731),
.B(n_1668),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1704),
.Y(n_1754)
);

AOI32xp33_ASAP7_75t_L g1755 ( 
.A1(n_1702),
.A2(n_1679),
.A3(n_1693),
.B1(n_1692),
.B2(n_1643),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1729),
.A2(n_1731),
.B1(n_1703),
.B2(n_1723),
.Y(n_1756)
);

INVxp67_ASAP7_75t_SL g1757 ( 
.A(n_1711),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1711),
.Y(n_1758)
);

O2A1O1Ixp33_ASAP7_75t_L g1759 ( 
.A1(n_1703),
.A2(n_1616),
.B(n_1618),
.C(n_1694),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1724),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1757),
.Y(n_1761)
);

OAI32xp33_ASAP7_75t_L g1762 ( 
.A1(n_1744),
.A2(n_1714),
.A3(n_1716),
.B1(n_1720),
.B2(n_1730),
.Y(n_1762)
);

NOR2x1_ASAP7_75t_L g1763 ( 
.A(n_1735),
.B(n_1729),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1751),
.Y(n_1764)
);

INVx5_ASAP7_75t_L g1765 ( 
.A(n_1740),
.Y(n_1765)
);

OAI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1743),
.A2(n_1731),
.B(n_1720),
.Y(n_1766)
);

O2A1O1Ixp5_ASAP7_75t_L g1767 ( 
.A1(n_1739),
.A2(n_1701),
.B(n_1719),
.C(n_1709),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1748),
.B(n_1723),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1752),
.A2(n_1709),
.B1(n_1719),
.B2(n_1701),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1748),
.B(n_1732),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1757),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1737),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1741),
.B(n_1710),
.Y(n_1773)
);

OAI32xp33_ASAP7_75t_L g1774 ( 
.A1(n_1742),
.A2(n_1714),
.A3(n_1716),
.B1(n_1727),
.B2(n_1730),
.Y(n_1774)
);

NAND3xp33_ASAP7_75t_L g1775 ( 
.A(n_1741),
.B(n_1728),
.C(n_1725),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1738),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1736),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1753),
.B(n_1710),
.Y(n_1778)
);

AOI221xp5_ASAP7_75t_L g1779 ( 
.A1(n_1759),
.A2(n_1726),
.B1(n_1725),
.B2(n_1724),
.C(n_1727),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1746),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1765),
.B(n_1745),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1761),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1765),
.B(n_1745),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1771),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1768),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1764),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1763),
.A2(n_1756),
.B1(n_1777),
.B2(n_1779),
.Y(n_1787)
);

CKINVDCx14_ASAP7_75t_R g1788 ( 
.A(n_1765),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1778),
.B(n_1750),
.Y(n_1789)
);

AOI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1762),
.A2(n_1774),
.B1(n_1772),
.B2(n_1775),
.C(n_1773),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1776),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1780),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1781),
.A2(n_1766),
.B(n_1775),
.Y(n_1793)
);

NAND3xp33_ASAP7_75t_L g1794 ( 
.A(n_1790),
.B(n_1767),
.C(n_1769),
.Y(n_1794)
);

INVx1_ASAP7_75t_SL g1795 ( 
.A(n_1783),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1786),
.B(n_1789),
.Y(n_1796)
);

NOR2x1_ASAP7_75t_L g1797 ( 
.A(n_1782),
.B(n_1749),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1790),
.B(n_1755),
.Y(n_1798)
);

NAND4xp25_ASAP7_75t_L g1799 ( 
.A(n_1787),
.B(n_1770),
.C(n_1747),
.D(n_1758),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1788),
.B(n_1754),
.Y(n_1800)
);

NAND4xp75_ASAP7_75t_L g1801 ( 
.A(n_1785),
.B(n_1760),
.C(n_1522),
.D(n_1695),
.Y(n_1801)
);

OAI21xp33_ASAP7_75t_SL g1802 ( 
.A1(n_1784),
.A2(n_1717),
.B(n_1682),
.Y(n_1802)
);

NAND3xp33_ASAP7_75t_L g1803 ( 
.A(n_1794),
.B(n_1792),
.C(n_1791),
.Y(n_1803)
);

OAI221xp5_ASAP7_75t_SL g1804 ( 
.A1(n_1793),
.A2(n_1717),
.B1(n_1682),
.B2(n_1618),
.C(n_1678),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_R g1805 ( 
.A(n_1796),
.B(n_1510),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1798),
.A2(n_1717),
.B(n_1676),
.Y(n_1806)
);

NAND3xp33_ASAP7_75t_L g1807 ( 
.A(n_1799),
.B(n_1717),
.C(n_1672),
.Y(n_1807)
);

NOR2x1_ASAP7_75t_L g1808 ( 
.A(n_1803),
.B(n_1797),
.Y(n_1808)
);

A2O1A1Ixp33_ASAP7_75t_L g1809 ( 
.A1(n_1807),
.A2(n_1806),
.B(n_1795),
.C(n_1804),
.Y(n_1809)
);

NAND3xp33_ASAP7_75t_SL g1810 ( 
.A(n_1805),
.B(n_1800),
.C(n_1801),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1807),
.A2(n_1802),
.B1(n_1694),
.B2(n_1689),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1806),
.B(n_1673),
.Y(n_1812)
);

XNOR2xp5_ASAP7_75t_L g1813 ( 
.A(n_1807),
.B(n_1538),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1808),
.Y(n_1814)
);

NOR2x1_ASAP7_75t_L g1815 ( 
.A(n_1810),
.B(n_1673),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1809),
.B(n_1632),
.Y(n_1816)
);

NOR2x1p5_ASAP7_75t_L g1817 ( 
.A(n_1812),
.B(n_1676),
.Y(n_1817)
);

OAI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1811),
.A2(n_1632),
.B1(n_1650),
.B2(n_1689),
.Y(n_1818)
);

OAI211xp5_ASAP7_75t_L g1819 ( 
.A1(n_1814),
.A2(n_1813),
.B(n_1688),
.C(n_1686),
.Y(n_1819)
);

NOR3xp33_ASAP7_75t_L g1820 ( 
.A(n_1815),
.B(n_1531),
.C(n_1667),
.Y(n_1820)
);

NAND4xp75_ASAP7_75t_L g1821 ( 
.A(n_1816),
.B(n_1683),
.C(n_1684),
.D(n_1677),
.Y(n_1821)
);

OAI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1819),
.A2(n_1818),
.B(n_1817),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1822),
.A2(n_1821),
.B1(n_1820),
.B2(n_1683),
.Y(n_1823)
);

OAI22x1_ASAP7_75t_L g1824 ( 
.A1(n_1823),
.A2(n_1677),
.B1(n_1684),
.B2(n_1685),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1823),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1825),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1824),
.A2(n_1688),
.B1(n_1686),
.B2(n_1685),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1826),
.B(n_1667),
.Y(n_1828)
);

AOI22x1_ASAP7_75t_L g1829 ( 
.A1(n_1827),
.A2(n_1688),
.B1(n_1686),
.B2(n_1685),
.Y(n_1829)
);

OAI21xp33_ASAP7_75t_L g1830 ( 
.A1(n_1828),
.A2(n_1672),
.B(n_1667),
.Y(n_1830)
);

AOI21xp33_ASAP7_75t_L g1831 ( 
.A1(n_1830),
.A2(n_1829),
.B(n_1678),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1831),
.Y(n_1832)
);

AOI221xp5_ASAP7_75t_L g1833 ( 
.A1(n_1832),
.A2(n_1678),
.B1(n_1672),
.B2(n_1654),
.C(n_1649),
.Y(n_1833)
);

AOI211xp5_ASAP7_75t_L g1834 ( 
.A1(n_1833),
.A2(n_1519),
.B(n_1485),
.C(n_1513),
.Y(n_1834)
);


endmodule