module fake_jpeg_14640_n_83 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_83);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_83;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx4f_ASAP7_75t_SL g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_22)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_2),
.B1(n_12),
.B2(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_15),
.B(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_14),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_19),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_21),
.B1(n_18),
.B2(n_2),
.Y(n_47)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_17),
.Y(n_40)
);

NOR2xp67_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_19),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_48),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_47),
.B(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_52),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_21),
.B1(n_18),
.B2(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_23),
.Y(n_52)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_43),
.Y(n_64)
);

OA21x2_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_32),
.B(n_27),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_29),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_11),
.C(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_64),
.B1(n_42),
.B2(n_26),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_45),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_59),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_57),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_57),
.B(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_62),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_70),
.C(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_71),
.B(n_61),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_75),
.B1(n_68),
.B2(n_65),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_69),
.C(n_35),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_76),
.B(n_77),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_72),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_35),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

AOI322xp5_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_80),
.A3(n_79),
.B1(n_27),
.B2(n_9),
.C1(n_4),
.C2(n_41),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_34),
.Y(n_83)
);


endmodule