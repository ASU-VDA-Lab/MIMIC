module fake_jpeg_23427_n_49 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_31;
wire n_17;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_1),
.B(n_8),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_19),
.A2(n_14),
.B(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_25),
.B(n_26),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_12),
.A2(n_0),
.B1(n_4),
.B2(n_6),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_6),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_26),
.B(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_31),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_32),
.B1(n_17),
.B2(n_7),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_10),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_20),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_32),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_8),
.B1(n_17),
.B2(n_31),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_34),
.B1(n_28),
.B2(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_29),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_43),
.B(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

BUFx24_ASAP7_75t_SL g48 ( 
.A(n_47),
.Y(n_48)
);

BUFx24_ASAP7_75t_SL g49 ( 
.A(n_48),
.Y(n_49)
);


endmodule