module fake_jpeg_2269_n_214 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_214);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_37),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_20),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_9),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_78),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_56),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_56),
.B(n_52),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_83),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_61),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_56),
.B1(n_73),
.B2(n_64),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_81),
.B1(n_79),
.B2(n_71),
.Y(n_108)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_94),
.Y(n_109)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_65),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_93),
.Y(n_98)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_71),
.B1(n_55),
.B2(n_61),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_97),
.B(n_106),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_87),
.B(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_99),
.B(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_110),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_63),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_105),
.Y(n_131)
);

OAI22x1_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_71),
.B1(n_81),
.B2(n_79),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_108),
.B1(n_96),
.B2(n_109),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_63),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_59),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_91),
.Y(n_110)
);

BUFx16f_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_52),
.B1(n_69),
.B2(n_70),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_23),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_108),
.B1(n_124),
.B2(n_126),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_117),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_129),
.B1(n_1),
.B2(n_3),
.Y(n_143)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_54),
.B(n_60),
.C(n_75),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_123),
.B(n_132),
.Y(n_150)
);

AO22x1_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_54),
.B1(n_67),
.B2(n_64),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_126),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_55),
.B1(n_67),
.B2(n_72),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_57),
.C(n_72),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_24),
.Y(n_136)
);

CKINVDCx12_ASAP7_75t_R g130 ( 
.A(n_100),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_4),
.Y(n_148)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_122),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_146),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_143),
.B1(n_157),
.B2(n_10),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_3),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

BUFx24_ASAP7_75t_SL g149 ( 
.A(n_135),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_129),
.B1(n_120),
.B2(n_8),
.Y(n_158)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_120),
.A2(n_26),
.B1(n_50),
.B2(n_49),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_175),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_125),
.C(n_117),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_167),
.C(n_171),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_163),
.B(n_161),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_117),
.B(n_25),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_174),
.B(n_27),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_138),
.C(n_155),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_51),
.B1(n_48),
.B2(n_46),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_44),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_43),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_141),
.C(n_144),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_9),
.B(n_10),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_160),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_179),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_145),
.C(n_141),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_159),
.C(n_28),
.Y(n_193)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_185),
.Y(n_192)
);

AOI321xp33_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_162),
.A3(n_159),
.B1(n_140),
.B2(n_16),
.C(n_18),
.Y(n_191)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_187),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_167),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_180),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_183),
.A2(n_168),
.B1(n_173),
.B2(n_140),
.Y(n_189)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_196),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_176),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_40),
.C(n_38),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_176),
.C(n_181),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_183),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_192),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_197),
.A2(n_188),
.B1(n_190),
.B2(n_194),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_201),
.C(n_202),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_204),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_195),
.C(n_193),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_205),
.A2(n_200),
.B1(n_199),
.B2(n_201),
.Y(n_206)
);

OAI321xp33_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_207),
.A3(n_203),
.B1(n_30),
.B2(n_31),
.C(n_35),
.Y(n_208)
);

AOI21x1_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_32),
.B(n_206),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_11),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_22),
.Y(n_212)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_18),
.A3(n_19),
.B1(n_20),
.B2(n_21),
.C1(n_22),
.C2(n_199),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_19),
.Y(n_214)
);


endmodule