module fake_jpeg_27457_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_37),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_43),
.B(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_47),
.B(n_48),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_23),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_35),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_20),
.B(n_32),
.C(n_28),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_48),
.B(n_23),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_59),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_64),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_32),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_16),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_26),
.B1(n_37),
.B2(n_19),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_67),
.B1(n_72),
.B2(n_50),
.Y(n_101)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_69),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_42),
.B1(n_37),
.B2(n_33),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_21),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_42),
.B1(n_49),
.B2(n_53),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_33),
.C(n_29),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_79),
.C(n_85),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_86),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_37),
.B1(n_34),
.B2(n_17),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_77),
.A2(n_91),
.B1(n_92),
.B2(n_16),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_24),
.B(n_19),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_24),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_43),
.B(n_29),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_44),
.B(n_33),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_52),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_60),
.A2(n_17),
.B1(n_25),
.B2(n_32),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_28),
.B1(n_25),
.B2(n_17),
.Y(n_92)
);

FAx1_ASAP7_75t_SL g93 ( 
.A(n_50),
.B(n_39),
.CI(n_38),
.CON(n_93),
.SN(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_39),
.B(n_22),
.C(n_21),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_95),
.A2(n_93),
.B(n_65),
.Y(n_134)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_31),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_108),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_76),
.C(n_90),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_95),
.C(n_121),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_120),
.B1(n_122),
.B2(n_19),
.Y(n_129)
);

AO21x1_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_25),
.B(n_28),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_103),
.A2(n_111),
.B(n_21),
.Y(n_148)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_31),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_109),
.B(n_99),
.Y(n_132)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_33),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_121),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_88),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_58),
.B1(n_16),
.B2(n_24),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_118),
.B1(n_116),
.B2(n_102),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_124),
.B(n_126),
.Y(n_181)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_88),
.B1(n_85),
.B2(n_78),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_129),
.B(n_132),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_78),
.B1(n_65),
.B2(n_66),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_139),
.B1(n_145),
.B2(n_125),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_107),
.C(n_52),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_149),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_134),
.A2(n_140),
.B(n_148),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_108),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_136),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_103),
.B(n_61),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_144),
.Y(n_160)
);

AND2x4_ASAP7_75t_SL g140 ( 
.A(n_100),
.B(n_93),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_73),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_141),
.Y(n_166)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

CKINVDCx10_ASAP7_75t_R g173 ( 
.A(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_81),
.Y(n_144)
);

AO22x1_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_68),
.B1(n_64),
.B2(n_87),
.Y(n_145)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_98),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_152),
.Y(n_167)
);

BUFx4f_ASAP7_75t_SL g147 ( 
.A(n_114),
.Y(n_147)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_114),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_70),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_151),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_86),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_111),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_146),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_144),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_170),
.Y(n_195)
);

BUFx24_ASAP7_75t_SL g158 ( 
.A(n_136),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_159),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_14),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_164),
.C(n_183),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_71),
.C(n_45),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_176),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_71),
.B(n_30),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_185),
.B(n_149),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_115),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_178),
.Y(n_209)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_96),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_171),
.B(n_172),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_96),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_30),
.Y(n_175)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_0),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_182),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_30),
.Y(n_180)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_45),
.C(n_68),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_140),
.A2(n_38),
.B(n_35),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_203),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_188),
.A2(n_200),
.B(n_189),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_185),
.A2(n_140),
.B(n_148),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_168),
.B(n_177),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_129),
.B1(n_145),
.B2(n_137),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_190),
.A2(n_206),
.B1(n_176),
.B2(n_182),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_183),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_194),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_128),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_199),
.C(n_202),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_132),
.C(n_128),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_179),
.A2(n_152),
.B(n_1),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_38),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_58),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_58),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_213),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_161),
.A2(n_143),
.B1(n_45),
.B2(n_7),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_7),
.C(n_15),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_208),
.B(n_211),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_212),
.B(n_155),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_143),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_157),
.A2(n_143),
.B1(n_1),
.B2(n_2),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_215),
.B1(n_176),
.B2(n_163),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_184),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_215)
);

NAND3xp33_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_166),
.C(n_160),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_220),
.B(n_231),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_219),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_177),
.Y(n_218)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_238),
.B1(n_215),
.B2(n_200),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_224),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_184),
.B1(n_159),
.B2(n_170),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_225),
.A2(n_235),
.B1(n_236),
.B2(n_198),
.Y(n_246)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_191),
.B(n_197),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_228),
.Y(n_258)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

FAx1_ASAP7_75t_L g231 ( 
.A(n_190),
.B(n_169),
.CI(n_167),
.CON(n_231),
.SN(n_231)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_204),
.B(n_178),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_234),
.A2(n_209),
.B(n_188),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_163),
.B1(n_167),
.B2(n_173),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_239),
.A2(n_254),
.B1(n_238),
.B2(n_237),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_227),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_246),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_198),
.C(n_199),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_247),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_194),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_205),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_256),
.Y(n_273)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_203),
.B1(n_196),
.B2(n_202),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_233),
.C(n_235),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_257),
.C(n_225),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_186),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_173),
.C(n_7),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_255),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_231),
.C(n_224),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_264),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_274),
.Y(n_283)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_272),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_244),
.B(n_242),
.Y(n_266)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_217),
.Y(n_267)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_239),
.A2(n_222),
.B1(n_231),
.B2(n_3),
.Y(n_268)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_8),
.Y(n_269)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

OAI21x1_ASAP7_75t_L g271 ( 
.A1(n_246),
.A2(n_8),
.B(n_13),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_257),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_250),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_251),
.A2(n_8),
.B(n_13),
.Y(n_274)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_285),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_273),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_247),
.C(n_243),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_248),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_286),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_261),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_273),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_290),
.B(n_295),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_270),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_293),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_249),
.B1(n_270),
.B2(n_254),
.Y(n_293)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_296),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_249),
.B1(n_262),
.B2(n_4),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_280),
.B(n_262),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_298),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_5),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_287),
.B(n_279),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_301),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_284),
.B(n_275),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_283),
.B1(n_9),
.B2(n_5),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_293),
.Y(n_307)
);

AOI221xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.C(n_12),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_303),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_304),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_SL g309 ( 
.A1(n_303),
.A2(n_291),
.B(n_290),
.C(n_6),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_309),
.Y(n_314)
);

AOI31xp67_ASAP7_75t_L g311 ( 
.A1(n_305),
.A2(n_9),
.A3(n_12),
.B(n_15),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_299),
.B(n_2),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_312),
.A2(n_313),
.B(n_310),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_314),
.B1(n_308),
.B2(n_306),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_0),
.B(n_312),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_317),
.Y(n_318)
);


endmodule