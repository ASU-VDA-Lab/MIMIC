module fake_jpeg_2234_n_485 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_485);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_485;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx11_ASAP7_75t_SL g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_59),
.B(n_64),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_60),
.B(n_63),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_16),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_65),
.B(n_70),
.Y(n_144)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g179 ( 
.A(n_66),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_34),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_67),
.B(n_107),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_69),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_21),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_28),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_71),
.A2(n_33),
.B1(n_53),
.B2(n_37),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_72),
.B(n_88),
.Y(n_159)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_34),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_73),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_35),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_74),
.Y(n_138)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_76),
.B(n_79),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_35),
.Y(n_77)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_77),
.Y(n_193)
);

BUFx24_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

CKINVDCx6p67_ASAP7_75t_R g197 ( 
.A(n_78),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_25),
.B(n_17),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

BUFx4f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_15),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_84),
.B(n_92),
.Y(n_166)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_85),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_1),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_87),
.A2(n_89),
.B(n_103),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_21),
.Y(n_88)
);

NAND2x1_ASAP7_75t_SL g89 ( 
.A(n_36),
.B(n_1),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_91),
.B(n_98),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_36),
.B(n_7),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_93),
.Y(n_188)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_95),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_97),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_24),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_24),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_99),
.B(n_108),
.Y(n_198)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_47),
.B(n_14),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

BUFx16f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_106),
.Y(n_182)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_54),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_27),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_27),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_27),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_113),
.B(n_120),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_30),
.B(n_7),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_114),
.B(n_118),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_30),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_30),
.Y(n_116)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_32),
.B(n_7),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g119 ( 
.A(n_32),
.Y(n_119)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_42),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_42),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_122),
.B(n_58),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_60),
.B(n_51),
.C(n_52),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_127),
.B(n_131),
.C(n_192),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_81),
.A2(n_51),
.B1(n_56),
.B2(n_33),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_130),
.A2(n_139),
.B(n_153),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_132),
.A2(n_145),
.B1(n_147),
.B2(n_154),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_56),
.B1(n_49),
.B2(n_42),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g268 ( 
.A1(n_134),
.A2(n_135),
.B1(n_149),
.B2(n_158),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_74),
.A2(n_49),
.B1(n_48),
.B2(n_31),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_104),
.A2(n_26),
.B1(n_41),
.B2(n_40),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_118),
.B1(n_71),
.B2(n_100),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_111),
.A2(n_62),
.B1(n_68),
.B2(n_82),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_74),
.A2(n_67),
.B1(n_101),
.B2(n_77),
.Y(n_149)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_87),
.A2(n_103),
.B1(n_80),
.B2(n_57),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_115),
.A2(n_49),
.B1(n_53),
.B2(n_26),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_94),
.A2(n_23),
.B1(n_31),
.B2(n_48),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_155),
.A2(n_156),
.B1(n_167),
.B2(n_169),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_87),
.A2(n_41),
.B1(n_40),
.B2(n_38),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_93),
.A2(n_38),
.B1(n_37),
.B2(n_9),
.Y(n_158)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_161),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_103),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_102),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_85),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_171),
.A2(n_175),
.B1(n_176),
.B2(n_196),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_90),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_83),
.A2(n_12),
.B1(n_14),
.B2(n_96),
.Y(n_176)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_117),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_107),
.A2(n_14),
.B1(n_117),
.B2(n_106),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_183),
.A2(n_195),
.B1(n_201),
.B2(n_162),
.Y(n_240)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_95),
.Y(n_184)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_184),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_186),
.B(n_187),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_83),
.A2(n_73),
.B1(n_66),
.B2(n_112),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_190),
.A2(n_196),
.B1(n_149),
.B2(n_176),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_105),
.A2(n_89),
.B1(n_73),
.B2(n_109),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_95),
.A2(n_96),
.B1(n_105),
.B2(n_78),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_69),
.A2(n_75),
.B1(n_121),
.B2(n_78),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_138),
.Y(n_204)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_204),
.Y(n_271)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_109),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_207),
.B(n_237),
.Y(n_280)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_125),
.Y(n_208)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_208),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_61),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_209),
.B(n_211),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_129),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_97),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_212),
.B(n_220),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_148),
.A2(n_172),
.B(n_170),
.C(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_213),
.B(n_239),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_124),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_214),
.Y(n_277)
);

INVx6_ASAP7_75t_SL g217 ( 
.A(n_197),
.Y(n_217)
);

INVx13_ASAP7_75t_L g276 ( 
.A(n_217),
.Y(n_276)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_218),
.Y(n_297)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_219),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_144),
.B(n_128),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_221),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_222),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_186),
.A2(n_172),
.B1(n_197),
.B2(n_185),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_SL g291 ( 
.A1(n_223),
.A2(n_240),
.B(n_244),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_224),
.B(n_229),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_148),
.A2(n_198),
.B(n_188),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_225),
.A2(n_213),
.B(n_261),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_134),
.A2(n_155),
.B1(n_135),
.B2(n_175),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_226),
.A2(n_242),
.B1(n_253),
.B2(n_216),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_126),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_227),
.B(n_241),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_228),
.A2(n_255),
.B1(n_226),
.B2(n_248),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_142),
.B(n_179),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_126),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_231),
.B(n_234),
.Y(n_296)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

INVx13_ASAP7_75t_L g279 ( 
.A(n_232),
.Y(n_279)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_140),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_233),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_179),
.B(n_163),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_154),
.A2(n_190),
.B1(n_158),
.B2(n_168),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_235),
.A2(n_228),
.B1(n_249),
.B2(n_207),
.Y(n_272)
);

BUFx6f_ASAP7_75t_SL g236 ( 
.A(n_162),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_133),
.B(n_182),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_165),
.Y(n_238)
);

INVx6_ASAP7_75t_L g307 ( 
.A(n_238),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_165),
.B(n_136),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_168),
.A2(n_180),
.B1(n_141),
.B2(n_181),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_243),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_202),
.A2(n_131),
.B1(n_192),
.B2(n_151),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_140),
.A2(n_177),
.B1(n_146),
.B2(n_189),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_245),
.A2(n_267),
.B1(n_246),
.B2(n_217),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_146),
.A2(n_177),
.B1(n_189),
.B2(n_160),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_246),
.A2(n_248),
.B1(n_249),
.B2(n_224),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_137),
.B(n_184),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_247),
.B(n_251),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_150),
.A2(n_160),
.B1(n_123),
.B2(n_161),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_123),
.A2(n_171),
.B1(n_151),
.B2(n_174),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_152),
.Y(n_250)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_250),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_178),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_253),
.B(n_270),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_199),
.B(n_191),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_254),
.B(n_256),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_202),
.A2(n_191),
.B1(n_199),
.B2(n_152),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_202),
.B(n_129),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_194),
.B(n_148),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_266),
.Y(n_304)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_193),
.Y(n_259)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_259),
.Y(n_313)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_197),
.Y(n_260)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_143),
.Y(n_262)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_262),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_126),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_263),
.Y(n_284)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_138),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_264),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_126),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_265),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_129),
.B(n_164),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_266),
.B(n_269),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_154),
.A2(n_132),
.B1(n_108),
.B2(n_91),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_129),
.B(n_164),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_138),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_272),
.A2(n_301),
.B1(n_314),
.B2(n_274),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_241),
.C(n_225),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_274),
.B(n_287),
.C(n_312),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_278),
.A2(n_302),
.B1(n_206),
.B2(n_259),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_285),
.B(n_275),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_216),
.A2(n_240),
.B1(n_215),
.B2(n_257),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_286),
.A2(n_242),
.B1(n_206),
.B2(n_252),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_237),
.B(n_253),
.C(n_218),
.Y(n_287)
);

INVx8_ASAP7_75t_L g290 ( 
.A(n_230),
.Y(n_290)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_290),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_304),
.B(n_280),
.Y(n_344)
);

AND2x6_ASAP7_75t_L g305 ( 
.A(n_214),
.B(n_261),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_268),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_306),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_221),
.B(n_208),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_251),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_231),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_310),
.B(n_318),
.Y(n_329)
);

AND2x2_ASAP7_75t_SL g311 ( 
.A(n_204),
.B(n_270),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_311),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_239),
.A2(n_268),
.B(n_205),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_314),
.A2(n_268),
.B(n_264),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_203),
.B(n_262),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_320),
.B(n_332),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_321),
.B(n_334),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_322),
.A2(n_326),
.B(n_339),
.Y(n_375)
);

OA22x2_ASAP7_75t_L g323 ( 
.A1(n_301),
.A2(n_268),
.B1(n_230),
.B2(n_243),
.Y(n_323)
);

A2O1A1Ixp33_ASAP7_75t_SL g382 ( 
.A1(n_323),
.A2(n_335),
.B(n_337),
.C(n_276),
.Y(n_382)
);

INVxp33_ASAP7_75t_L g373 ( 
.A(n_324),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_294),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_327),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_330),
.A2(n_348),
.B1(n_299),
.B2(n_295),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_331),
.A2(n_354),
.B1(n_299),
.B2(n_303),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_315),
.B(n_219),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_333),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_315),
.B(n_210),
.Y(n_334)
);

A2O1A1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_286),
.A2(n_232),
.B(n_260),
.C(n_236),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_308),
.Y(n_336)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_336),
.Y(n_367)
);

AO22x2_ASAP7_75t_L g337 ( 
.A1(n_278),
.A2(n_252),
.B1(n_250),
.B2(n_227),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_277),
.B(n_210),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_338),
.B(n_343),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_285),
.A2(n_238),
.B(n_233),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_311),
.Y(n_340)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_340),
.Y(n_371)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_271),
.Y(n_341)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_341),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_275),
.A2(n_304),
.B(n_288),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_342),
.A2(n_326),
.B(n_343),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_280),
.B(n_281),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_298),
.Y(n_357)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_317),
.Y(n_345)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_345),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_300),
.Y(n_346)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_346),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_281),
.B(n_287),
.Y(n_347)
);

A2O1A1O1Ixp25_ASAP7_75t_L g369 ( 
.A1(n_347),
.A2(n_349),
.B(n_279),
.C(n_276),
.D(n_313),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_291),
.A2(n_312),
.B1(n_288),
.B2(n_305),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_312),
.B(n_277),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_297),
.Y(n_350)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_350),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_352),
.C(n_353),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_282),
.B(n_288),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_289),
.B(n_311),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_271),
.A2(n_273),
.B1(n_318),
.B2(n_309),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_273),
.Y(n_355)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_355),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_297),
.B(n_298),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_283),
.C(n_316),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_357),
.B(n_354),
.Y(n_411)
);

OAI22xp33_ASAP7_75t_L g358 ( 
.A1(n_330),
.A2(n_284),
.B1(n_309),
.B2(n_292),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_358),
.A2(n_386),
.B1(n_337),
.B2(n_335),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_325),
.A2(n_284),
.B1(n_310),
.B2(n_292),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_360),
.A2(n_376),
.B(n_377),
.Y(n_401)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_341),
.Y(n_364)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_364),
.Y(n_389)
);

NOR4xp25_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_347),
.C(n_328),
.D(n_321),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_369),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_370),
.Y(n_406)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_355),
.Y(n_374)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_374),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_326),
.A2(n_303),
.B(n_279),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_322),
.A2(n_313),
.B(n_283),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_378),
.B(n_352),
.C(n_353),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_339),
.A2(n_276),
.B(n_307),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_381),
.A2(n_375),
.B(n_382),
.Y(n_403)
);

INVx4_ASAP7_75t_SL g407 ( 
.A(n_382),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_337),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_348),
.A2(n_290),
.B1(n_293),
.B2(n_295),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_363),
.B(n_344),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_387),
.B(n_390),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_362),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_362),
.B(n_327),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_391),
.B(n_397),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_376),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_392),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_351),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_402),
.C(n_409),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_377),
.B(n_342),
.Y(n_394)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_394),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_395),
.Y(n_415)
);

OAI21xp33_ASAP7_75t_L g397 ( 
.A1(n_371),
.A2(n_349),
.B(n_346),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_364),
.Y(n_398)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_398),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_399),
.A2(n_403),
.B(n_369),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_333),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_400),
.B(n_408),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_361),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_410),
.Y(n_418)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_380),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_363),
.B(n_329),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_368),
.B(n_356),
.C(n_323),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_365),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_367),
.B(n_323),
.Y(n_412)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_412),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_393),
.B(n_378),
.C(n_357),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_424),
.C(n_427),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_411),
.Y(n_434)
);

XOR2x2_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_399),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_359),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_401),
.A2(n_375),
.B(n_381),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_425),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_401),
.A2(n_360),
.B(n_325),
.Y(n_426)
);

CKINVDCx14_ASAP7_75t_R g445 ( 
.A(n_426),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_370),
.C(n_361),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_406),
.A2(n_383),
.B1(n_358),
.B2(n_386),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_430),
.A2(n_432),
.B1(n_412),
.B2(n_407),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_390),
.B(n_374),
.Y(n_431)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_431),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_395),
.A2(n_373),
.B1(n_382),
.B2(n_323),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_403),
.A2(n_382),
.B(n_373),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_433),
.A2(n_335),
.B(n_396),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_439),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_435),
.A2(n_448),
.B1(n_415),
.B2(n_418),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_425),
.A2(n_388),
.B(n_394),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_437),
.A2(n_442),
.B1(n_444),
.B2(n_421),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_429),
.B(n_400),
.Y(n_438)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_438),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_414),
.B(n_394),
.C(n_387),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_439),
.B(n_419),
.C(n_414),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_420),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_408),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_431),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_443),
.B(n_449),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_422),
.A2(n_407),
.B1(n_382),
.B2(n_391),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_428),
.B(n_410),
.Y(n_446)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_446),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_422),
.A2(n_407),
.B1(n_405),
.B2(n_398),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_458),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_456),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_455),
.A2(n_444),
.B(n_426),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_434),
.B(n_427),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_457),
.B(n_459),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_443),
.A2(n_430),
.B1(n_432),
.B2(n_418),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_436),
.B(n_424),
.C(n_416),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_460),
.B(n_461),
.C(n_437),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_421),
.C(n_423),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_469),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_441),
.C(n_445),
.Y(n_466)
);

CKINVDCx14_ASAP7_75t_R g467 ( 
.A(n_454),
.Y(n_467)
);

INVx11_ASAP7_75t_L g471 ( 
.A(n_467),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_452),
.A2(n_441),
.B(n_447),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_468),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_465),
.B(n_456),
.C(n_457),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_466),
.A2(n_459),
.B1(n_453),
.B2(n_415),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_465),
.B(n_446),
.C(n_451),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_470),
.A2(n_463),
.B1(n_446),
.B2(n_413),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_476),
.B(n_477),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_475),
.B(n_464),
.C(n_462),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_475),
.B(n_462),
.C(n_448),
.Y(n_478)
);

AOI21x1_ASAP7_75t_L g479 ( 
.A1(n_478),
.A2(n_474),
.B(n_473),
.Y(n_479)
);

AOI322xp5_ASAP7_75t_L g482 ( 
.A1(n_479),
.A2(n_472),
.A3(n_440),
.B1(n_417),
.B2(n_389),
.C1(n_319),
.C2(n_379),
.Y(n_482)
);

AOI322xp5_ASAP7_75t_L g481 ( 
.A1(n_480),
.A2(n_471),
.A3(n_433),
.B1(n_449),
.B2(n_417),
.C1(n_396),
.C2(n_389),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_481),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_483),
.A2(n_482),
.B1(n_372),
.B2(n_385),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_484),
.B(n_384),
.Y(n_485)
);


endmodule