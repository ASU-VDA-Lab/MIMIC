module fake_jpeg_21564_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_0),
.C(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_16),
.B(n_24),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_48),
.Y(n_61)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_SL g46 ( 
.A1(n_29),
.A2(n_28),
.B(n_17),
.C(n_18),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_49),
.B1(n_50),
.B2(n_30),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_16),
.B(n_24),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_32),
.A2(n_21),
.B1(n_13),
.B2(n_25),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_21),
.B1(n_17),
.B2(n_13),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_27),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_53),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_27),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_65),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

BUFx2_ASAP7_75t_SL g62 ( 
.A(n_42),
.Y(n_62)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_70),
.Y(n_77)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_25),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_47),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_68),
.C(n_40),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_31),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

CKINVDCx11_ASAP7_75t_R g71 ( 
.A(n_69),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_58),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_76),
.B(n_81),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_41),
.C(n_52),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_58),
.C(n_59),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_51),
.B1(n_46),
.B2(n_53),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_46),
.B(n_53),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_50),
.B(n_1),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_85),
.B(n_18),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_61),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_89),
.C(n_90),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_58),
.B(n_69),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_97),
.B(n_74),
.Y(n_101)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_92),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_64),
.C(n_60),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_80),
.C(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_96),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_20),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_104),
.B1(n_106),
.B2(n_103),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_31),
.C(n_14),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_73),
.B1(n_86),
.B2(n_90),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_78),
.B1(n_77),
.B2(n_83),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_89),
.A2(n_83),
.B1(n_82),
.B2(n_78),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_112),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_91),
.B(n_82),
.C(n_63),
.D(n_28),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_107),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_111),
.C(n_99),
.Y(n_119)
);

AO221x1_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_75),
.B1(n_98),
.B2(n_3),
.C(n_1),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_3),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_116),
.Y(n_121)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_117),
.A2(n_120),
.B(n_19),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_75),
.A3(n_26),
.B1(n_19),
.B2(n_15),
.C1(n_4),
.C2(n_8),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_99),
.C(n_15),
.Y(n_120)
);

AOI221xp5_ASAP7_75t_SL g122 ( 
.A1(n_118),
.A2(n_113),
.B1(n_14),
.B2(n_26),
.C(n_20),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_123),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_115),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_4),
.A3(n_5),
.B1(n_7),
.B2(n_11),
.C1(n_75),
.C2(n_126),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_127),
.C(n_128),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_7),
.Y(n_131)
);


endmodule