module fake_netlist_6_1643_n_191 (n_41, n_52, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_54, n_27, n_3, n_14, n_38, n_0, n_39, n_60, n_59, n_32, n_4, n_36, n_22, n_26, n_55, n_13, n_35, n_11, n_28, n_17, n_23, n_58, n_12, n_20, n_50, n_49, n_7, n_30, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_31, n_25, n_40, n_57, n_53, n_51, n_44, n_56, n_191);

input n_41;
input n_52;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_54;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_39;
input n_60;
input n_59;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_55;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_58;
input n_12;
input n_20;
input n_50;
input n_49;
input n_7;
input n_30;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_31;
input n_25;
input n_40;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_191;

wire n_91;
wire n_119;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_158;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_87;
wire n_189;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_155;
wire n_62;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_140;
wire n_70;
wire n_120;
wire n_67;
wire n_82;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_181;
wire n_76;
wire n_182;
wire n_124;
wire n_126;
wire n_97;
wire n_108;
wire n_94;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_65;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_190;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_171;
wire n_169;

INVxp67_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_13),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_8),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_35),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_14),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_7),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_12),
.Y(n_83)
);

NOR2xp67_ASAP7_75t_L g84 ( 
.A(n_16),
.B(n_50),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_31),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_9),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_22),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_53),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_28),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

BUFx8_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_72),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_65),
.B(n_0),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVxp67_ASAP7_75t_SL g116 ( 
.A(n_110),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_109),
.B(n_69),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_84),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_111),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_61),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_85),
.Y(n_126)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_80),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

AND2x4_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_130),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

AND2x4_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_96),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_91),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_88),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NAND2x1p5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_81),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_83),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

AND2x4_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_123),
.Y(n_145)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_86),
.B1(n_87),
.B2(n_92),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_125),
.C(n_89),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_133),
.Y(n_152)
);

BUFx4f_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

NAND2x2_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_143),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

AND2x4_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_82),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

AO21x2_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_93),
.B(n_94),
.Y(n_162)
);

AOI221xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_127),
.B1(n_5),
.B2(n_6),
.Y(n_164)
);

AOI221xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_144),
.B1(n_153),
.B2(n_147),
.C(n_148),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_154),
.B1(n_146),
.B2(n_157),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_17),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

AOI221xp5_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.C(n_26),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_162),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_169),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_166),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_170),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_172),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_179),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_181),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_59),
.Y(n_184)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_33),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_185),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_34),
.B(n_37),
.C(n_38),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

AOI222xp33_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.C1(n_46),
.C2(n_47),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_57),
.B(n_58),
.Y(n_191)
);


endmodule