module real_jpeg_12152_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_3),
.A2(n_27),
.B1(n_31),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_3),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_3),
.A2(n_41),
.B1(n_50),
.B2(n_52),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_3),
.A2(n_41),
.B1(n_63),
.B2(n_66),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_5),
.A2(n_50),
.B1(n_52),
.B2(n_56),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_5),
.A2(n_56),
.B1(n_63),
.B2(n_66),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_5),
.A2(n_27),
.B1(n_31),
.B2(n_56),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_6),
.A2(n_50),
.B1(n_52),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_6),
.A2(n_63),
.B1(n_66),
.B2(n_71),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_71),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_6),
.A2(n_27),
.B1(n_31),
.B2(n_71),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_8),
.A2(n_63),
.B1(n_66),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_8),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_8),
.A2(n_50),
.B1(n_52),
.B2(n_78),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_8),
.A2(n_37),
.B1(n_38),
.B2(n_78),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_8),
.A2(n_27),
.B1(n_31),
.B2(n_78),
.Y(n_286)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_10),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_10),
.A2(n_31),
.B(n_34),
.C(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_10),
.B(n_39),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_10),
.A2(n_30),
.B1(n_50),
.B2(n_52),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_10),
.A2(n_87),
.B1(n_116),
.B2(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_10),
.B(n_54),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_11),
.A2(n_63),
.B1(n_66),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_11),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_11),
.A2(n_50),
.B1(n_52),
.B2(n_80),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_11),
.A2(n_37),
.B1(n_38),
.B2(n_80),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_11),
.A2(n_27),
.B1(n_31),
.B2(n_80),
.Y(n_296)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_13),
.A2(n_27),
.B1(n_31),
.B2(n_45),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_13),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_13),
.A2(n_45),
.B1(n_63),
.B2(n_66),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_14),
.A2(n_50),
.B1(n_52),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_14),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_68),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_14),
.A2(n_63),
.B1(n_66),
.B2(n_68),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_14),
.A2(n_27),
.B1(n_31),
.B2(n_68),
.Y(n_246)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_315),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_307),
.B(n_314),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_273),
.B(n_304),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_251),
.B(n_272),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_224),
.B(n_250),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_125),
.B(n_203),
.C(n_223),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_98),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_23),
.B(n_98),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_72),
.C(n_85),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_24),
.B(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_42),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_25),
.B(n_43),
.C(n_57),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_39),
.B2(n_40),
.Y(n_25)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_30),
.A2(n_35),
.B(n_37),
.Y(n_82)
);

HAxp5_ASAP7_75t_SL g135 ( 
.A(n_30),
.B(n_38),
.CON(n_135),
.SN(n_135)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_30),
.B(n_61),
.C(n_66),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_30),
.B(n_87),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_30),
.B(n_62),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_32),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_32),
.A2(n_39),
.B1(n_107),
.B2(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_32),
.B(n_269),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_32),
.A2(n_39),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_36),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_36),
.A2(n_286),
.B(n_287),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_38),
.B1(n_48),
.B2(n_49),
.Y(n_53)
);

NOR3xp33_ASAP7_75t_L g136 ( 
.A(n_37),
.B(n_49),
.C(n_50),
.Y(n_136)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_39),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_39),
.B(n_269),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_57),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_54),
.B2(n_55),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_44),
.Y(n_97)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_46),
.A2(n_54),
.B1(n_95),
.B2(n_135),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_46),
.A2(n_111),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_46),
.B(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_46),
.A2(n_54),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_46),
.A2(n_54),
.B(n_111),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_53),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_47),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_47),
.B(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_47),
.A2(n_240),
.B(n_241),
.Y(n_239)
);

OA22x2_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_48),
.A2(n_52),
.B(n_134),
.C(n_136),
.Y(n_133)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_50),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_52),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_52),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_54),
.B(n_111),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_55),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_67),
.B(n_69),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_58),
.B(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_58),
.A2(n_142),
.B1(n_144),
.B2(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_58),
.A2(n_144),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_58),
.A2(n_144),
.B1(n_152),
.B2(n_162),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_58),
.A2(n_144),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_58),
.A2(n_69),
.B(n_212),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_58),
.A2(n_67),
.B(n_144),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_66),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_62),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

CKINVDCx6p67_ASAP7_75t_R g66 ( 
.A(n_63),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_66),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_67),
.B(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_72),
.B(n_85),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_74),
.A2(n_119),
.B(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_74),
.A2(n_75),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_75),
.B(n_138),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_79),
.Y(n_117)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_83),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_91),
.C(n_93),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_86),
.A2(n_91),
.B1(n_92),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_90),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_87),
.A2(n_116),
.B1(n_167),
.B2(n_175),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_87),
.A2(n_116),
.B(n_231),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_88),
.B(n_185),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_93),
.B(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g280 ( 
.A1(n_96),
.A2(n_281),
.B(n_282),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_113),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_99),
.B(n_114),
.C(n_124),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_112),
.Y(n_99)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_103),
.B(n_108),
.C(n_112),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_104),
.A2(n_244),
.B(n_245),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_104),
.A2(n_267),
.B(n_268),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_104),
.A2(n_268),
.B(n_311),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_110),
.B(n_241),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_124),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_115),
.B(n_120),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_116),
.A2(n_169),
.B(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_121),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_122),
.B(n_143),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_198),
.B(n_202),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_153),
.B(n_197),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_148),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_130),
.B(n_148),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_145),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_139),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_132),
.B(n_139),
.C(n_145),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_137),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_138),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B(n_143),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.C(n_151),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_151),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_192),
.B(n_196),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_181),
.B(n_191),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_170),
.B(n_180),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_165),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_165),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_163),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_176),
.B(n_179),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_183),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_187),
.C(n_190),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_189),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_195),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_201),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_222),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_222),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_207),
.C(n_214),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_214),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_213),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_213),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_210),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_217),
.C(n_220),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_218),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_221),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_226),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_249),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_234),
.B1(n_247),
.B2(n_248),
.Y(n_227)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_248),
.C(n_249),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_229),
.A2(n_230),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_232),
.Y(n_263)
);

AOI21xp33_ASAP7_75t_L g289 ( 
.A1(n_230),
.A2(n_263),
.B(n_265),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_239),
.C(n_243),
.Y(n_254)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_243),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_240),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_245),
.B(n_287),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_246),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_271),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_271),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_270),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_253),
.B(n_256),
.C(n_262),
.Y(n_302)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_262),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_260),
.B(n_261),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_257),
.B(n_260),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_259),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_276),
.C(n_289),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g303 ( 
.A(n_261),
.B(n_276),
.CI(n_289),
.CON(n_303),
.SN(n_303)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_301),
.Y(n_273)
);

AOI21xp33_ASAP7_75t_L g304 ( 
.A1(n_274),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_290),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_290),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_285),
.B2(n_288),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_283),
.B2(n_284),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_284),
.C(n_285),
.Y(n_291)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_284),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_294),
.C(n_299),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_285),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_285),
.A2(n_288),
.B1(n_293),
.B2(n_300),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_291),
.C(n_300),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_286),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_297),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_296),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_298),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_303),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_313),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_308),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_318),
.Y(n_320)
);

FAx1_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_310),
.CI(n_312),
.CON(n_308),
.SN(n_308)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_320),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);


endmodule