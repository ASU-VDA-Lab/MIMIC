module fake_jpeg_14502_n_592 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_592);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_592;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_10),
.B(n_5),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx2_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_6),
.B(n_10),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_13),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_60),
.Y(n_212)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_62),
.Y(n_164)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_64),
.Y(n_173)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_65),
.Y(n_172)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_67),
.Y(n_157)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g209 ( 
.A(n_68),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_26),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_69),
.B(n_71),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_70),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_26),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_72),
.Y(n_182)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_74),
.Y(n_205)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_76),
.B(n_78),
.Y(n_147)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_23),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_79),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_80),
.Y(n_218)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_81),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_23),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_82),
.B(n_87),
.Y(n_161)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_84),
.Y(n_168)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_85),
.Y(n_200)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_86),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_17),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_88),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_89),
.Y(n_199)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_91),
.Y(n_206)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_53),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_92),
.Y(n_198)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_94),
.Y(n_201)
);

INVx6_ASAP7_75t_SL g95 ( 
.A(n_53),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_95),
.B(n_98),
.Y(n_162)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_97),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_23),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_99),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_39),
.B(n_0),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_107),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_23),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_101),
.B(n_103),
.Y(n_165)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_19),
.Y(n_102)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_55),
.B(n_0),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_117),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_106),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_39),
.B(n_15),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_19),
.Y(n_108)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_23),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_110),
.B(n_114),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_45),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_45),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_116),
.B(n_118),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_22),
.B(n_1),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_45),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_40),
.Y(n_122)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g171 ( 
.A(n_123),
.Y(n_171)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_47),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_124),
.B(n_38),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_22),
.B(n_1),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_125),
.B(n_52),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_40),
.Y(n_126)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_126),
.Y(n_215)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_27),
.Y(n_127)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_46),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_2),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_67),
.A2(n_28),
.B1(n_27),
.B2(n_53),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_133),
.A2(n_136),
.B1(n_149),
.B2(n_153),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_24),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_135),
.B(n_151),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_72),
.A2(n_90),
.B1(n_62),
.B2(n_64),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_70),
.A2(n_24),
.B1(n_33),
.B2(n_56),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_139),
.A2(n_145),
.B1(n_163),
.B2(n_202),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_88),
.A2(n_28),
.B1(n_42),
.B2(n_51),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_89),
.A2(n_42),
.B1(n_51),
.B2(n_54),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_76),
.B(n_33),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_97),
.A2(n_29),
.B1(n_57),
.B2(n_56),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_128),
.A2(n_28),
.B1(n_42),
.B2(n_54),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_156),
.A2(n_176),
.B1(n_181),
.B2(n_187),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_60),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_158),
.B(n_183),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_111),
.A2(n_29),
.B1(n_57),
.B2(n_52),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_167),
.B(n_9),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g237 ( 
.A(n_174),
.B(n_179),
.C(n_197),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_112),
.A2(n_50),
.B1(n_48),
.B2(n_43),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g178 ( 
.A1(n_127),
.A2(n_50),
.B(n_48),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g276 ( 
.A1(n_178),
.A2(n_133),
.B(n_156),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_59),
.B(n_43),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_80),
.A2(n_38),
.B1(n_37),
.B2(n_30),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_61),
.B(n_37),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_192),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_115),
.A2(n_30),
.B1(n_58),
.B2(n_45),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_74),
.B(n_58),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_106),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_194),
.A2(n_211),
.B1(n_213),
.B2(n_216),
.Y(n_280)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_104),
.Y(n_195)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_79),
.B(n_5),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_196),
.B(n_204),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_65),
.B(n_5),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_123),
.A2(n_45),
.B1(n_7),
.B2(n_8),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_60),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_126),
.A2(n_122),
.B1(n_99),
.B2(n_84),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_113),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_119),
.B(n_7),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_214),
.B(n_212),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_93),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_85),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_217),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_136),
.A2(n_109),
.B1(n_102),
.B2(n_91),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_219),
.A2(n_239),
.B1(n_265),
.B2(n_280),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_167),
.A2(n_91),
.B1(n_68),
.B2(n_13),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_220),
.A2(n_221),
.B(n_243),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_221),
.B(n_276),
.Y(n_326)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_222),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_162),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_223),
.B(n_231),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_134),
.B(n_12),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_224),
.Y(n_347)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_225),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_226),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_230),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_209),
.Y(n_231)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

INVx3_ASAP7_75t_SL g310 ( 
.A(n_232),
.Y(n_310)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_144),
.Y(n_233)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_233),
.Y(n_308)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_130),
.Y(n_234)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_234),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_129),
.B(n_14),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_235),
.B(n_257),
.Y(n_302)
);

INVx11_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_193),
.Y(n_238)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_238),
.Y(n_312)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_154),
.Y(n_240)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_240),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_147),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_242),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_140),
.A2(n_14),
.B(n_216),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_243),
.A2(n_220),
.B(n_221),
.Y(n_338)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_160),
.Y(n_244)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_244),
.Y(n_342)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_142),
.Y(n_245)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_245),
.Y(n_298)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_157),
.Y(n_246)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_246),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_148),
.B(n_188),
.C(n_169),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_247),
.B(n_260),
.C(n_264),
.Y(n_323)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_207),
.Y(n_248)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_165),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_249),
.B(n_272),
.Y(n_296)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_157),
.Y(n_250)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_250),
.Y(n_311)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_164),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_251),
.Y(n_314)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_168),
.Y(n_252)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_252),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_198),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_253),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_173),
.Y(n_254)
);

INVx8_ASAP7_75t_L g339 ( 
.A(n_254),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_173),
.Y(n_255)
);

INVx8_ASAP7_75t_L g349 ( 
.A(n_255),
.Y(n_349)
);

INVx11_ASAP7_75t_L g256 ( 
.A(n_206),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_256),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_166),
.B(n_180),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_155),
.A2(n_210),
.B1(n_218),
.B2(n_215),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_258),
.A2(n_267),
.B1(n_283),
.B2(n_290),
.Y(n_321)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_146),
.Y(n_259)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_259),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_137),
.B(n_161),
.Y(n_260)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_177),
.Y(n_261)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_261),
.Y(n_324)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_146),
.Y(n_262)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_262),
.Y(n_325)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_170),
.Y(n_263)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_263),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_209),
.B(n_175),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_266),
.B(n_273),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_155),
.A2(n_218),
.B1(n_215),
.B2(n_171),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_176),
.B(n_181),
.Y(n_268)
);

AOI21xp33_ASAP7_75t_L g299 ( 
.A1(n_268),
.A2(n_282),
.B(n_285),
.Y(n_299)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_132),
.Y(n_269)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_269),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_149),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_212),
.B(n_208),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_131),
.Y(n_274)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_274),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_177),
.Y(n_275)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_275),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_145),
.A2(n_150),
.B1(n_159),
.B2(n_203),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_277),
.A2(n_281),
.B1(n_293),
.B2(n_213),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_138),
.B(n_205),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_278),
.B(n_279),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_143),
.B(n_191),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_150),
.A2(n_159),
.B1(n_203),
.B2(n_190),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_132),
.B(n_191),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_171),
.A2(n_172),
.B1(n_184),
.B2(n_152),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_131),
.B(n_141),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_286),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_190),
.B(n_141),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_217),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_152),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_287),
.B(n_291),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_182),
.B(n_184),
.Y(n_288)
);

AND2x2_ASAP7_75t_SL g315 ( 
.A(n_288),
.B(n_289),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_182),
.B(n_186),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_200),
.Y(n_290)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_290),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_186),
.B(n_199),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_199),
.B(n_194),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_294),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_189),
.A2(n_71),
.B1(n_69),
.B2(n_176),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_200),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_301),
.A2(n_321),
.B1(n_252),
.B2(n_251),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_305),
.B(n_224),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_268),
.A2(n_292),
.B1(n_219),
.B2(n_270),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_306),
.A2(n_307),
.B1(n_333),
.B2(n_305),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_270),
.A2(n_234),
.B1(n_225),
.B2(n_245),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_316),
.A2(n_338),
.B(n_300),
.Y(n_351)
);

FAx1_ASAP7_75t_SL g322 ( 
.A(n_235),
.B(n_260),
.CI(n_247),
.CON(n_322),
.SN(n_322)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_322),
.B(n_341),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_253),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_327),
.B(n_334),
.Y(n_357)
);

O2A1O1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_264),
.A2(n_242),
.B(n_282),
.C(n_241),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_329),
.A2(n_304),
.B(n_311),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_224),
.A2(n_264),
.B1(n_240),
.B2(n_233),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_285),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_257),
.B(n_227),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_236),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_346),
.B(n_274),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_351),
.A2(n_358),
.B(n_362),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_315),
.B(n_229),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_352),
.B(n_360),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_353),
.A2(n_371),
.B1(n_373),
.B2(n_380),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_299),
.B(n_288),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_354),
.B(n_361),
.Y(n_400)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_295),
.Y(n_355)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_355),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_326),
.B(n_271),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_356),
.B(n_363),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_332),
.A2(n_250),
.B1(n_246),
.B2(n_248),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_314),
.Y(n_359)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_359),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_289),
.Y(n_360)
);

NAND2xp33_ASAP7_75t_SL g362 ( 
.A(n_337),
.B(n_222),
.Y(n_362)
);

AND2x2_ASAP7_75t_SL g363 ( 
.A(n_306),
.B(n_291),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_332),
.A2(n_238),
.B1(n_259),
.B2(n_262),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_365),
.A2(n_388),
.B(n_328),
.Y(n_427)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_295),
.Y(n_366)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_366),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_296),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_367),
.B(n_374),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_301),
.A2(n_269),
.B1(n_263),
.B2(n_244),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_368),
.A2(n_376),
.B1(n_382),
.B2(n_310),
.Y(n_405)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_298),
.Y(n_369)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_369),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_326),
.B(n_323),
.C(n_315),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_370),
.B(n_383),
.C(n_384),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_320),
.A2(n_261),
.B1(n_232),
.B2(n_275),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_372),
.A2(n_310),
.B1(n_339),
.B2(n_349),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_338),
.A2(n_254),
.B1(n_255),
.B2(n_237),
.Y(n_373)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_340),
.Y(n_375)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_375),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_315),
.A2(n_228),
.B1(n_256),
.B2(n_226),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_298),
.Y(n_377)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_377),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_302),
.B(n_228),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_379),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_322),
.B(n_302),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_316),
.A2(n_347),
.B1(n_319),
.B2(n_329),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_347),
.A2(n_326),
.B1(n_322),
.B2(n_323),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_381),
.B(n_389),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_330),
.A2(n_303),
.B1(n_350),
.B2(n_327),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_297),
.B(n_318),
.C(n_313),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_313),
.B(n_350),
.C(n_325),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_317),
.B(n_325),
.C(n_343),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_385),
.B(n_387),
.C(n_342),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_304),
.B(n_346),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_386),
.B(n_390),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_317),
.B(n_343),
.C(n_336),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_308),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_311),
.B(n_331),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_340),
.B(n_336),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_391),
.B(n_392),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_324),
.A2(n_310),
.B1(n_344),
.B2(n_314),
.Y(n_392)
);

OAI21xp33_ASAP7_75t_L g393 ( 
.A1(n_309),
.A2(n_345),
.B(n_324),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_345),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_308),
.Y(n_394)
);

INVx13_ASAP7_75t_L g412 ( 
.A(n_394),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_391),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_395),
.B(n_417),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_309),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_396),
.B(n_422),
.C(n_387),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_388),
.A2(n_362),
.B(n_357),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_397),
.A2(n_410),
.B(n_416),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_401),
.B(n_405),
.Y(n_431)
);

OA21x2_ASAP7_75t_L g404 ( 
.A1(n_363),
.A2(n_331),
.B(n_312),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_404),
.B(n_408),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_357),
.B(n_335),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_378),
.B(n_335),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_409),
.B(n_411),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_386),
.A2(n_348),
.B(n_328),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_360),
.B(n_379),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_352),
.B(n_342),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_413),
.B(n_385),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_382),
.Y(n_417)
);

XNOR2x1_ASAP7_75t_L g443 ( 
.A(n_420),
.B(n_354),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_370),
.B(n_312),
.C(n_344),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_427),
.A2(n_365),
.B(n_351),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_374),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_430),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_384),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_429),
.Y(n_432)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_432),
.Y(n_480)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_429),
.Y(n_434)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_434),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_398),
.B(n_363),
.Y(n_435)
);

CKINVDCx14_ASAP7_75t_R g468 ( 
.A(n_435),
.Y(n_468)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_406),
.Y(n_436)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_436),
.Y(n_477)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_403),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_437),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_399),
.B(n_354),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_439),
.B(n_451),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_398),
.B(n_363),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_441),
.B(n_445),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_442),
.B(n_443),
.C(n_446),
.Y(n_473)
);

NOR2x1_ASAP7_75t_R g479 ( 
.A(n_444),
.B(n_401),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_402),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_414),
.B(n_356),
.C(n_380),
.Y(n_446)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_403),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_448),
.A2(n_450),
.B1(n_452),
.B2(n_453),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_367),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_449),
.Y(n_471)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_419),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_397),
.A2(n_364),
.B(n_353),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_419),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_417),
.A2(n_361),
.B1(n_353),
.B2(n_373),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_406),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_454),
.A2(n_461),
.B1(n_462),
.B2(n_377),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_418),
.A2(n_368),
.B1(n_364),
.B2(n_376),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_456),
.A2(n_457),
.B1(n_400),
.B2(n_404),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_418),
.A2(n_358),
.B1(n_383),
.B2(n_369),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_402),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_458),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_411),
.B(n_428),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_459),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_396),
.B(n_356),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_420),
.C(n_422),
.Y(n_474)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_421),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_464),
.A2(n_475),
.B1(n_491),
.B2(n_453),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_414),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_465),
.B(n_472),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_432),
.A2(n_423),
.B1(n_395),
.B2(n_415),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_466),
.A2(n_483),
.B1(n_431),
.B2(n_440),
.Y(n_492)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_469),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_423),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_474),
.B(n_479),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_456),
.A2(n_400),
.B1(n_404),
.B2(n_427),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_446),
.B(n_399),
.C(n_400),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_478),
.B(n_481),
.C(n_482),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_399),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_439),
.B(n_451),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_434),
.A2(n_415),
.B1(n_416),
.B2(n_400),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_447),
.B(n_413),
.C(n_407),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_486),
.C(n_487),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_407),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_431),
.B(n_408),
.C(n_404),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_431),
.B(n_409),
.C(n_424),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_490),
.B(n_444),
.C(n_424),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_457),
.A2(n_405),
.B1(n_371),
.B2(n_421),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_492),
.A2(n_505),
.B1(n_513),
.B2(n_516),
.Y(n_530)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_477),
.Y(n_493)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_493),
.Y(n_528)
);

XOR2x2_ASAP7_75t_L g494 ( 
.A(n_472),
.B(n_435),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_500),
.Y(n_524)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_485),
.Y(n_495)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_495),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_497),
.A2(n_433),
.B1(n_488),
.B2(n_464),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_465),
.B(n_474),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_470),
.B(n_458),
.Y(n_501)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_501),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_471),
.B(n_438),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_502),
.B(n_506),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_463),
.B(n_445),
.Y(n_503)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_503),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_483),
.A2(n_467),
.B1(n_466),
.B2(n_468),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_476),
.B(n_390),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_489),
.Y(n_508)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_508),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_487),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_509),
.B(n_511),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_510),
.B(n_515),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_480),
.B(n_455),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_484),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_512),
.B(n_514),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_490),
.A2(n_440),
.B1(n_433),
.B2(n_455),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_486),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_491),
.B(n_441),
.Y(n_515)
);

FAx1_ASAP7_75t_SL g516 ( 
.A(n_478),
.B(n_488),
.CI(n_482),
.CON(n_516),
.SN(n_516)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_517),
.A2(n_513),
.B1(n_510),
.B2(n_511),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_501),
.A2(n_475),
.B(n_479),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_518),
.A2(n_519),
.B(n_520),
.Y(n_538)
);

BUFx12f_ASAP7_75t_SL g519 ( 
.A(n_516),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_503),
.A2(n_410),
.B(n_473),
.Y(n_520)
);

A2O1A1Ixp33_ASAP7_75t_SL g521 ( 
.A1(n_492),
.A2(n_461),
.B(n_452),
.C(n_450),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_521),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_505),
.A2(n_473),
.B(n_437),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_526),
.A2(n_532),
.B(n_507),
.Y(n_544)
);

BUFx12f_ASAP7_75t_SL g532 ( 
.A(n_516),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_526),
.B(n_500),
.C(n_504),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_535),
.B(n_539),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_527),
.A2(n_496),
.B1(n_509),
.B2(n_515),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_536),
.A2(n_541),
.B1(n_533),
.B2(n_520),
.Y(n_554)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_529),
.Y(n_537)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_537),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_523),
.B(n_504),
.C(n_499),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_540),
.A2(n_525),
.B1(n_533),
.B2(n_518),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_530),
.A2(n_494),
.B1(n_507),
.B2(n_499),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_517),
.B(n_498),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_542),
.B(n_543),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_530),
.B(n_498),
.Y(n_543)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_544),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_523),
.B(n_481),
.C(n_425),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_545),
.B(n_547),
.C(n_548),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_522),
.B(n_425),
.C(n_448),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_524),
.B(n_525),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_524),
.B(n_493),
.C(n_426),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_549),
.B(n_521),
.C(n_528),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_550),
.B(n_556),
.Y(n_563)
);

OA21x2_ASAP7_75t_L g552 ( 
.A1(n_536),
.A2(n_519),
.B(n_532),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_552),
.A2(n_521),
.B1(n_348),
.B2(n_436),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_554),
.B(n_562),
.Y(n_572)
);

AOI22x1_ASAP7_75t_L g555 ( 
.A1(n_538),
.A2(n_546),
.B1(n_521),
.B2(n_548),
.Y(n_555)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_555),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_547),
.A2(n_531),
.B1(n_528),
.B2(n_534),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_535),
.B(n_366),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_559),
.B(n_560),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_549),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_561),
.A2(n_541),
.B(n_543),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_564),
.A2(n_565),
.B(n_551),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g565 ( 
.A1(n_557),
.A2(n_539),
.B(n_545),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_550),
.B(n_542),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_567),
.B(n_568),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_553),
.B(n_426),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_SL g578 ( 
.A1(n_570),
.A2(n_355),
.B(n_412),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_552),
.B(n_359),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_571),
.B(n_566),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_573),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_575),
.B(n_576),
.C(n_578),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_572),
.B(n_558),
.C(n_551),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_564),
.A2(n_562),
.B(n_552),
.Y(n_577)
);

A2O1A1O1Ixp25_ASAP7_75t_L g581 ( 
.A1(n_577),
.A2(n_569),
.B(n_555),
.C(n_572),
.D(n_568),
.Y(n_581)
);

INVxp67_ASAP7_75t_SL g579 ( 
.A(n_563),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_579),
.B(n_570),
.C(n_558),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_581),
.B(n_583),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_574),
.B(n_454),
.C(n_392),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_584),
.B(n_389),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_580),
.A2(n_412),
.B(n_375),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_586),
.B(n_582),
.C(n_394),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_587),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_588),
.B(n_585),
.C(n_589),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_590),
.B(n_339),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_591),
.B(n_349),
.Y(n_592)
);


endmodule