module fake_jpeg_8877_n_334 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_31),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_27),
.B1(n_30),
.B2(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_18),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_18),
.B(n_2),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_50),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx5_ASAP7_75t_SL g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx5_ASAP7_75t_SL g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_62),
.Y(n_72)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_65),
.B1(n_27),
.B2(n_33),
.Y(n_71)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_63),
.B(n_19),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_43),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_71),
.A2(n_37),
.B1(n_33),
.B2(n_22),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_76),
.B(n_77),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_45),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_79),
.A2(n_22),
.B(n_25),
.Y(n_120)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_85),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_39),
.C(n_44),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_37),
.Y(n_114)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_87),
.Y(n_121)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_95),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_60),
.Y(n_103)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_39),
.B1(n_35),
.B2(n_58),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_85),
.B1(n_41),
.B2(n_91),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_74),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_100),
.B(n_101),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_74),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_30),
.B1(n_33),
.B2(n_22),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_102),
.A2(n_111),
.B1(n_112),
.B2(n_119),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_103),
.B(n_106),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_35),
.B1(n_48),
.B2(n_47),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_125)
);

AOI32xp33_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_59),
.A3(n_41),
.B1(n_30),
.B2(n_55),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_107),
.C(n_114),
.Y(n_151)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_44),
.C(n_39),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_35),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_43),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_77),
.A2(n_41),
.B1(n_37),
.B2(n_66),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_118),
.B1(n_73),
.B2(n_34),
.Y(n_134)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_34),
.A3(n_19),
.B1(n_28),
.B2(n_25),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_76),
.A2(n_67),
.B(n_19),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_25),
.B(n_21),
.Y(n_146)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_128),
.B1(n_132),
.B2(n_139),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_41),
.B1(n_57),
.B2(n_78),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_43),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_142),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_SL g178 ( 
.A1(n_134),
.A2(n_26),
.B(n_23),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_98),
.A2(n_73),
.B1(n_80),
.B2(n_78),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_135),
.A2(n_150),
.B1(n_97),
.B2(n_101),
.Y(n_157)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_137),
.B(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_105),
.B1(n_114),
.B2(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_120),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_87),
.B1(n_80),
.B2(n_33),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_149),
.B1(n_23),
.B2(n_26),
.Y(n_166)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_144),
.B(n_145),
.Y(n_179)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_146),
.A2(n_121),
.B(n_96),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_57),
.C(n_40),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_70),
.C(n_123),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_40),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_100),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_118),
.A2(n_40),
.B1(n_34),
.B2(n_28),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_40),
.B1(n_21),
.B2(n_28),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_146),
.B(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_160),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_165),
.B1(n_178),
.B2(n_125),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_140),
.B(n_106),
.Y(n_158)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_110),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_167),
.C(n_169),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_172),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_136),
.A2(n_109),
.B1(n_97),
.B2(n_40),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_166),
.A2(n_168),
.B1(n_23),
.B2(n_29),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_152),
.A2(n_108),
.B1(n_29),
.B2(n_26),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_108),
.C(n_20),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_142),
.B(n_20),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_170),
.B(n_177),
.CI(n_32),
.CON(n_203),
.SN(n_203)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_140),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_171),
.A2(n_174),
.B(n_175),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_127),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_2),
.Y(n_174)
);

NAND2xp33_ASAP7_75t_SL g175 ( 
.A(n_136),
.B(n_2),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_134),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_176),
.A2(n_180),
.B(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_32),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_139),
.C(n_132),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_192),
.C(n_197),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_180),
.A2(n_129),
.B1(n_143),
.B2(n_137),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_186),
.A2(n_187),
.B(n_203),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_200),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_129),
.B(n_135),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_189),
.A2(n_193),
.B(n_198),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_179),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_190),
.B(n_196),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_128),
.Y(n_192)
);

AOI21x1_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_149),
.B(n_150),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_144),
.C(n_145),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_130),
.B(n_14),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_161),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_20),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_167),
.C(n_165),
.Y(n_215)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_204),
.Y(n_218)
);

OAI22x1_ASAP7_75t_SL g205 ( 
.A1(n_156),
.A2(n_141),
.B1(n_24),
.B2(n_32),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_3),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_156),
.A2(n_131),
.B1(n_29),
.B2(n_24),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_206),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_160),
.A2(n_24),
.B1(n_32),
.B2(n_11),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_157),
.A2(n_131),
.B1(n_24),
.B2(n_5),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_172),
.B1(n_153),
.B2(n_163),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_191),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_225),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_177),
.Y(n_212)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_192),
.C(n_201),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_154),
.B(n_168),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_216),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_166),
.B1(n_158),
.B2(n_174),
.Y(n_219)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_174),
.B1(n_4),
.B2(n_5),
.Y(n_220)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_9),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_222),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_9),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_3),
.Y(n_223)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_224)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_207),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_227),
.B(n_228),
.Y(n_253)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_183),
.B(n_209),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_230),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_182),
.B(n_9),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_184),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_199),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_234),
.B1(n_193),
.B2(n_209),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_188),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_235),
.Y(n_237)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_226),
.B(n_216),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_245),
.C(n_246),
.Y(n_261)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

FAx1_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_187),
.CI(n_189),
.CON(n_242),
.SN(n_242)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_184),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_251),
.C(n_254),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_203),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_203),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_194),
.C(n_6),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_258),
.C(n_220),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_13),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_249),
.A2(n_233),
.B1(n_228),
.B2(n_232),
.Y(n_259)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_259),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_227),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_265),
.Y(n_282)
);

INVxp67_ASAP7_75t_SL g264 ( 
.A(n_241),
.Y(n_264)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_253),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_270),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_269),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_222),
.C(n_231),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_274),
.C(n_261),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_212),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_230),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_271),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_234),
.B1(n_213),
.B2(n_218),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_237),
.B1(n_257),
.B2(n_238),
.Y(n_281)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_273),
.B(n_276),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_218),
.C(n_211),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_271),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_263),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_285),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_251),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_242),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_258),
.C(n_244),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_286),
.C(n_291),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_217),
.B(n_250),
.Y(n_284)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_254),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_272),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_291),
.B(n_229),
.Y(n_292)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_277),
.A2(n_275),
.B1(n_262),
.B2(n_260),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_294),
.A2(n_287),
.B(n_288),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_242),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_283),
.C(n_280),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_286),
.C(n_244),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_301),
.Y(n_313)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_270),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_303),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_223),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_219),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_217),
.B(n_235),
.Y(n_309)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_293),
.B(n_268),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_308),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

OAI21x1_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_295),
.B(n_300),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_293),
.B(n_224),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_7),
.B(n_8),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_13),
.Y(n_312)
);

AOI21xp33_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_7),
.B(n_8),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_SL g324 ( 
.A1(n_316),
.A2(n_322),
.B(n_8),
.C(n_10),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_305),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_317),
.B(n_318),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_296),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_14),
.Y(n_327)
);

AOI21x1_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_310),
.B(n_314),
.Y(n_323)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_324),
.C(n_327),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_308),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_325),
.A2(n_321),
.B(n_315),
.Y(n_329)
);

A2O1A1O1Ixp25_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_324),
.B(n_326),
.C(n_15),
.D(n_16),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_14),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_328),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_15),
.B(n_6),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_333),
.B(n_15),
.Y(n_334)
);


endmodule