module fake_netlist_6_802_n_4303 (n_992, n_1, n_801, n_1234, n_1199, n_741, n_1027, n_1351, n_625, n_1189, n_223, n_1212, n_226, n_208, n_68, n_726, n_212, n_700, n_50, n_1307, n_1038, n_578, n_1003, n_365, n_168, n_1237, n_1061, n_1357, n_77, n_783, n_798, n_188, n_509, n_1342, n_245, n_1209, n_1348, n_1387, n_677, n_805, n_1151, n_396, n_350, n_78, n_1380, n_442, n_480, n_142, n_1009, n_62, n_1160, n_883, n_1238, n_1032, n_1247, n_893, n_1099, n_1264, n_1192, n_471, n_424, n_1370, n_369, n_287, n_415, n_830, n_65, n_230, n_461, n_873, n_141, n_383, n_1285, n_1371, n_200, n_447, n_1172, n_852, n_71, n_229, n_1393, n_1078, n_250, n_544, n_1140, n_35, n_1263, n_836, n_375, n_522, n_1261, n_945, n_1143, n_1232, n_616, n_658, n_1119, n_428, n_1300, n_641, n_822, n_693, n_1313, n_1056, n_758, n_516, n_1163, n_1180, n_943, n_491, n_42, n_772, n_1344, n_666, n_371, n_940, n_770, n_567, n_405, n_213, n_538, n_1106, n_886, n_343, n_953, n_1094, n_1345, n_494, n_539, n_493, n_155, n_45, n_454, n_638, n_1211, n_381, n_887, n_112, n_1280, n_713, n_1400, n_126, n_58, n_976, n_224, n_48, n_734, n_1088, n_196, n_1231, n_917, n_574, n_9, n_907, n_6, n_14, n_659, n_407, n_913, n_808, n_867, n_1230, n_473, n_1193, n_1054, n_559, n_1333, n_44, n_163, n_281, n_551, n_699, n_564, n_451, n_824, n_279, n_686, n_757, n_594, n_577, n_166, n_619, n_1367, n_1336, n_521, n_572, n_395, n_813, n_323, n_606, n_818, n_1123, n_1309, n_92, n_513, n_645, n_1381, n_331, n_916, n_483, n_102, n_608, n_261, n_630, n_32, n_541, n_512, n_121, n_433, n_792, n_476, n_2, n_1328, n_219, n_264, n_263, n_1162, n_860, n_788, n_939, n_821, n_938, n_1302, n_1068, n_329, n_982, n_549, n_1075, n_408, n_932, n_61, n_237, n_243, n_979, n_905, n_117, n_175, n_322, n_993, n_689, n_354, n_1330, n_134, n_1278, n_547, n_558, n_1064, n_1396, n_634, n_136, n_966, n_764, n_692, n_733, n_1233, n_1289, n_487, n_241, n_30, n_1107, n_1014, n_1290, n_882, n_1354, n_586, n_423, n_318, n_1111, n_715, n_1251, n_1265, n_88, n_530, n_277, n_618, n_1297, n_1312, n_199, n_1167, n_1359, n_674, n_871, n_922, n_268, n_1335, n_210, n_1069, n_5, n_612, n_178, n_247, n_1165, n_355, n_702, n_347, n_1175, n_328, n_1386, n_429, n_1012, n_195, n_780, n_675, n_903, n_286, n_254, n_242, n_835, n_1214, n_928, n_47, n_690, n_850, n_816, n_1157, n_1188, n_877, n_604, n_825, n_728, n_1063, n_26, n_55, n_267, n_1124, n_515, n_598, n_696, n_961, n_437, n_1082, n_1317, n_593, n_514, n_687, n_697, n_890, n_637, n_295, n_701, n_950, n_388, n_190, n_484, n_170, n_891, n_949, n_678, n_283, n_91, n_507, n_968, n_909, n_1369, n_881, n_1008, n_760, n_590, n_63, n_362, n_148, n_161, n_22, n_462, n_1033, n_1052, n_1296, n_304, n_694, n_1294, n_125, n_297, n_595, n_627, n_524, n_342, n_1044, n_1391, n_449, n_131, n_1208, n_1164, n_1295, n_1072, n_495, n_815, n_1100, n_585, n_840, n_874, n_1128, n_382, n_673, n_1071, n_1067, n_898, n_255, n_284, n_865, n_925, n_1101, n_15, n_1026, n_38, n_289, n_1364, n_615, n_1249, n_59, n_1293, n_1127, n_320, n_108, n_639, n_963, n_794, n_727, n_894, n_685, n_353, n_605, n_826, n_872, n_1139, n_86, n_104, n_718, n_1018, n_1366, n_542, n_847, n_644, n_682, n_851, n_305, n_72, n_996, n_532, n_173, n_1308, n_1376, n_413, n_791, n_510, n_837, n_79, n_948, n_704, n_977, n_1005, n_536, n_622, n_147, n_581, n_765, n_432, n_987, n_1340, n_631, n_720, n_153, n_842, n_156, n_145, n_843, n_656, n_989, n_1277, n_797, n_1246, n_899, n_189, n_738, n_1304, n_1035, n_294, n_499, n_705, n_11, n_1004, n_1176, n_1022, n_614, n_529, n_425, n_684, n_1181, n_37, n_486, n_947, n_1117, n_1087, n_648, n_657, n_1049, n_803, n_290, n_118, n_926, n_927, n_919, n_478, n_929, n_107, n_1228, n_417, n_446, n_89, n_777, n_1299, n_272, n_526, n_1183, n_1384, n_69, n_293, n_53, n_458, n_1070, n_998, n_16, n_717, n_18, n_154, n_1383, n_1178, n_98, n_1073, n_1000, n_796, n_252, n_1195, n_184, n_552, n_1358, n_1388, n_216, n_912, n_745, n_1284, n_1142, n_716, n_623, n_1048, n_1201, n_1398, n_884, n_1395, n_731, n_755, n_931, n_1021, n_474, n_527, n_683, n_811, n_1207, n_312, n_1368, n_66, n_958, n_292, n_1250, n_100, n_1137, n_880, n_889, n_150, n_589, n_1310, n_819, n_1363, n_1334, n_767, n_1314, n_600, n_964, n_831, n_477, n_954, n_864, n_1110, n_399, n_124, n_1382, n_211, n_1372, n_231, n_40, n_505, n_319, n_1339, n_537, n_311, n_10, n_403, n_1080, n_723, n_596, n_123, n_546, n_562, n_1141, n_1268, n_386, n_1220, n_556, n_162, n_1136, n_128, n_1125, n_970, n_642, n_995, n_276, n_1159, n_1092, n_441, n_221, n_1060, n_444, n_146, n_1252, n_1223, n_303, n_511, n_193, n_1286, n_1053, n_416, n_520, n_418, n_1093, n_113, n_4, n_266, n_296, n_775, n_651, n_1153, n_439, n_217, n_518, n_1185, n_453, n_215, n_914, n_759, n_426, n_317, n_90, n_54, n_488, n_497, n_773, n_920, n_99, n_1374, n_1315, n_13, n_1224, n_1135, n_1169, n_1179, n_401, n_324, n_335, n_463, n_1243, n_848, n_120, n_301, n_274, n_1096, n_1091, n_36, n_1267, n_1281, n_983, n_427, n_496, n_906, n_1390, n_688, n_1077, n_351, n_259, n_177, n_385, n_1323, n_858, n_1331, n_613, n_736, n_501, n_956, n_960, n_663, n_856, n_379, n_778, n_1134, n_410, n_1129, n_554, n_602, n_664, n_171, n_169, n_435, n_793, n_326, n_587, n_580, n_762, n_1030, n_1202, n_465, n_1079, n_341, n_828, n_607, n_316, n_419, n_28, n_1103, n_144, n_1203, n_820, n_951, n_106, n_725, n_952, n_999, n_358, n_1254, n_160, n_186, n_0, n_368, n_575, n_994, n_732, n_974, n_392, n_724, n_1020, n_1042, n_628, n_1273, n_557, n_349, n_617, n_845, n_807, n_1036, n_140, n_1138, n_1275, n_485, n_67, n_443, n_892, n_768, n_421, n_238, n_1095, n_202, n_597, n_280, n_1270, n_1187, n_610, n_1024, n_198, n_179, n_248, n_517, n_667, n_1206, n_621, n_1037, n_1397, n_1279, n_1115, n_750, n_901, n_468, n_923, n_504, n_183, n_1015, n_466, n_1057, n_603, n_991, n_235, n_1126, n_340, n_710, n_1108, n_1182, n_1298, n_39, n_73, n_785, n_746, n_609, n_101, n_167, n_1356, n_127, n_1168, n_1216, n_133, n_1320, n_96, n_1316, n_1287, n_302, n_380, n_137, n_20, n_1190, n_397, n_122, n_34, n_1262, n_218, n_1213, n_70, n_1350, n_172, n_1272, n_239, n_97, n_782, n_490, n_220, n_809, n_1043, n_986, n_80, n_1081, n_402, n_352, n_800, n_1084, n_1171, n_460, n_1361, n_662, n_374, n_1152, n_450, n_921, n_1346, n_711, n_579, n_1352, n_937, n_370, n_650, n_1046, n_1145, n_330, n_1121, n_1102, n_972, n_258, n_456, n_1332, n_260, n_313, n_624, n_962, n_1041, n_565, n_356, n_936, n_1288, n_1186, n_1062, n_885, n_896, n_83, n_654, n_411, n_152, n_1222, n_599, n_776, n_321, n_105, n_227, n_204, n_482, n_934, n_420, n_1341, n_394, n_164, n_23, n_942, n_543, n_1271, n_1355, n_1225, n_325, n_804, n_464, n_533, n_806, n_879, n_959, n_584, n_244, n_1343, n_76, n_548, n_94, n_282, n_833, n_523, n_1319, n_707, n_345, n_799, n_1155, n_139, n_41, n_273, n_787, n_1146, n_159, n_1086, n_1066, n_157, n_1282, n_550, n_275, n_652, n_560, n_1241, n_1321, n_569, n_737, n_1318, n_1235, n_1229, n_306, n_1292, n_1373, n_21, n_346, n_3, n_1029, n_790, n_138, n_1210, n_49, n_299, n_1248, n_902, n_333, n_1047, n_1385, n_431, n_24, n_459, n_1269, n_502, n_672, n_1257, n_285, n_1375, n_85, n_655, n_706, n_1045, n_786, n_1236, n_834, n_19, n_29, n_75, n_743, n_766, n_430, n_1325, n_1002, n_545, n_489, n_251, n_1019, n_636, n_729, n_110, n_151, n_876, n_774, n_1337, n_660, n_438, n_1360, n_1200, n_479, n_1353, n_869, n_1154, n_1113, n_646, n_528, n_391, n_1098, n_1329, n_817, n_262, n_187, n_897, n_846, n_841, n_1001, n_508, n_1050, n_1177, n_332, n_1150, n_398, n_1191, n_566, n_1023, n_1076, n_1118, n_194, n_57, n_1007, n_1378, n_855, n_52, n_591, n_1377, n_256, n_853, n_440, n_695, n_875, n_209, n_367, n_680, n_661, n_278, n_1256, n_671, n_7, n_933, n_740, n_703, n_978, n_384, n_1291, n_1217, n_751, n_749, n_310, n_1324, n_1399, n_969, n_988, n_1065, n_84, n_1401, n_1255, n_568, n_143, n_180, n_1204, n_823, n_1132, n_643, n_233, n_698, n_1074, n_1394, n_1327, n_1326, n_739, n_400, n_955, n_337, n_1379, n_214, n_246, n_1338, n_1097, n_935, n_781, n_789, n_1130, n_181, n_182, n_573, n_769, n_676, n_327, n_1120, n_832, n_555, n_389, n_814, n_669, n_176, n_114, n_300, n_222, n_747, n_74, n_1389, n_1105, n_721, n_742, n_535, n_691, n_372, n_111, n_314, n_378, n_1196, n_377, n_863, n_601, n_338, n_1283, n_918, n_748, n_506, n_1114, n_56, n_763, n_1147, n_360, n_119, n_957, n_895, n_866, n_1227, n_191, n_387, n_452, n_744, n_971, n_946, n_344, n_761, n_1303, n_1205, n_1258, n_1392, n_174, n_1173, n_525, n_1116, n_611, n_1219, n_8, n_1174, n_1016, n_1347, n_795, n_1221, n_1245, n_838, n_129, n_647, n_197, n_844, n_17, n_448, n_1017, n_1083, n_109, n_445, n_930, n_888, n_1112, n_234, n_910, n_911, n_82, n_27, n_236, n_653, n_752, n_908, n_944, n_576, n_1028, n_472, n_270, n_414, n_563, n_1011, n_1215, n_25, n_93, n_839, n_708, n_668, n_626, n_990, n_779, n_1104, n_854, n_1058, n_498, n_1122, n_870, n_904, n_1253, n_709, n_1266, n_366, n_103, n_1109, n_185, n_712, n_348, n_1276, n_376, n_390, n_1148, n_31, n_334, n_1161, n_1085, n_232, n_46, n_1239, n_771, n_470, n_475, n_924, n_298, n_492, n_1149, n_265, n_1184, n_228, n_719, n_455, n_363, n_1090, n_592, n_829, n_1156, n_1362, n_393, n_984, n_503, n_132, n_868, n_570, n_859, n_406, n_735, n_878, n_620, n_130, n_519, n_307, n_469, n_1218, n_500, n_981, n_714, n_1349, n_291, n_1144, n_357, n_985, n_481, n_997, n_1301, n_802, n_561, n_33, n_980, n_1306, n_1198, n_436, n_116, n_409, n_1244, n_240, n_756, n_810, n_1133, n_635, n_95, n_1194, n_1051, n_253, n_583, n_249, n_201, n_1039, n_1034, n_1158, n_754, n_941, n_975, n_1031, n_115, n_1305, n_553, n_43, n_849, n_753, n_467, n_269, n_359, n_973, n_1055, n_582, n_861, n_857, n_967, n_571, n_271, n_404, n_158, n_206, n_679, n_633, n_1170, n_665, n_588, n_225, n_1260, n_308, n_309, n_1010, n_149, n_1040, n_915, n_632, n_1166, n_812, n_1131, n_534, n_1006, n_373, n_87, n_257, n_730, n_1311, n_670, n_203, n_207, n_1089, n_1365, n_205, n_1242, n_681, n_1226, n_1274, n_412, n_640, n_1322, n_81, n_965, n_339, n_784, n_315, n_434, n_64, n_288, n_1059, n_1197, n_422, n_722, n_862, n_135, n_165, n_540, n_457, n_364, n_629, n_900, n_531, n_827, n_60, n_361, n_1025, n_336, n_12, n_1013, n_1259, n_192, n_51, n_649, n_1240, n_4303);

input n_992;
input n_1;
input n_801;
input n_1234;
input n_1199;
input n_741;
input n_1027;
input n_1351;
input n_625;
input n_1189;
input n_223;
input n_1212;
input n_226;
input n_208;
input n_68;
input n_726;
input n_212;
input n_700;
input n_50;
input n_1307;
input n_1038;
input n_578;
input n_1003;
input n_365;
input n_168;
input n_1237;
input n_1061;
input n_1357;
input n_77;
input n_783;
input n_798;
input n_188;
input n_509;
input n_1342;
input n_245;
input n_1209;
input n_1348;
input n_1387;
input n_677;
input n_805;
input n_1151;
input n_396;
input n_350;
input n_78;
input n_1380;
input n_442;
input n_480;
input n_142;
input n_1009;
input n_62;
input n_1160;
input n_883;
input n_1238;
input n_1032;
input n_1247;
input n_893;
input n_1099;
input n_1264;
input n_1192;
input n_471;
input n_424;
input n_1370;
input n_369;
input n_287;
input n_415;
input n_830;
input n_65;
input n_230;
input n_461;
input n_873;
input n_141;
input n_383;
input n_1285;
input n_1371;
input n_200;
input n_447;
input n_1172;
input n_852;
input n_71;
input n_229;
input n_1393;
input n_1078;
input n_250;
input n_544;
input n_1140;
input n_35;
input n_1263;
input n_836;
input n_375;
input n_522;
input n_1261;
input n_945;
input n_1143;
input n_1232;
input n_616;
input n_658;
input n_1119;
input n_428;
input n_1300;
input n_641;
input n_822;
input n_693;
input n_1313;
input n_1056;
input n_758;
input n_516;
input n_1163;
input n_1180;
input n_943;
input n_491;
input n_42;
input n_772;
input n_1344;
input n_666;
input n_371;
input n_940;
input n_770;
input n_567;
input n_405;
input n_213;
input n_538;
input n_1106;
input n_886;
input n_343;
input n_953;
input n_1094;
input n_1345;
input n_494;
input n_539;
input n_493;
input n_155;
input n_45;
input n_454;
input n_638;
input n_1211;
input n_381;
input n_887;
input n_112;
input n_1280;
input n_713;
input n_1400;
input n_126;
input n_58;
input n_976;
input n_224;
input n_48;
input n_734;
input n_1088;
input n_196;
input n_1231;
input n_917;
input n_574;
input n_9;
input n_907;
input n_6;
input n_14;
input n_659;
input n_407;
input n_913;
input n_808;
input n_867;
input n_1230;
input n_473;
input n_1193;
input n_1054;
input n_559;
input n_1333;
input n_44;
input n_163;
input n_281;
input n_551;
input n_699;
input n_564;
input n_451;
input n_824;
input n_279;
input n_686;
input n_757;
input n_594;
input n_577;
input n_166;
input n_619;
input n_1367;
input n_1336;
input n_521;
input n_572;
input n_395;
input n_813;
input n_323;
input n_606;
input n_818;
input n_1123;
input n_1309;
input n_92;
input n_513;
input n_645;
input n_1381;
input n_331;
input n_916;
input n_483;
input n_102;
input n_608;
input n_261;
input n_630;
input n_32;
input n_541;
input n_512;
input n_121;
input n_433;
input n_792;
input n_476;
input n_2;
input n_1328;
input n_219;
input n_264;
input n_263;
input n_1162;
input n_860;
input n_788;
input n_939;
input n_821;
input n_938;
input n_1302;
input n_1068;
input n_329;
input n_982;
input n_549;
input n_1075;
input n_408;
input n_932;
input n_61;
input n_237;
input n_243;
input n_979;
input n_905;
input n_117;
input n_175;
input n_322;
input n_993;
input n_689;
input n_354;
input n_1330;
input n_134;
input n_1278;
input n_547;
input n_558;
input n_1064;
input n_1396;
input n_634;
input n_136;
input n_966;
input n_764;
input n_692;
input n_733;
input n_1233;
input n_1289;
input n_487;
input n_241;
input n_30;
input n_1107;
input n_1014;
input n_1290;
input n_882;
input n_1354;
input n_586;
input n_423;
input n_318;
input n_1111;
input n_715;
input n_1251;
input n_1265;
input n_88;
input n_530;
input n_277;
input n_618;
input n_1297;
input n_1312;
input n_199;
input n_1167;
input n_1359;
input n_674;
input n_871;
input n_922;
input n_268;
input n_1335;
input n_210;
input n_1069;
input n_5;
input n_612;
input n_178;
input n_247;
input n_1165;
input n_355;
input n_702;
input n_347;
input n_1175;
input n_328;
input n_1386;
input n_429;
input n_1012;
input n_195;
input n_780;
input n_675;
input n_903;
input n_286;
input n_254;
input n_242;
input n_835;
input n_1214;
input n_928;
input n_47;
input n_690;
input n_850;
input n_816;
input n_1157;
input n_1188;
input n_877;
input n_604;
input n_825;
input n_728;
input n_1063;
input n_26;
input n_55;
input n_267;
input n_1124;
input n_515;
input n_598;
input n_696;
input n_961;
input n_437;
input n_1082;
input n_1317;
input n_593;
input n_514;
input n_687;
input n_697;
input n_890;
input n_637;
input n_295;
input n_701;
input n_950;
input n_388;
input n_190;
input n_484;
input n_170;
input n_891;
input n_949;
input n_678;
input n_283;
input n_91;
input n_507;
input n_968;
input n_909;
input n_1369;
input n_881;
input n_1008;
input n_760;
input n_590;
input n_63;
input n_362;
input n_148;
input n_161;
input n_22;
input n_462;
input n_1033;
input n_1052;
input n_1296;
input n_304;
input n_694;
input n_1294;
input n_125;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_1044;
input n_1391;
input n_449;
input n_131;
input n_1208;
input n_1164;
input n_1295;
input n_1072;
input n_495;
input n_815;
input n_1100;
input n_585;
input n_840;
input n_874;
input n_1128;
input n_382;
input n_673;
input n_1071;
input n_1067;
input n_898;
input n_255;
input n_284;
input n_865;
input n_925;
input n_1101;
input n_15;
input n_1026;
input n_38;
input n_289;
input n_1364;
input n_615;
input n_1249;
input n_59;
input n_1293;
input n_1127;
input n_320;
input n_108;
input n_639;
input n_963;
input n_794;
input n_727;
input n_894;
input n_685;
input n_353;
input n_605;
input n_826;
input n_872;
input n_1139;
input n_86;
input n_104;
input n_718;
input n_1018;
input n_1366;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_305;
input n_72;
input n_996;
input n_532;
input n_173;
input n_1308;
input n_1376;
input n_413;
input n_791;
input n_510;
input n_837;
input n_79;
input n_948;
input n_704;
input n_977;
input n_1005;
input n_536;
input n_622;
input n_147;
input n_581;
input n_765;
input n_432;
input n_987;
input n_1340;
input n_631;
input n_720;
input n_153;
input n_842;
input n_156;
input n_145;
input n_843;
input n_656;
input n_989;
input n_1277;
input n_797;
input n_1246;
input n_899;
input n_189;
input n_738;
input n_1304;
input n_1035;
input n_294;
input n_499;
input n_705;
input n_11;
input n_1004;
input n_1176;
input n_1022;
input n_614;
input n_529;
input n_425;
input n_684;
input n_1181;
input n_37;
input n_486;
input n_947;
input n_1117;
input n_1087;
input n_648;
input n_657;
input n_1049;
input n_803;
input n_290;
input n_118;
input n_926;
input n_927;
input n_919;
input n_478;
input n_929;
input n_107;
input n_1228;
input n_417;
input n_446;
input n_89;
input n_777;
input n_1299;
input n_272;
input n_526;
input n_1183;
input n_1384;
input n_69;
input n_293;
input n_53;
input n_458;
input n_1070;
input n_998;
input n_16;
input n_717;
input n_18;
input n_154;
input n_1383;
input n_1178;
input n_98;
input n_1073;
input n_1000;
input n_796;
input n_252;
input n_1195;
input n_184;
input n_552;
input n_1358;
input n_1388;
input n_216;
input n_912;
input n_745;
input n_1284;
input n_1142;
input n_716;
input n_623;
input n_1048;
input n_1201;
input n_1398;
input n_884;
input n_1395;
input n_731;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_683;
input n_811;
input n_1207;
input n_312;
input n_1368;
input n_66;
input n_958;
input n_292;
input n_1250;
input n_100;
input n_1137;
input n_880;
input n_889;
input n_150;
input n_589;
input n_1310;
input n_819;
input n_1363;
input n_1334;
input n_767;
input n_1314;
input n_600;
input n_964;
input n_831;
input n_477;
input n_954;
input n_864;
input n_1110;
input n_399;
input n_124;
input n_1382;
input n_211;
input n_1372;
input n_231;
input n_40;
input n_505;
input n_319;
input n_1339;
input n_537;
input n_311;
input n_10;
input n_403;
input n_1080;
input n_723;
input n_596;
input n_123;
input n_546;
input n_562;
input n_1141;
input n_1268;
input n_386;
input n_1220;
input n_556;
input n_162;
input n_1136;
input n_128;
input n_1125;
input n_970;
input n_642;
input n_995;
input n_276;
input n_1159;
input n_1092;
input n_441;
input n_221;
input n_1060;
input n_444;
input n_146;
input n_1252;
input n_1223;
input n_303;
input n_511;
input n_193;
input n_1286;
input n_1053;
input n_416;
input n_520;
input n_418;
input n_1093;
input n_113;
input n_4;
input n_266;
input n_296;
input n_775;
input n_651;
input n_1153;
input n_439;
input n_217;
input n_518;
input n_1185;
input n_453;
input n_215;
input n_914;
input n_759;
input n_426;
input n_317;
input n_90;
input n_54;
input n_488;
input n_497;
input n_773;
input n_920;
input n_99;
input n_1374;
input n_1315;
input n_13;
input n_1224;
input n_1135;
input n_1169;
input n_1179;
input n_401;
input n_324;
input n_335;
input n_463;
input n_1243;
input n_848;
input n_120;
input n_301;
input n_274;
input n_1096;
input n_1091;
input n_36;
input n_1267;
input n_1281;
input n_983;
input n_427;
input n_496;
input n_906;
input n_1390;
input n_688;
input n_1077;
input n_351;
input n_259;
input n_177;
input n_385;
input n_1323;
input n_858;
input n_1331;
input n_613;
input n_736;
input n_501;
input n_956;
input n_960;
input n_663;
input n_856;
input n_379;
input n_778;
input n_1134;
input n_410;
input n_1129;
input n_554;
input n_602;
input n_664;
input n_171;
input n_169;
input n_435;
input n_793;
input n_326;
input n_587;
input n_580;
input n_762;
input n_1030;
input n_1202;
input n_465;
input n_1079;
input n_341;
input n_828;
input n_607;
input n_316;
input n_419;
input n_28;
input n_1103;
input n_144;
input n_1203;
input n_820;
input n_951;
input n_106;
input n_725;
input n_952;
input n_999;
input n_358;
input n_1254;
input n_160;
input n_186;
input n_0;
input n_368;
input n_575;
input n_994;
input n_732;
input n_974;
input n_392;
input n_724;
input n_1020;
input n_1042;
input n_628;
input n_1273;
input n_557;
input n_349;
input n_617;
input n_845;
input n_807;
input n_1036;
input n_140;
input n_1138;
input n_1275;
input n_485;
input n_67;
input n_443;
input n_892;
input n_768;
input n_421;
input n_238;
input n_1095;
input n_202;
input n_597;
input n_280;
input n_1270;
input n_1187;
input n_610;
input n_1024;
input n_198;
input n_179;
input n_248;
input n_517;
input n_667;
input n_1206;
input n_621;
input n_1037;
input n_1397;
input n_1279;
input n_1115;
input n_750;
input n_901;
input n_468;
input n_923;
input n_504;
input n_183;
input n_1015;
input n_466;
input n_1057;
input n_603;
input n_991;
input n_235;
input n_1126;
input n_340;
input n_710;
input n_1108;
input n_1182;
input n_1298;
input n_39;
input n_73;
input n_785;
input n_746;
input n_609;
input n_101;
input n_167;
input n_1356;
input n_127;
input n_1168;
input n_1216;
input n_133;
input n_1320;
input n_96;
input n_1316;
input n_1287;
input n_302;
input n_380;
input n_137;
input n_20;
input n_1190;
input n_397;
input n_122;
input n_34;
input n_1262;
input n_218;
input n_1213;
input n_70;
input n_1350;
input n_172;
input n_1272;
input n_239;
input n_97;
input n_782;
input n_490;
input n_220;
input n_809;
input n_1043;
input n_986;
input n_80;
input n_1081;
input n_402;
input n_352;
input n_800;
input n_1084;
input n_1171;
input n_460;
input n_1361;
input n_662;
input n_374;
input n_1152;
input n_450;
input n_921;
input n_1346;
input n_711;
input n_579;
input n_1352;
input n_937;
input n_370;
input n_650;
input n_1046;
input n_1145;
input n_330;
input n_1121;
input n_1102;
input n_972;
input n_258;
input n_456;
input n_1332;
input n_260;
input n_313;
input n_624;
input n_962;
input n_1041;
input n_565;
input n_356;
input n_936;
input n_1288;
input n_1186;
input n_1062;
input n_885;
input n_896;
input n_83;
input n_654;
input n_411;
input n_152;
input n_1222;
input n_599;
input n_776;
input n_321;
input n_105;
input n_227;
input n_204;
input n_482;
input n_934;
input n_420;
input n_1341;
input n_394;
input n_164;
input n_23;
input n_942;
input n_543;
input n_1271;
input n_1355;
input n_1225;
input n_325;
input n_804;
input n_464;
input n_533;
input n_806;
input n_879;
input n_959;
input n_584;
input n_244;
input n_1343;
input n_76;
input n_548;
input n_94;
input n_282;
input n_833;
input n_523;
input n_1319;
input n_707;
input n_345;
input n_799;
input n_1155;
input n_139;
input n_41;
input n_273;
input n_787;
input n_1146;
input n_159;
input n_1086;
input n_1066;
input n_157;
input n_1282;
input n_550;
input n_275;
input n_652;
input n_560;
input n_1241;
input n_1321;
input n_569;
input n_737;
input n_1318;
input n_1235;
input n_1229;
input n_306;
input n_1292;
input n_1373;
input n_21;
input n_346;
input n_3;
input n_1029;
input n_790;
input n_138;
input n_1210;
input n_49;
input n_299;
input n_1248;
input n_902;
input n_333;
input n_1047;
input n_1385;
input n_431;
input n_24;
input n_459;
input n_1269;
input n_502;
input n_672;
input n_1257;
input n_285;
input n_1375;
input n_85;
input n_655;
input n_706;
input n_1045;
input n_786;
input n_1236;
input n_834;
input n_19;
input n_29;
input n_75;
input n_743;
input n_766;
input n_430;
input n_1325;
input n_1002;
input n_545;
input n_489;
input n_251;
input n_1019;
input n_636;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_1337;
input n_660;
input n_438;
input n_1360;
input n_1200;
input n_479;
input n_1353;
input n_869;
input n_1154;
input n_1113;
input n_646;
input n_528;
input n_391;
input n_1098;
input n_1329;
input n_817;
input n_262;
input n_187;
input n_897;
input n_846;
input n_841;
input n_1001;
input n_508;
input n_1050;
input n_1177;
input n_332;
input n_1150;
input n_398;
input n_1191;
input n_566;
input n_1023;
input n_1076;
input n_1118;
input n_194;
input n_57;
input n_1007;
input n_1378;
input n_855;
input n_52;
input n_591;
input n_1377;
input n_256;
input n_853;
input n_440;
input n_695;
input n_875;
input n_209;
input n_367;
input n_680;
input n_661;
input n_278;
input n_1256;
input n_671;
input n_7;
input n_933;
input n_740;
input n_703;
input n_978;
input n_384;
input n_1291;
input n_1217;
input n_751;
input n_749;
input n_310;
input n_1324;
input n_1399;
input n_969;
input n_988;
input n_1065;
input n_84;
input n_1401;
input n_1255;
input n_568;
input n_143;
input n_180;
input n_1204;
input n_823;
input n_1132;
input n_643;
input n_233;
input n_698;
input n_1074;
input n_1394;
input n_1327;
input n_1326;
input n_739;
input n_400;
input n_955;
input n_337;
input n_1379;
input n_214;
input n_246;
input n_1338;
input n_1097;
input n_935;
input n_781;
input n_789;
input n_1130;
input n_181;
input n_182;
input n_573;
input n_769;
input n_676;
input n_327;
input n_1120;
input n_832;
input n_555;
input n_389;
input n_814;
input n_669;
input n_176;
input n_114;
input n_300;
input n_222;
input n_747;
input n_74;
input n_1389;
input n_1105;
input n_721;
input n_742;
input n_535;
input n_691;
input n_372;
input n_111;
input n_314;
input n_378;
input n_1196;
input n_377;
input n_863;
input n_601;
input n_338;
input n_1283;
input n_918;
input n_748;
input n_506;
input n_1114;
input n_56;
input n_763;
input n_1147;
input n_360;
input n_119;
input n_957;
input n_895;
input n_866;
input n_1227;
input n_191;
input n_387;
input n_452;
input n_744;
input n_971;
input n_946;
input n_344;
input n_761;
input n_1303;
input n_1205;
input n_1258;
input n_1392;
input n_174;
input n_1173;
input n_525;
input n_1116;
input n_611;
input n_1219;
input n_8;
input n_1174;
input n_1016;
input n_1347;
input n_795;
input n_1221;
input n_1245;
input n_838;
input n_129;
input n_647;
input n_197;
input n_844;
input n_17;
input n_448;
input n_1017;
input n_1083;
input n_109;
input n_445;
input n_930;
input n_888;
input n_1112;
input n_234;
input n_910;
input n_911;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_908;
input n_944;
input n_576;
input n_1028;
input n_472;
input n_270;
input n_414;
input n_563;
input n_1011;
input n_1215;
input n_25;
input n_93;
input n_839;
input n_708;
input n_668;
input n_626;
input n_990;
input n_779;
input n_1104;
input n_854;
input n_1058;
input n_498;
input n_1122;
input n_870;
input n_904;
input n_1253;
input n_709;
input n_1266;
input n_366;
input n_103;
input n_1109;
input n_185;
input n_712;
input n_348;
input n_1276;
input n_376;
input n_390;
input n_1148;
input n_31;
input n_334;
input n_1161;
input n_1085;
input n_232;
input n_46;
input n_1239;
input n_771;
input n_470;
input n_475;
input n_924;
input n_298;
input n_492;
input n_1149;
input n_265;
input n_1184;
input n_228;
input n_719;
input n_455;
input n_363;
input n_1090;
input n_592;
input n_829;
input n_1156;
input n_1362;
input n_393;
input n_984;
input n_503;
input n_132;
input n_868;
input n_570;
input n_859;
input n_406;
input n_735;
input n_878;
input n_620;
input n_130;
input n_519;
input n_307;
input n_469;
input n_1218;
input n_500;
input n_981;
input n_714;
input n_1349;
input n_291;
input n_1144;
input n_357;
input n_985;
input n_481;
input n_997;
input n_1301;
input n_802;
input n_561;
input n_33;
input n_980;
input n_1306;
input n_1198;
input n_436;
input n_116;
input n_409;
input n_1244;
input n_240;
input n_756;
input n_810;
input n_1133;
input n_635;
input n_95;
input n_1194;
input n_1051;
input n_253;
input n_583;
input n_249;
input n_201;
input n_1039;
input n_1034;
input n_1158;
input n_754;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_1305;
input n_553;
input n_43;
input n_849;
input n_753;
input n_467;
input n_269;
input n_359;
input n_973;
input n_1055;
input n_582;
input n_861;
input n_857;
input n_967;
input n_571;
input n_271;
input n_404;
input n_158;
input n_206;
input n_679;
input n_633;
input n_1170;
input n_665;
input n_588;
input n_225;
input n_1260;
input n_308;
input n_309;
input n_1010;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_1166;
input n_812;
input n_1131;
input n_534;
input n_1006;
input n_373;
input n_87;
input n_257;
input n_730;
input n_1311;
input n_670;
input n_203;
input n_207;
input n_1089;
input n_1365;
input n_205;
input n_1242;
input n_681;
input n_1226;
input n_1274;
input n_412;
input n_640;
input n_1322;
input n_81;
input n_965;
input n_339;
input n_784;
input n_315;
input n_434;
input n_64;
input n_288;
input n_1059;
input n_1197;
input n_422;
input n_722;
input n_862;
input n_135;
input n_165;
input n_540;
input n_457;
input n_364;
input n_629;
input n_900;
input n_531;
input n_827;
input n_60;
input n_361;
input n_1025;
input n_336;
input n_12;
input n_1013;
input n_1259;
input n_192;
input n_51;
input n_649;
input n_1240;

output n_4303;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1674;
wire n_3392;
wire n_3266;
wire n_3574;
wire n_3152;
wire n_4154;
wire n_3579;
wire n_4251;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_3783;
wire n_4177;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1581;
wire n_3844;
wire n_2534;
wire n_2353;
wire n_3301;
wire n_3089;
wire n_4099;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4168;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_3911;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_2647;
wire n_2997;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_4092;
wire n_1724;
wire n_3708;
wire n_2336;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4087;
wire n_1700;
wire n_2211;
wire n_1415;
wire n_1555;
wire n_1786;
wire n_3487;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_2291;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_2886;
wire n_2974;
wire n_3946;
wire n_1985;
wire n_4213;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1867;
wire n_1517;
wire n_2926;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_3106;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_2356;
wire n_1511;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1572;
wire n_1874;
wire n_3165;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2510;
wire n_2739;
wire n_1735;
wire n_1954;
wire n_1541;
wire n_2480;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_2791;
wire n_3750;
wire n_3607;
wire n_3251;
wire n_3877;
wire n_3316;
wire n_2212;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_2729;
wire n_3063;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_4187;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1471;
wire n_3737;
wire n_3624;
wire n_3077;
wire n_3979;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_1404;
wire n_2124;
wire n_2378;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_3765;
wire n_2655;
wire n_4125;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_4262;
wire n_1894;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_4071;
wire n_4255;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_3413;
wire n_3850;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_3943;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4102;
wire n_4297;
wire n_2113;
wire n_1641;
wire n_2190;
wire n_1918;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_3959;
wire n_2268;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_1441;
wire n_3373;
wire n_2104;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_3910;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4296;
wire n_2633;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_3949;
wire n_2792;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_1530;
wire n_3798;
wire n_3488;
wire n_1543;
wire n_2811;
wire n_1599;
wire n_3732;
wire n_4257;
wire n_2674;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_3980;
wire n_2831;
wire n_2998;
wire n_3446;
wire n_4158;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_4259;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_2692;
wire n_3842;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_3099;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_3888;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4161;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_3403;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_3092;
wire n_2714;
wire n_2245;
wire n_3055;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_2068;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3734;
wire n_3686;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_3746;
wire n_1713;
wire n_2971;
wire n_3599;
wire n_2678;
wire n_3384;
wire n_3935;
wire n_4277;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_3012;
wire n_1662;
wire n_3772;
wire n_3875;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_3247;
wire n_3069;
wire n_3921;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_2664;
wire n_2641;
wire n_1722;
wire n_1664;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_3933;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_3273;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_3691;
wire n_3861;
wire n_2624;
wire n_4066;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_2347;
wire n_1801;
wire n_1886;
wire n_3917;
wire n_2092;
wire n_1654;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3428;
wire n_3153;
wire n_3410;
wire n_3689;
wire n_1752;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_4043;
wire n_2916;
wire n_3415;
wire n_4292;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_3434;
wire n_1515;
wire n_3510;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_4169;
wire n_4055;
wire n_2377;
wire n_3271;
wire n_2178;
wire n_4248;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_1630;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_3578;
wire n_3885;
wire n_2271;
wire n_3192;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_2794;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_3073;
wire n_2431;
wire n_4018;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_3253;
wire n_3337;
wire n_3431;
wire n_3450;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_4002;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2893;
wire n_2775;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_4289;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4288;
wire n_2712;
wire n_2684;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_3953;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_2913;
wire n_3614;
wire n_1756;
wire n_3183;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_1952;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_1932;
wire n_2535;
wire n_1880;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_4191;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_2870;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_2767;
wire n_3793;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_1514;
wire n_1863;
wire n_3385;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1714;
wire n_3922;
wire n_3179;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_4000;
wire n_2897;
wire n_2537;
wire n_3970;
wire n_2554;
wire n_2089;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_3171;
wire n_1913;
wire n_4216;
wire n_3608;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_2339;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3426;
wire n_3158;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2643;
wire n_2590;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_3435;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_1432;
wire n_2208;
wire n_2604;
wire n_2407;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_2012;
wire n_3497;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_2134;
wire n_2335;
wire n_1529;
wire n_2473;
wire n_3887;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_4096;
wire n_1431;
wire n_4123;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_4286;
wire n_1809;
wire n_3119;
wire n_4280;
wire n_2958;
wire n_1577;
wire n_2948;
wire n_3735;
wire n_2297;
wire n_2119;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_4218;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_3832;
wire n_2520;
wire n_4264;
wire n_2857;
wire n_3693;
wire n_3788;
wire n_2372;
wire n_1490;
wire n_1568;
wire n_2896;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_4175;
wire n_3200;
wire n_1665;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3867;
wire n_3341;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_2482;
wire n_1507;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1811;
wire n_3661;
wire n_3006;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_2424;
wire n_1604;
wire n_2296;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_3971;
wire n_2849;
wire n_1774;
wire n_1475;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_3393;
wire n_2442;
wire n_3627;
wire n_3451;
wire n_1791;
wire n_3480;
wire n_1418;
wire n_3331;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_2545;
wire n_3577;
wire n_3540;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_3606;
wire n_3142;
wire n_3598;
wire n_2966;
wire n_2294;
wire n_2581;
wire n_3641;
wire n_1966;
wire n_1942;
wire n_3591;
wire n_3777;
wire n_2218;
wire n_1837;
wire n_2788;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1534;
wire n_3892;
wire n_1564;
wire n_1736;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_3944;
wire n_3909;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_3270;
wire n_2618;
wire n_2357;
wire n_2025;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_3755;
wire n_4042;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_3481;
wire n_2329;
wire n_2237;
wire n_3026;
wire n_2250;
wire n_1951;
wire n_3090;
wire n_4299;
wire n_3033;
wire n_3724;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_3913;
wire n_4276;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3323;
wire n_3226;
wire n_3364;
wire n_4020;
wire n_4176;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_1618;
wire n_3407;
wire n_1531;
wire n_2828;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_4261;
wire n_1745;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_2920;
wire n_4015;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_3742;
wire n_2462;
wire n_1933;
wire n_3243;
wire n_2889;
wire n_3683;
wire n_4034;
wire n_4056;
wire n_1617;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_3736;
wire n_2732;
wire n_2928;
wire n_4206;
wire n_2249;
wire n_1917;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_1881;
wire n_1806;
wire n_3284;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_2289;
wire n_2315;
wire n_1733;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_3663;
wire n_4132;
wire n_2995;
wire n_2955;
wire n_1731;
wire n_2158;
wire n_3360;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4001;
wire n_1687;
wire n_2328;
wire n_1439;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_4149;
wire n_2627;
wire n_2276;
wire n_3234;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_3016;
wire n_1668;
wire n_2777;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4030;
wire n_4003;
wire n_3870;
wire n_4126;
wire n_1696;
wire n_2829;
wire n_2181;
wire n_1594;
wire n_1995;
wire n_3751;
wire n_1869;
wire n_3625;
wire n_2911;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_2448;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_2327;
wire n_2201;
wire n_3919;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_2984;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_2983;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3276;
wire n_1934;
wire n_3250;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_1728;
wire n_3973;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_3886;
wire n_2924;
wire n_3595;
wire n_3414;
wire n_1661;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_2549;
wire n_4234;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_4211;
wire n_4182;
wire n_1667;
wire n_3230;
wire n_4016;
wire n_3236;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_1409;
wire n_4230;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_4274;
wire n_2423;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4270;
wire n_4151;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_3730;
wire n_2404;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_4155;
wire n_2740;
wire n_4238;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_3042;
wire n_1589;
wire n_3213;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1943;
wire n_3228;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_2472;
wire n_3238;
wire n_1891;
wire n_2171;
wire n_3529;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4109;
wire n_4192;
wire n_1443;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_2808;
wire n_2037;
wire n_3710;
wire n_4159;
wire n_4195;
wire n_3784;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_2373;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_3628;
wire n_4144;
wire n_1870;
wire n_2964;
wire n_4174;
wire n_1692;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3475;
wire n_3501;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1642;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_2257;
wire n_3692;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_4258;
wire n_3597;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_2670;
wire n_2700;
wire n_2346;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_3045;
wire n_3821;
wire n_3115;
wire n_1883;
wire n_4300;
wire n_3318;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_3439;
wire n_3588;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_4135;
wire n_4209;
wire n_2871;
wire n_4279;
wire n_2688;
wire n_1456;
wire n_1845;
wire n_3858;
wire n_4183;
wire n_1489;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_1544;
wire n_2258;
wire n_1485;
wire n_1640;
wire n_4040;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_2390;
wire n_4007;
wire n_3712;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1522;
wire n_4239;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_3562;
wire n_3044;
wire n_2973;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_2154;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1672;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1914;
wire n_3457;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_3762;
wire n_3932;
wire n_3469;
wire n_3958;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1556;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_3713;
wire n_3379;
wire n_3156;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_1650;
wire n_1794;
wire n_1962;
wire n_3506;
wire n_2398;
wire n_1559;
wire n_1928;
wire n_1725;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_3124;
wire n_1741;
wire n_1746;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_3524;
wire n_2671;
wire n_2761;
wire n_2888;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_2885;
wire n_3711;
wire n_3776;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_2070;
wire n_2588;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_3308;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_3694;
wire n_2937;
wire n_2045;
wire n_2261;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_1800;
wire n_2241;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_4203;
wire n_3808;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1826;
wire n_1882;
wire n_2951;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_3758;
wire n_1879;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_3585;
wire n_3565;
wire n_1953;
wire n_3343;
wire n_3303;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_1976;
wire n_4229;
wire n_2905;
wire n_3990;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_3890;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_2358;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_3951;
wire n_3034;
wire n_3569;
wire n_3874;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_3027;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_4295;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_2020;
wire n_1643;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_3117;
wire n_1461;
wire n_3432;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_3774;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_2910;
wire n_2385;
wire n_4112;
wire n_1848;
wire n_1785;
wire n_3268;
wire n_4009;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_3473;
wire n_2485;
wire n_2450;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_2769;
wire n_3622;
wire n_2492;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1570;
wire n_1702;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_2180;
wire n_1689;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_3573;
wire n_1944;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_3334;
wire n_4027;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_3553;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_2275;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_3811;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_2255;
wire n_2112;
wire n_3494;
wire n_1464;
wire n_2430;
wire n_1737;
wire n_3486;
wire n_1414;
wire n_4086;
wire n_2649;
wire n_2721;
wire n_3556;
wire n_2034;
wire n_3836;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_4068;
wire n_2032;
wire n_2744;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_4166;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_3404;
wire n_3745;
wire n_3362;
wire n_2242;
wire n_4059;
wire n_1509;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_3523;
wire n_2222;
wire n_3256;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4142;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_2505;
wire n_2188;
wire n_2609;
wire n_1989;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_3643;
wire n_3697;
wire n_1584;
wire n_2425;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_2666;
wire n_4105;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_2147;
wire n_2564;
wire n_4244;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_3123;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_3038;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_2531;
wire n_1789;
wire n_1770;
wire n_3285;
wire n_4208;
wire n_2523;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_3596;
wire n_3478;
wire n_3936;
wire n_4089;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3521;
wire n_3233;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_2805;
wire n_3310;
wire n_2681;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_3989;
wire n_2478;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_4108;
wire n_3374;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_4051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_2909;
wire n_2248;
wire n_4293;
wire n_3552;
wire n_3206;
wire n_2363;
wire n_2578;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_3709;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_3187;
wire n_2540;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_2217;
wire n_1675;
wire n_2197;
wire n_2065;
wire n_2879;
wire n_3717;
wire n_4148;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_4057;
wire n_2968;
wire n_4201;
wire n_1629;
wire n_2221;
wire n_4263;
wire n_2055;
wire n_1819;
wire n_3555;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_3059;
wire n_2038;
wire n_2891;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_1578;
wire n_1861;
wire n_3110;
wire n_1890;
wire n_1632;
wire n_3017;
wire n_3955;
wire n_2477;
wire n_1805;
wire n_1888;
wire n_2280;
wire n_1557;
wire n_1833;
wire n_3903;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_2333;
wire n_1868;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_4138;
wire n_1417;
wire n_2185;
wire n_2086;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_3740;
wire n_3162;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3333;
wire n_3274;
wire n_3186;
wire n_4129;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3584;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_4275;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_2912;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_3182;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;

INVx1_ASAP7_75t_L g1402 ( 
.A(n_909),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_837),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_989),
.Y(n_1404)
);

BUFx10_ASAP7_75t_L g1405 ( 
.A(n_999),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_752),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1346),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1076),
.Y(n_1408)
);

CKINVDCx16_ASAP7_75t_R g1409 ( 
.A(n_288),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_138),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1291),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_846),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1146),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_128),
.Y(n_1414)
);

INVx2_ASAP7_75t_SL g1415 ( 
.A(n_537),
.Y(n_1415)
);

CKINVDCx20_ASAP7_75t_R g1416 ( 
.A(n_1126),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_887),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_720),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1318),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_250),
.Y(n_1420)
);

INVxp67_ASAP7_75t_SL g1421 ( 
.A(n_1273),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_462),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1166),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_7),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_242),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1105),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1312),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_706),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_138),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_247),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1303),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1324),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_502),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1270),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1264),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_781),
.Y(n_1436)
);

INVx2_ASAP7_75t_SL g1437 ( 
.A(n_1396),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1326),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1087),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1240),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_668),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_368),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1039),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_571),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_307),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1313),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_849),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_15),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1342),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1309),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_308),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_574),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1348),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1102),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_670),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_787),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1308),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_604),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_145),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_311),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_476),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1279),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_511),
.Y(n_1463)
);

INVxp33_ASAP7_75t_L g1464 ( 
.A(n_742),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1032),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_213),
.Y(n_1466)
);

CKINVDCx20_ASAP7_75t_R g1467 ( 
.A(n_943),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_754),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_505),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_797),
.Y(n_1470)
);

BUFx10_ASAP7_75t_L g1471 ( 
.A(n_1003),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_736),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_654),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_497),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_697),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_648),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_948),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_185),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_393),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_564),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1361),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1144),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1352),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_869),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_618),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_527),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1335),
.Y(n_1487)
);

CKINVDCx16_ASAP7_75t_R g1488 ( 
.A(n_970),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_510),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_36),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1276),
.Y(n_1491)
);

BUFx8_ASAP7_75t_SL g1492 ( 
.A(n_998),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_372),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_382),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_539),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1142),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1379),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_520),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_444),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_822),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1388),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_726),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_528),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1038),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_533),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_791),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1248),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_924),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_550),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_426),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_1086),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_297),
.Y(n_1512)
);

INVx1_ASAP7_75t_SL g1513 ( 
.A(n_1269),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_181),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_1054),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_496),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_503),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_997),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_320),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1400),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1152),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_682),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_352),
.Y(n_1523)
);

INVx1_ASAP7_75t_SL g1524 ( 
.A(n_507),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_67),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1271),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1021),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1323),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1136),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_213),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1318),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_897),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_639),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1317),
.Y(n_1534)
);

CKINVDCx14_ASAP7_75t_R g1535 ( 
.A(n_834),
.Y(n_1535)
);

CKINVDCx20_ASAP7_75t_R g1536 ( 
.A(n_743),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1297),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_872),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1280),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1022),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_271),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1349),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1081),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1397),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_950),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1266),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1343),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1162),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_939),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_601),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1384),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_1322),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_866),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_365),
.Y(n_1554)
);

INVxp67_ASAP7_75t_L g1555 ( 
.A(n_698),
.Y(n_1555)
);

INVxp33_ASAP7_75t_R g1556 ( 
.A(n_657),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_865),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_309),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_946),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_260),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_58),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_240),
.Y(n_1562)
);

CKINVDCx20_ASAP7_75t_R g1563 ( 
.A(n_1319),
.Y(n_1563)
);

CKINVDCx14_ASAP7_75t_R g1564 ( 
.A(n_1344),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1282),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_925),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1058),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1257),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1361),
.Y(n_1569)
);

CKINVDCx20_ASAP7_75t_R g1570 ( 
.A(n_724),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1325),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1340),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1047),
.Y(n_1573)
);

BUFx10_ASAP7_75t_L g1574 ( 
.A(n_549),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_70),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1115),
.Y(n_1576)
);

CKINVDCx14_ASAP7_75t_R g1577 ( 
.A(n_454),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_882),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_932),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1197),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1353),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1146),
.Y(n_1582)
);

BUFx5_ASAP7_75t_L g1583 ( 
.A(n_494),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_1167),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_889),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_900),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_249),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_463),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_231),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_984),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_321),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_687),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1107),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_659),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_48),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_72),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_294),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_1020),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1307),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_391),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_158),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_297),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1395),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_295),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1071),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_359),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_780),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1210),
.Y(n_1608)
);

BUFx10_ASAP7_75t_L g1609 ( 
.A(n_1293),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_184),
.Y(n_1610)
);

CKINVDCx20_ASAP7_75t_R g1611 ( 
.A(n_796),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_806),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_888),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1334),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_183),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_103),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1217),
.Y(n_1617)
);

CKINVDCx16_ASAP7_75t_R g1618 ( 
.A(n_334),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1316),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_808),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_553),
.Y(n_1621)
);

CKINVDCx20_ASAP7_75t_R g1622 ( 
.A(n_1386),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1292),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1267),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1216),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1311),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1274),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_426),
.Y(n_1628)
);

CKINVDCx20_ASAP7_75t_R g1629 ( 
.A(n_680),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_122),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_838),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_391),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_785),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_388),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_1077),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1112),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_677),
.Y(n_1637)
);

CKINVDCx20_ASAP7_75t_R g1638 ( 
.A(n_1346),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_32),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_905),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_334),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_721),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1048),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_28),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1372),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_430),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1234),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1398),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_847),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_583),
.Y(n_1650)
);

CKINVDCx20_ASAP7_75t_R g1651 ( 
.A(n_1333),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1088),
.Y(n_1652)
);

CKINVDCx20_ASAP7_75t_R g1653 ( 
.A(n_365),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_275),
.Y(n_1654)
);

CKINVDCx20_ASAP7_75t_R g1655 ( 
.A(n_493),
.Y(n_1655)
);

BUFx10_ASAP7_75t_L g1656 ( 
.A(n_1265),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_121),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_146),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_551),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1313),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_87),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1109),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1128),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1290),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1298),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_491),
.Y(n_1666)
);

BUFx10_ASAP7_75t_L g1667 ( 
.A(n_861),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_985),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1258),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_486),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1027),
.Y(n_1671)
);

CKINVDCx20_ASAP7_75t_R g1672 ( 
.A(n_123),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1028),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1046),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_461),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1068),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_987),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_6),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_922),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_3),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1043),
.Y(n_1681)
);

BUFx2_ASAP7_75t_SL g1682 ( 
.A(n_1193),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_81),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_783),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_784),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_245),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1357),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_248),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1030),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_696),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_838),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_383),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_546),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_643),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_129),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_173),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1031),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_13),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1284),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1161),
.Y(n_1700)
);

CKINVDCx20_ASAP7_75t_R g1701 ( 
.A(n_389),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1156),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1399),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1039),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1239),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_867),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_16),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_168),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_1302),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1299),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_732),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_332),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1347),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1350),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1330),
.Y(n_1715)
);

CKINVDCx20_ASAP7_75t_R g1716 ( 
.A(n_974),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1336),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_1393),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1277),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1278),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_479),
.Y(n_1721)
);

BUFx2_ASAP7_75t_L g1722 ( 
.A(n_855),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1145),
.Y(n_1723)
);

CKINVDCx20_ASAP7_75t_R g1724 ( 
.A(n_818),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_940),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_740),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_668),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_576),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_546),
.Y(n_1729)
);

CKINVDCx20_ASAP7_75t_R g1730 ( 
.A(n_1331),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_968),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_674),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_850),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_585),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1148),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1053),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1343),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_170),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1294),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_807),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1055),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_471),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_651),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_930),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_997),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_516),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1072),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_594),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_969),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_240),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_835),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_635),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_290),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1208),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_896),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1121),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1286),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_596),
.Y(n_1758)
);

CKINVDCx14_ASAP7_75t_R g1759 ( 
.A(n_828),
.Y(n_1759)
);

CKINVDCx20_ASAP7_75t_R g1760 ( 
.A(n_868),
.Y(n_1760)
);

BUFx10_ASAP7_75t_L g1761 ( 
.A(n_588),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_1085),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1272),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_88),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_1392),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_113),
.Y(n_1766)
);

INVxp67_ASAP7_75t_SL g1767 ( 
.A(n_1277),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_420),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_314),
.Y(n_1769)
);

CKINVDCx20_ASAP7_75t_R g1770 ( 
.A(n_462),
.Y(n_1770)
);

BUFx6f_ASAP7_75t_L g1771 ( 
.A(n_545),
.Y(n_1771)
);

BUFx2_ASAP7_75t_L g1772 ( 
.A(n_257),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1315),
.Y(n_1773)
);

BUFx10_ASAP7_75t_L g1774 ( 
.A(n_82),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_1055),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1196),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_338),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_403),
.Y(n_1778)
);

BUFx6f_ASAP7_75t_L g1779 ( 
.A(n_451),
.Y(n_1779)
);

CKINVDCx20_ASAP7_75t_R g1780 ( 
.A(n_1370),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_1263),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1338),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_133),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_700),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1268),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_89),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_715),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1349),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_513),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_631),
.Y(n_1790)
);

CKINVDCx20_ASAP7_75t_R g1791 ( 
.A(n_1063),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_744),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_729),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1165),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_1243),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1027),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1045),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_548),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1119),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1295),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1329),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_417),
.Y(n_1802)
);

CKINVDCx14_ASAP7_75t_R g1803 ( 
.A(n_770),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_1351),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1209),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_692),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_1341),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1052),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_429),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_786),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_50),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_88),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_636),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1306),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_1358),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_282),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1304),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1195),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_827),
.Y(n_1819)
);

CKINVDCx16_ASAP7_75t_R g1820 ( 
.A(n_474),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_559),
.Y(n_1821)
);

BUFx3_ASAP7_75t_L g1822 ( 
.A(n_213),
.Y(n_1822)
);

CKINVDCx20_ASAP7_75t_R g1823 ( 
.A(n_177),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_595),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_1241),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_1222),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1371),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_647),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1292),
.Y(n_1829)
);

CKINVDCx16_ASAP7_75t_R g1830 ( 
.A(n_12),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_653),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_662),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_430),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_456),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1090),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_195),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_385),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_286),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_594),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_171),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_347),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_224),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1317),
.Y(n_1843)
);

CKINVDCx14_ASAP7_75t_R g1844 ( 
.A(n_780),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_530),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_309),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_187),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_61),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_1309),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_1310),
.Y(n_1850)
);

BUFx10_ASAP7_75t_L g1851 ( 
.A(n_893),
.Y(n_1851)
);

CKINVDCx20_ASAP7_75t_R g1852 ( 
.A(n_318),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1394),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_449),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_965),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1074),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_57),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_371),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1192),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_538),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_28),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_629),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_788),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_335),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_978),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1005),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_271),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_1260),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1211),
.Y(n_1869)
);

BUFx3_ASAP7_75t_L g1870 ( 
.A(n_1324),
.Y(n_1870)
);

BUFx2_ASAP7_75t_L g1871 ( 
.A(n_1331),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_71),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_602),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_533),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_907),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_859),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_90),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_577),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_162),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_568),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1296),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_257),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_914),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_448),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1314),
.Y(n_1885)
);

CKINVDCx20_ASAP7_75t_R g1886 ( 
.A(n_627),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_28),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_234),
.Y(n_1888)
);

BUFx2_ASAP7_75t_L g1889 ( 
.A(n_90),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_274),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1227),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_1327),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_1355),
.Y(n_1893)
);

CKINVDCx20_ASAP7_75t_R g1894 ( 
.A(n_545),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_188),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_821),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_833),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1259),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1149),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_842),
.Y(n_1900)
);

CKINVDCx20_ASAP7_75t_R g1901 ( 
.A(n_283),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_688),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_1212),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_11),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1320),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1332),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_190),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_562),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1169),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_962),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_901),
.Y(n_1911)
);

CKINVDCx20_ASAP7_75t_R g1912 ( 
.A(n_582),
.Y(n_1912)
);

BUFx8_ASAP7_75t_SL g1913 ( 
.A(n_182),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1294),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_856),
.Y(n_1915)
);

CKINVDCx20_ASAP7_75t_R g1916 ( 
.A(n_817),
.Y(n_1916)
);

HB1xp67_ASAP7_75t_L g1917 ( 
.A(n_794),
.Y(n_1917)
);

CKINVDCx20_ASAP7_75t_R g1918 ( 
.A(n_540),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_481),
.Y(n_1919)
);

BUFx10_ASAP7_75t_L g1920 ( 
.A(n_682),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_326),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_1203),
.Y(n_1922)
);

INVx3_ASAP7_75t_L g1923 ( 
.A(n_614),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_992),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_315),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_1275),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_177),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1164),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1062),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_877),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_42),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_489),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_341),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_1200),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_1139),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_501),
.Y(n_1936)
);

BUFx6f_ASAP7_75t_L g1937 ( 
.A(n_761),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_827),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_1328),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_917),
.Y(n_1940)
);

CKINVDCx5p33_ASAP7_75t_R g1941 ( 
.A(n_714),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1168),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1069),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_1285),
.Y(n_1944)
);

BUFx6f_ASAP7_75t_L g1945 ( 
.A(n_1101),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1301),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_945),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1339),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_1315),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1269),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_821),
.Y(n_1951)
);

CKINVDCx20_ASAP7_75t_R g1952 ( 
.A(n_1229),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_890),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_795),
.Y(n_1954)
);

BUFx6f_ASAP7_75t_L g1955 ( 
.A(n_1262),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_83),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_974),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1111),
.Y(n_1958)
);

BUFx2_ASAP7_75t_SL g1959 ( 
.A(n_1283),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_844),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1321),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_959),
.Y(n_1962)
);

BUFx2_ASAP7_75t_SL g1963 ( 
.A(n_1163),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_277),
.Y(n_1964)
);

CKINVDCx5p33_ASAP7_75t_R g1965 ( 
.A(n_440),
.Y(n_1965)
);

CKINVDCx5p33_ASAP7_75t_R g1966 ( 
.A(n_35),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_186),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1004),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1001),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_938),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_337),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_1161),
.Y(n_1972)
);

BUFx10_ASAP7_75t_L g1973 ( 
.A(n_1116),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1356),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_900),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_915),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_100),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1221),
.Y(n_1978)
);

CKINVDCx20_ASAP7_75t_R g1979 ( 
.A(n_347),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_150),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_423),
.Y(n_1981)
);

BUFx6f_ASAP7_75t_L g1982 ( 
.A(n_1219),
.Y(n_1982)
);

INVx1_ASAP7_75t_SL g1983 ( 
.A(n_870),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1305),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_1042),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_375),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_566),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1288),
.Y(n_1988)
);

CKINVDCx5p33_ASAP7_75t_R g1989 ( 
.A(n_683),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_531),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_857),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1051),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_575),
.Y(n_1993)
);

BUFx8_ASAP7_75t_SL g1994 ( 
.A(n_1345),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1374),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_531),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_705),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_159),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_976),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_13),
.Y(n_2000)
);

INVx1_ASAP7_75t_SL g2001 ( 
.A(n_115),
.Y(n_2001)
);

BUFx3_ASAP7_75t_L g2002 ( 
.A(n_893),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1026),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_1100),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_820),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_650),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1337),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1131),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1359),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1009),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_1383),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_128),
.Y(n_2012)
);

INVx1_ASAP7_75t_SL g2013 ( 
.A(n_216),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_447),
.Y(n_2014)
);

CKINVDCx16_ASAP7_75t_R g2015 ( 
.A(n_921),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1341),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_429),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_798),
.Y(n_2018)
);

BUFx3_ASAP7_75t_L g2019 ( 
.A(n_1261),
.Y(n_2019)
);

CKINVDCx5p33_ASAP7_75t_R g2020 ( 
.A(n_318),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_1070),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_1281),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_1289),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_716),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_1300),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_167),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_731),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_577),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_685),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1354),
.Y(n_2030)
);

INVx1_ASAP7_75t_SL g2031 ( 
.A(n_210),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_313),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_461),
.Y(n_2033)
);

BUFx3_ASAP7_75t_L g2034 ( 
.A(n_789),
.Y(n_2034)
);

BUFx2_ASAP7_75t_L g2035 ( 
.A(n_279),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_635),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1265),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1094),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1360),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1091),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_477),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1006),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_440),
.Y(n_2043)
);

CKINVDCx5p33_ASAP7_75t_R g2044 ( 
.A(n_1390),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_639),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1366),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1131),
.Y(n_2047)
);

BUFx2_ASAP7_75t_L g2048 ( 
.A(n_704),
.Y(n_2048)
);

CKINVDCx20_ASAP7_75t_R g2049 ( 
.A(n_328),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_762),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_1100),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_1287),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_1375),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_584),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_397),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_362),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_730),
.Y(n_2057)
);

CKINVDCx16_ASAP7_75t_R g2058 ( 
.A(n_1409),
.Y(n_2058)
);

INVxp33_ASAP7_75t_SL g2059 ( 
.A(n_1693),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1583),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_L g2061 ( 
.A(n_1535),
.B(n_0),
.Y(n_2061)
);

CKINVDCx20_ASAP7_75t_R g2062 ( 
.A(n_1564),
.Y(n_2062)
);

BUFx3_ASAP7_75t_L g2063 ( 
.A(n_1558),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1583),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1583),
.Y(n_2065)
);

HB1xp67_ASAP7_75t_L g2066 ( 
.A(n_1913),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1583),
.Y(n_2067)
);

CKINVDCx20_ASAP7_75t_R g2068 ( 
.A(n_1577),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1583),
.Y(n_2069)
);

BUFx2_ASAP7_75t_L g2070 ( 
.A(n_1492),
.Y(n_2070)
);

CKINVDCx16_ASAP7_75t_R g2071 ( 
.A(n_1830),
.Y(n_2071)
);

INVxp67_ASAP7_75t_L g2072 ( 
.A(n_1772),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1445),
.Y(n_2073)
);

INVx1_ASAP7_75t_SL g2074 ( 
.A(n_1889),
.Y(n_2074)
);

CKINVDCx20_ASAP7_75t_R g2075 ( 
.A(n_1759),
.Y(n_2075)
);

CKINVDCx20_ASAP7_75t_R g2076 ( 
.A(n_1803),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1448),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1478),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_1994),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1519),
.Y(n_2080)
);

CKINVDCx20_ASAP7_75t_R g2081 ( 
.A(n_1844),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1530),
.Y(n_2082)
);

INVxp33_ASAP7_75t_L g2083 ( 
.A(n_2035),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1575),
.Y(n_2084)
);

BUFx2_ASAP7_75t_L g2085 ( 
.A(n_1501),
.Y(n_2085)
);

CKINVDCx20_ASAP7_75t_R g2086 ( 
.A(n_1488),
.Y(n_2086)
);

CKINVDCx20_ASAP7_75t_R g2087 ( 
.A(n_1618),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1595),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1596),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1602),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1610),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1630),
.Y(n_2092)
);

INVx1_ASAP7_75t_SL g2093 ( 
.A(n_1502),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1639),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1644),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1661),
.Y(n_2096)
);

INVxp33_ASAP7_75t_SL g2097 ( 
.A(n_1699),
.Y(n_2097)
);

INVxp67_ASAP7_75t_SL g2098 ( 
.A(n_1809),
.Y(n_2098)
);

BUFx6f_ASAP7_75t_L g2099 ( 
.A(n_1683),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1678),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1686),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1695),
.Y(n_2102)
);

CKINVDCx5p33_ASAP7_75t_R g2103 ( 
.A(n_1820),
.Y(n_2103)
);

BUFx2_ASAP7_75t_L g2104 ( 
.A(n_1636),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1786),
.Y(n_2105)
);

CKINVDCx20_ASAP7_75t_R g2106 ( 
.A(n_2015),
.Y(n_2106)
);

BUFx5_ASAP7_75t_L g2107 ( 
.A(n_1402),
.Y(n_2107)
);

BUFx3_ASAP7_75t_L g2108 ( 
.A(n_1822),
.Y(n_2108)
);

CKINVDCx14_ASAP7_75t_R g2109 ( 
.A(n_1714),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1840),
.Y(n_2110)
);

HB1xp67_ASAP7_75t_L g2111 ( 
.A(n_1810),
.Y(n_2111)
);

CKINVDCx5p33_ASAP7_75t_R g2112 ( 
.A(n_1410),
.Y(n_2112)
);

CKINVDCx20_ASAP7_75t_R g2113 ( 
.A(n_1403),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1847),
.Y(n_2114)
);

INVxp67_ASAP7_75t_SL g2115 ( 
.A(n_1809),
.Y(n_2115)
);

NOR2xp67_ASAP7_75t_L g2116 ( 
.A(n_1923),
.B(n_0),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1867),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1877),
.Y(n_2118)
);

INVxp33_ASAP7_75t_SL g2119 ( 
.A(n_1917),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1888),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1895),
.Y(n_2121)
);

INVxp33_ASAP7_75t_SL g2122 ( 
.A(n_1943),
.Y(n_2122)
);

CKINVDCx20_ASAP7_75t_R g2123 ( 
.A(n_1416),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1907),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_1414),
.Y(n_2125)
);

CKINVDCx20_ASAP7_75t_R g2126 ( 
.A(n_1431),
.Y(n_2126)
);

BUFx2_ASAP7_75t_L g2127 ( 
.A(n_1722),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1931),
.Y(n_2128)
);

INVxp33_ASAP7_75t_L g2129 ( 
.A(n_1871),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1964),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1977),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1980),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1998),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_1420),
.Y(n_2134)
);

CKINVDCx20_ASAP7_75t_R g2135 ( 
.A(n_1467),
.Y(n_2135)
);

INVxp67_ASAP7_75t_SL g2136 ( 
.A(n_1683),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1430),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1783),
.Y(n_2138)
);

INVx3_ASAP7_75t_L g2139 ( 
.A(n_1569),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1783),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1783),
.Y(n_2141)
);

CKINVDCx5p33_ASAP7_75t_R g2142 ( 
.A(n_1424),
.Y(n_2142)
);

CKINVDCx20_ASAP7_75t_R g2143 ( 
.A(n_1515),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2012),
.Y(n_2144)
);

CKINVDCx5p33_ASAP7_75t_R g2145 ( 
.A(n_1425),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2012),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1459),
.Y(n_2147)
);

INVxp67_ASAP7_75t_SL g2148 ( 
.A(n_1569),
.Y(n_2148)
);

BUFx3_ASAP7_75t_L g2149 ( 
.A(n_1456),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1460),
.Y(n_2150)
);

CKINVDCx14_ASAP7_75t_R g2151 ( 
.A(n_2048),
.Y(n_2151)
);

CKINVDCx5p33_ASAP7_75t_R g2152 ( 
.A(n_1429),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1466),
.Y(n_2153)
);

INVxp67_ASAP7_75t_L g2154 ( 
.A(n_1774),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1490),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1512),
.Y(n_2156)
);

CKINVDCx14_ASAP7_75t_R g2157 ( 
.A(n_1405),
.Y(n_2157)
);

INVxp67_ASAP7_75t_SL g2158 ( 
.A(n_1569),
.Y(n_2158)
);

HB1xp67_ASAP7_75t_L g2159 ( 
.A(n_1451),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1698),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1708),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1836),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2032),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1614),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1614),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1614),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1674),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1771),
.Y(n_2168)
);

CKINVDCx20_ASAP7_75t_R g2169 ( 
.A(n_1536),
.Y(n_2169)
);

CKINVDCx20_ASAP7_75t_R g2170 ( 
.A(n_1563),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1779),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1824),
.Y(n_2172)
);

HB1xp67_ASAP7_75t_L g2173 ( 
.A(n_1514),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1824),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1937),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1937),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1937),
.Y(n_2177)
);

CKINVDCx5p33_ASAP7_75t_R g2178 ( 
.A(n_1525),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1945),
.Y(n_2179)
);

CKINVDCx16_ASAP7_75t_R g2180 ( 
.A(n_1471),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1945),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_1541),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1955),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1955),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1982),
.Y(n_2185)
);

BUFx6f_ASAP7_75t_L g2186 ( 
.A(n_1982),
.Y(n_2186)
);

CKINVDCx16_ASAP7_75t_R g2187 ( 
.A(n_1471),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1517),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1551),
.Y(n_2189)
);

CKINVDCx5p33_ASAP7_75t_R g2190 ( 
.A(n_1560),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1647),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1650),
.Y(n_2192)
);

CKINVDCx16_ASAP7_75t_R g2193 ( 
.A(n_1574),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1705),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_1561),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1870),
.Y(n_2196)
);

CKINVDCx20_ASAP7_75t_R g2197 ( 
.A(n_1570),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2002),
.Y(n_2198)
);

CKINVDCx5p33_ASAP7_75t_R g2199 ( 
.A(n_1562),
.Y(n_2199)
);

CKINVDCx20_ASAP7_75t_R g2200 ( 
.A(n_1592),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2019),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2034),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2054),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2055),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2057),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1406),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1407),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1412),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1413),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1417),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1418),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1426),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1434),
.Y(n_2213)
);

CKINVDCx5p33_ASAP7_75t_R g2214 ( 
.A(n_1587),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1438),
.Y(n_2215)
);

INVxp33_ASAP7_75t_L g2216 ( 
.A(n_1464),
.Y(n_2216)
);

CKINVDCx5p33_ASAP7_75t_R g2217 ( 
.A(n_1589),
.Y(n_2217)
);

INVxp33_ASAP7_75t_L g2218 ( 
.A(n_1440),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1441),
.Y(n_2219)
);

INVxp67_ASAP7_75t_SL g2220 ( 
.A(n_1696),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1449),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1452),
.Y(n_2222)
);

BUFx6f_ASAP7_75t_L g2223 ( 
.A(n_2099),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2165),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2148),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2098),
.B(n_1415),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2158),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2115),
.B(n_1419),
.Y(n_2228)
);

AOI22xp5_ASAP7_75t_L g2229 ( 
.A1(n_2059),
.A2(n_1591),
.B1(n_1601),
.B2(n_1597),
.Y(n_2229)
);

BUFx6f_ASAP7_75t_L g2230 ( 
.A(n_2099),
.Y(n_2230)
);

AOI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2097),
.A2(n_1604),
.B1(n_1616),
.B2(n_1615),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2136),
.Y(n_2232)
);

AND2x2_ASAP7_75t_SL g2233 ( 
.A(n_2058),
.B(n_1447),
.Y(n_2233)
);

BUFx3_ASAP7_75t_L g2234 ( 
.A(n_2063),
.Y(n_2234)
);

BUFx6f_ASAP7_75t_L g2235 ( 
.A(n_2099),
.Y(n_2235)
);

BUFx6f_ASAP7_75t_L g2236 ( 
.A(n_2186),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2216),
.B(n_1421),
.Y(n_2237)
);

AND2x2_ASAP7_75t_R g2238 ( 
.A(n_2086),
.B(n_1556),
.Y(n_2238)
);

INVx4_ASAP7_75t_L g2239 ( 
.A(n_2112),
.Y(n_2239)
);

BUFx12f_ASAP7_75t_L g2240 ( 
.A(n_2079),
.Y(n_2240)
);

AND2x4_ASAP7_75t_L g2241 ( 
.A(n_2072),
.B(n_1437),
.Y(n_2241)
);

OAI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_2119),
.A2(n_2122),
.B1(n_2093),
.B2(n_2109),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2186),
.Y(n_2243)
);

BUFx6f_ASAP7_75t_L g2244 ( 
.A(n_2186),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2138),
.Y(n_2245)
);

BUFx6f_ASAP7_75t_L g2246 ( 
.A(n_2139),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2140),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2141),
.Y(n_2248)
);

INVx4_ASAP7_75t_L g2249 ( 
.A(n_2125),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_2144),
.Y(n_2250)
);

OA21x2_ASAP7_75t_L g2251 ( 
.A1(n_2060),
.A2(n_1470),
.B(n_1450),
.Y(n_2251)
);

BUFx8_ASAP7_75t_L g2252 ( 
.A(n_2070),
.Y(n_2252)
);

BUFx6f_ASAP7_75t_L g2253 ( 
.A(n_2108),
.Y(n_2253)
);

CKINVDCx5p33_ASAP7_75t_R g2254 ( 
.A(n_2134),
.Y(n_2254)
);

NAND2xp33_ASAP7_75t_L g2255 ( 
.A(n_2142),
.B(n_2145),
.Y(n_2255)
);

AOI22xp5_ASAP7_75t_L g2256 ( 
.A1(n_2061),
.A2(n_1657),
.B1(n_1658),
.B2(n_1654),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2146),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2164),
.Y(n_2258)
);

INVx3_ASAP7_75t_L g2259 ( 
.A(n_2149),
.Y(n_2259)
);

BUFx8_ASAP7_75t_L g2260 ( 
.A(n_2085),
.Y(n_2260)
);

INVx4_ASAP7_75t_L g2261 ( 
.A(n_2152),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2166),
.Y(n_2262)
);

OAI22xp5_ASAP7_75t_L g2263 ( 
.A1(n_2151),
.A2(n_1688),
.B1(n_1707),
.B2(n_1680),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2167),
.Y(n_2264)
);

BUFx6f_ASAP7_75t_L g2265 ( 
.A(n_2091),
.Y(n_2265)
);

INVx6_ASAP7_75t_L g2266 ( 
.A(n_2180),
.Y(n_2266)
);

BUFx3_ASAP7_75t_L g2267 ( 
.A(n_2192),
.Y(n_2267)
);

OA21x2_ASAP7_75t_L g2268 ( 
.A1(n_2064),
.A2(n_1544),
.B(n_1477),
.Y(n_2268)
);

AOI22xp5_ASAP7_75t_L g2269 ( 
.A1(n_2103),
.A2(n_1738),
.B1(n_1753),
.B2(n_1750),
.Y(n_2269)
);

INVxp67_ASAP7_75t_L g2270 ( 
.A(n_2159),
.Y(n_2270)
);

OAI21x1_ASAP7_75t_L g2271 ( 
.A1(n_2065),
.A2(n_1578),
.B(n_1548),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_2096),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_L g2273 ( 
.A(n_2102),
.Y(n_2273)
);

AOI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_2071),
.A2(n_1764),
.B1(n_1769),
.B2(n_1766),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2168),
.Y(n_2275)
);

BUFx6f_ASAP7_75t_L g2276 ( 
.A(n_2110),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2220),
.B(n_1691),
.Y(n_2277)
);

BUFx6f_ASAP7_75t_L g2278 ( 
.A(n_2121),
.Y(n_2278)
);

INVx3_ASAP7_75t_L g2279 ( 
.A(n_2137),
.Y(n_2279)
);

OAI21x1_ASAP7_75t_L g2280 ( 
.A1(n_2067),
.A2(n_1585),
.B(n_1581),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2171),
.Y(n_2281)
);

BUFx6f_ASAP7_75t_L g2282 ( 
.A(n_2128),
.Y(n_2282)
);

BUFx3_ASAP7_75t_L g2283 ( 
.A(n_2188),
.Y(n_2283)
);

BUFx6f_ASAP7_75t_L g2284 ( 
.A(n_2156),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2173),
.B(n_1767),
.Y(n_2285)
);

OAI22xp5_ASAP7_75t_SL g2286 ( 
.A1(n_2087),
.A2(n_1823),
.B1(n_1852),
.B2(n_1672),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2172),
.Y(n_2287)
);

BUFx3_ASAP7_75t_L g2288 ( 
.A(n_2189),
.Y(n_2288)
);

BUFx3_ASAP7_75t_L g2289 ( 
.A(n_2191),
.Y(n_2289)
);

BUFx6f_ASAP7_75t_L g2290 ( 
.A(n_2174),
.Y(n_2290)
);

BUFx6f_ASAP7_75t_L g2291 ( 
.A(n_2175),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2176),
.Y(n_2292)
);

NOR2xp33_ASAP7_75t_L g2293 ( 
.A(n_2178),
.B(n_1811),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2177),
.Y(n_2294)
);

CKINVDCx16_ASAP7_75t_R g2295 ( 
.A(n_2062),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2179),
.Y(n_2296)
);

OAI21x1_ASAP7_75t_L g2297 ( 
.A1(n_2069),
.A2(n_2183),
.B(n_2181),
.Y(n_2297)
);

BUFx6f_ASAP7_75t_L g2298 ( 
.A(n_2184),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2182),
.B(n_1816),
.Y(n_2299)
);

BUFx8_ASAP7_75t_L g2300 ( 
.A(n_2104),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2185),
.Y(n_2301)
);

OAI22xp5_ASAP7_75t_L g2302 ( 
.A1(n_2074),
.A2(n_1842),
.B1(n_1846),
.B2(n_1838),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2068),
.A2(n_1857),
.B1(n_1861),
.B2(n_1848),
.Y(n_2303)
);

NOR2x1_ASAP7_75t_L g2304 ( 
.A(n_2116),
.B(n_1586),
.Y(n_2304)
);

HB1xp67_ASAP7_75t_L g2305 ( 
.A(n_2190),
.Y(n_2305)
);

AOI22xp5_ASAP7_75t_L g2306 ( 
.A1(n_2075),
.A2(n_1872),
.B1(n_1882),
.B2(n_1879),
.Y(n_2306)
);

OA21x2_ASAP7_75t_L g2307 ( 
.A1(n_2203),
.A2(n_1608),
.B(n_1603),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2204),
.Y(n_2308)
);

OA21x2_ASAP7_75t_L g2309 ( 
.A1(n_2205),
.A2(n_2207),
.B(n_2206),
.Y(n_2309)
);

HB1xp67_ASAP7_75t_L g2310 ( 
.A(n_2195),
.Y(n_2310)
);

INVx4_ASAP7_75t_L g2311 ( 
.A(n_2199),
.Y(n_2311)
);

AOI22xp5_ASAP7_75t_L g2312 ( 
.A1(n_2076),
.A2(n_1890),
.B1(n_1904),
.B2(n_1887),
.Y(n_2312)
);

INVx3_ASAP7_75t_L g2313 ( 
.A(n_2222),
.Y(n_2313)
);

BUFx6f_ASAP7_75t_L g2314 ( 
.A(n_2073),
.Y(n_2314)
);

INVx5_ASAP7_75t_L g2315 ( 
.A(n_2187),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_2111),
.B(n_2154),
.Y(n_2316)
);

INVxp33_ASAP7_75t_SL g2317 ( 
.A(n_2066),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_SL g2318 ( 
.A(n_2193),
.B(n_1921),
.Y(n_2318)
);

INVx1_ASAP7_75t_SL g2319 ( 
.A(n_2081),
.Y(n_2319)
);

BUFx8_ASAP7_75t_SL g2320 ( 
.A(n_2113),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2214),
.B(n_1925),
.Y(n_2321)
);

BUFx2_ASAP7_75t_L g2322 ( 
.A(n_2106),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2208),
.Y(n_2323)
);

BUFx6f_ASAP7_75t_L g2324 ( 
.A(n_2077),
.Y(n_2324)
);

OA21x2_ASAP7_75t_L g2325 ( 
.A1(n_2209),
.A2(n_1641),
.B(n_1621),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2217),
.B(n_1609),
.Y(n_2326)
);

OAI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_2129),
.A2(n_1956),
.B1(n_1966),
.B2(n_1927),
.Y(n_2327)
);

BUFx8_ASAP7_75t_L g2328 ( 
.A(n_2127),
.Y(n_2328)
);

BUFx3_ASAP7_75t_L g2329 ( 
.A(n_2194),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_L g2330 ( 
.A(n_2083),
.B(n_1967),
.Y(n_2330)
);

OAI22x1_ASAP7_75t_R g2331 ( 
.A1(n_2123),
.A2(n_2049),
.B1(n_1901),
.B2(n_1622),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2157),
.B(n_1609),
.Y(n_2332)
);

OAI22x1_ASAP7_75t_R g2333 ( 
.A1(n_2126),
.A2(n_1629),
.B1(n_1638),
.B2(n_1611),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2107),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2078),
.Y(n_2335)
);

OA21x2_ASAP7_75t_L g2336 ( 
.A1(n_2210),
.A2(n_2212),
.B(n_2211),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2218),
.B(n_1656),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2080),
.Y(n_2338)
);

OA21x2_ASAP7_75t_L g2339 ( 
.A1(n_2213),
.A2(n_1689),
.B(n_1675),
.Y(n_2339)
);

NAND2xp33_ASAP7_75t_L g2340 ( 
.A(n_2196),
.B(n_2000),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2082),
.Y(n_2341)
);

OAI22xp5_ASAP7_75t_SL g2342 ( 
.A1(n_2135),
.A2(n_1653),
.B1(n_1655),
.B2(n_1651),
.Y(n_2342)
);

OAI21x1_ASAP7_75t_L g2343 ( 
.A1(n_2215),
.A2(n_1719),
.B(n_1704),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2084),
.Y(n_2344)
);

OA21x2_ASAP7_75t_L g2345 ( 
.A1(n_2219),
.A2(n_1743),
.B(n_1739),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2198),
.B(n_2020),
.Y(n_2346)
);

NOR2xp33_ASAP7_75t_L g2347 ( 
.A(n_2201),
.B(n_2026),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2088),
.Y(n_2348)
);

INVx5_ASAP7_75t_L g2349 ( 
.A(n_2089),
.Y(n_2349)
);

AND2x4_ASAP7_75t_L g2350 ( 
.A(n_2202),
.B(n_1787),
.Y(n_2350)
);

BUFx6f_ASAP7_75t_L g2351 ( 
.A(n_2090),
.Y(n_2351)
);

BUFx6f_ASAP7_75t_L g2352 ( 
.A(n_2092),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2094),
.Y(n_2353)
);

HB1xp67_ASAP7_75t_L g2354 ( 
.A(n_2095),
.Y(n_2354)
);

CKINVDCx5p33_ASAP7_75t_R g2355 ( 
.A(n_2143),
.Y(n_2355)
);

CKINVDCx5p33_ASAP7_75t_R g2356 ( 
.A(n_2320),
.Y(n_2356)
);

CKINVDCx5p33_ASAP7_75t_R g2357 ( 
.A(n_2254),
.Y(n_2357)
);

CKINVDCx20_ASAP7_75t_R g2358 ( 
.A(n_2355),
.Y(n_2358)
);

CKINVDCx20_ASAP7_75t_R g2359 ( 
.A(n_2295),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2308),
.Y(n_2360)
);

CKINVDCx16_ASAP7_75t_R g2361 ( 
.A(n_2333),
.Y(n_2361)
);

OAI21x1_ASAP7_75t_L g2362 ( 
.A1(n_2297),
.A2(n_2221),
.B(n_2101),
.Y(n_2362)
);

CKINVDCx5p33_ASAP7_75t_R g2363 ( 
.A(n_2240),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2243),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2337),
.B(n_2100),
.Y(n_2365)
);

CKINVDCx5p33_ASAP7_75t_R g2366 ( 
.A(n_2239),
.Y(n_2366)
);

CKINVDCx5p33_ASAP7_75t_R g2367 ( 
.A(n_2249),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2224),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_2261),
.Y(n_2369)
);

CKINVDCx5p33_ASAP7_75t_R g2370 ( 
.A(n_2311),
.Y(n_2370)
);

AND2x6_ASAP7_75t_L g2371 ( 
.A(n_2332),
.B(n_2304),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2225),
.B(n_2227),
.Y(n_2372)
);

AO21x2_ASAP7_75t_L g2373 ( 
.A1(n_2299),
.A2(n_1457),
.B(n_1454),
.Y(n_2373)
);

CKINVDCx5p33_ASAP7_75t_R g2374 ( 
.A(n_2305),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_2310),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2323),
.Y(n_2376)
);

CKINVDCx5p33_ASAP7_75t_R g2377 ( 
.A(n_2322),
.Y(n_2377)
);

CKINVDCx5p33_ASAP7_75t_R g2378 ( 
.A(n_2315),
.Y(n_2378)
);

CKINVDCx20_ASAP7_75t_R g2379 ( 
.A(n_2319),
.Y(n_2379)
);

CKINVDCx20_ASAP7_75t_R g2380 ( 
.A(n_2266),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2237),
.B(n_2330),
.Y(n_2381)
);

CKINVDCx16_ASAP7_75t_R g2382 ( 
.A(n_2331),
.Y(n_2382)
);

CKINVDCx5p33_ASAP7_75t_R g2383 ( 
.A(n_2315),
.Y(n_2383)
);

BUFx6f_ASAP7_75t_SL g2384 ( 
.A(n_2233),
.Y(n_2384)
);

CKINVDCx5p33_ASAP7_75t_R g2385 ( 
.A(n_2317),
.Y(n_2385)
);

INVx3_ASAP7_75t_L g2386 ( 
.A(n_2309),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_R g2387 ( 
.A(n_2255),
.B(n_2169),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2265),
.Y(n_2388)
);

CKINVDCx20_ASAP7_75t_R g2389 ( 
.A(n_2342),
.Y(n_2389)
);

CKINVDCx5p33_ASAP7_75t_R g2390 ( 
.A(n_2293),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2314),
.Y(n_2391)
);

NOR2xp33_ASAP7_75t_R g2392 ( 
.A(n_2232),
.B(n_2170),
.Y(n_2392)
);

CKINVDCx5p33_ASAP7_75t_R g2393 ( 
.A(n_2252),
.Y(n_2393)
);

CKINVDCx5p33_ASAP7_75t_R g2394 ( 
.A(n_2234),
.Y(n_2394)
);

INVxp33_ASAP7_75t_L g2395 ( 
.A(n_2286),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2324),
.Y(n_2396)
);

BUFx8_ASAP7_75t_L g2397 ( 
.A(n_2326),
.Y(n_2397)
);

INVx3_ASAP7_75t_L g2398 ( 
.A(n_2336),
.Y(n_2398)
);

INVx3_ASAP7_75t_L g2399 ( 
.A(n_2251),
.Y(n_2399)
);

AND2x2_ASAP7_75t_L g2400 ( 
.A(n_2270),
.B(n_2105),
.Y(n_2400)
);

BUFx6f_ASAP7_75t_SL g2401 ( 
.A(n_2316),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2351),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2352),
.Y(n_2403)
);

CKINVDCx5p33_ASAP7_75t_R g2404 ( 
.A(n_2321),
.Y(n_2404)
);

CKINVDCx5p33_ASAP7_75t_R g2405 ( 
.A(n_2253),
.Y(n_2405)
);

CKINVDCx5p33_ASAP7_75t_R g2406 ( 
.A(n_2242),
.Y(n_2406)
);

CKINVDCx5p33_ASAP7_75t_R g2407 ( 
.A(n_2260),
.Y(n_2407)
);

HB1xp67_ASAP7_75t_L g2408 ( 
.A(n_2259),
.Y(n_2408)
);

CKINVDCx5p33_ASAP7_75t_R g2409 ( 
.A(n_2300),
.Y(n_2409)
);

CKINVDCx20_ASAP7_75t_R g2410 ( 
.A(n_2328),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_2263),
.Y(n_2411)
);

BUFx6f_ASAP7_75t_L g2412 ( 
.A(n_2236),
.Y(n_2412)
);

CKINVDCx20_ASAP7_75t_R g2413 ( 
.A(n_2303),
.Y(n_2413)
);

XOR2xp5_ASAP7_75t_L g2414 ( 
.A(n_2306),
.B(n_2197),
.Y(n_2414)
);

CKINVDCx5p33_ASAP7_75t_R g2415 ( 
.A(n_2269),
.Y(n_2415)
);

INVx1_ASAP7_75t_SL g2416 ( 
.A(n_2238),
.Y(n_2416)
);

CKINVDCx20_ASAP7_75t_R g2417 ( 
.A(n_2312),
.Y(n_2417)
);

INVx2_ASAP7_75t_SL g2418 ( 
.A(n_2285),
.Y(n_2418)
);

CKINVDCx5p33_ASAP7_75t_R g2419 ( 
.A(n_2256),
.Y(n_2419)
);

CKINVDCx5p33_ASAP7_75t_R g2420 ( 
.A(n_2327),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2272),
.Y(n_2421)
);

NOR2xp33_ASAP7_75t_R g2422 ( 
.A(n_2340),
.B(n_2200),
.Y(n_2422)
);

INVxp67_ASAP7_75t_L g2423 ( 
.A(n_2347),
.Y(n_2423)
);

CKINVDCx5p33_ASAP7_75t_R g2424 ( 
.A(n_2274),
.Y(n_2424)
);

CKINVDCx20_ASAP7_75t_R g2425 ( 
.A(n_2318),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2273),
.Y(n_2426)
);

OAI22xp5_ASAP7_75t_SL g2427 ( 
.A1(n_2229),
.A2(n_1716),
.B1(n_1724),
.B2(n_1701),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2283),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2288),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2276),
.Y(n_2430)
);

CKINVDCx5p33_ASAP7_75t_R g2431 ( 
.A(n_2231),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2289),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_2329),
.Y(n_2433)
);

NOR2xp33_ASAP7_75t_L g2434 ( 
.A(n_2226),
.B(n_1508),
.Y(n_2434)
);

BUFx6f_ASAP7_75t_L g2435 ( 
.A(n_2244),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_2302),
.Y(n_2436)
);

AND2x6_ASAP7_75t_L g2437 ( 
.A(n_2334),
.B(n_1458),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2343),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2278),
.Y(n_2439)
);

CKINVDCx5p33_ASAP7_75t_R g2440 ( 
.A(n_2354),
.Y(n_2440)
);

BUFx6f_ASAP7_75t_L g2441 ( 
.A(n_2223),
.Y(n_2441)
);

AO22x2_ASAP7_75t_L g2442 ( 
.A1(n_2241),
.A2(n_1959),
.B1(n_1963),
.B2(n_1682),
.Y(n_2442)
);

CKINVDCx5p33_ASAP7_75t_R g2443 ( 
.A(n_2228),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2282),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2245),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2335),
.Y(n_2446)
);

INVx3_ASAP7_75t_L g2447 ( 
.A(n_2268),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_2277),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2247),
.Y(n_2449)
);

INVx3_ASAP7_75t_L g2450 ( 
.A(n_2290),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2248),
.Y(n_2451)
);

CKINVDCx5p33_ASAP7_75t_R g2452 ( 
.A(n_2346),
.Y(n_2452)
);

NOR2xp33_ASAP7_75t_L g2453 ( 
.A(n_2230),
.B(n_1528),
.Y(n_2453)
);

CKINVDCx5p33_ASAP7_75t_R g2454 ( 
.A(n_2246),
.Y(n_2454)
);

CKINVDCx5p33_ASAP7_75t_R g2455 ( 
.A(n_2291),
.Y(n_2455)
);

BUFx6f_ASAP7_75t_L g2456 ( 
.A(n_2235),
.Y(n_2456)
);

CKINVDCx5p33_ASAP7_75t_R g2457 ( 
.A(n_2298),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2338),
.Y(n_2458)
);

INVx8_ASAP7_75t_L g2459 ( 
.A(n_2350),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2250),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2341),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2344),
.Y(n_2462)
);

NOR2xp33_ASAP7_75t_R g2463 ( 
.A(n_2313),
.B(n_1730),
.Y(n_2463)
);

CKINVDCx5p33_ASAP7_75t_R g2464 ( 
.A(n_2348),
.Y(n_2464)
);

CKINVDCx20_ASAP7_75t_R g2465 ( 
.A(n_2353),
.Y(n_2465)
);

HB1xp67_ASAP7_75t_L g2466 ( 
.A(n_2307),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_SL g2467 ( 
.A(n_2349),
.B(n_1404),
.Y(n_2467)
);

BUFx3_ASAP7_75t_L g2468 ( 
.A(n_2325),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2257),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_2279),
.Y(n_2470)
);

CKINVDCx5p33_ASAP7_75t_R g2471 ( 
.A(n_2349),
.Y(n_2471)
);

HB1xp67_ASAP7_75t_L g2472 ( 
.A(n_2339),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2271),
.Y(n_2473)
);

CKINVDCx20_ASAP7_75t_R g2474 ( 
.A(n_2345),
.Y(n_2474)
);

NOR2xp33_ASAP7_75t_R g2475 ( 
.A(n_2258),
.B(n_1760),
.Y(n_2475)
);

CKINVDCx20_ASAP7_75t_R g2476 ( 
.A(n_2262),
.Y(n_2476)
);

CKINVDCx5p33_ASAP7_75t_R g2477 ( 
.A(n_2287),
.Y(n_2477)
);

CKINVDCx5p33_ASAP7_75t_R g2478 ( 
.A(n_2296),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2264),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_2275),
.Y(n_2480)
);

CKINVDCx20_ASAP7_75t_R g2481 ( 
.A(n_2281),
.Y(n_2481)
);

CKINVDCx5p33_ASAP7_75t_R g2482 ( 
.A(n_2292),
.Y(n_2482)
);

CKINVDCx20_ASAP7_75t_R g2483 ( 
.A(n_2294),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2301),
.Y(n_2484)
);

CKINVDCx5p33_ASAP7_75t_R g2485 ( 
.A(n_2280),
.Y(n_2485)
);

NOR2xp33_ASAP7_75t_L g2486 ( 
.A(n_2299),
.B(n_1555),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2284),
.Y(n_2487)
);

BUFx3_ASAP7_75t_L g2488 ( 
.A(n_2234),
.Y(n_2488)
);

CKINVDCx5p33_ASAP7_75t_R g2489 ( 
.A(n_2320),
.Y(n_2489)
);

CKINVDCx5p33_ASAP7_75t_R g2490 ( 
.A(n_2320),
.Y(n_2490)
);

CKINVDCx5p33_ASAP7_75t_R g2491 ( 
.A(n_2320),
.Y(n_2491)
);

AND2x2_ASAP7_75t_L g2492 ( 
.A(n_2337),
.B(n_2114),
.Y(n_2492)
);

CKINVDCx5p33_ASAP7_75t_R g2493 ( 
.A(n_2320),
.Y(n_2493)
);

CKINVDCx20_ASAP7_75t_R g2494 ( 
.A(n_2320),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2267),
.Y(n_2495)
);

CKINVDCx5p33_ASAP7_75t_R g2496 ( 
.A(n_2320),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2404),
.B(n_2117),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2360),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2381),
.B(n_2118),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2443),
.B(n_2120),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2376),
.Y(n_2501)
);

BUFx10_ASAP7_75t_L g2502 ( 
.A(n_2356),
.Y(n_2502)
);

OAI22xp33_ASAP7_75t_L g2503 ( 
.A1(n_2419),
.A2(n_1483),
.B1(n_1513),
.B2(n_1495),
.Y(n_2503)
);

INVx4_ASAP7_75t_SL g2504 ( 
.A(n_2401),
.Y(n_2504)
);

INVx4_ASAP7_75t_L g2505 ( 
.A(n_2405),
.Y(n_2505)
);

AND2x4_ASAP7_75t_L g2506 ( 
.A(n_2488),
.B(n_2124),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2445),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2449),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2451),
.Y(n_2509)
);

AND2x6_ASAP7_75t_L g2510 ( 
.A(n_2438),
.B(n_1461),
.Y(n_2510)
);

INVxp67_ASAP7_75t_SL g2511 ( 
.A(n_2466),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2460),
.Y(n_2512)
);

INVx3_ASAP7_75t_L g2513 ( 
.A(n_2412),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2469),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2479),
.Y(n_2515)
);

AND2x6_ASAP7_75t_L g2516 ( 
.A(n_2473),
.B(n_1463),
.Y(n_2516)
);

INVx5_ASAP7_75t_L g2517 ( 
.A(n_2412),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_L g2518 ( 
.A(n_2423),
.B(n_1520),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_SL g2519 ( 
.A(n_2452),
.B(n_1408),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2484),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2446),
.Y(n_2521)
);

AOI22xp5_ASAP7_75t_L g2522 ( 
.A1(n_2474),
.A2(n_1770),
.B1(n_1791),
.B2(n_1780),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_SL g2523 ( 
.A(n_2418),
.B(n_1411),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2492),
.B(n_2130),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2458),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2461),
.Y(n_2526)
);

AND2x4_ASAP7_75t_L g2527 ( 
.A(n_2388),
.B(n_2131),
.Y(n_2527)
);

BUFx6f_ASAP7_75t_L g2528 ( 
.A(n_2435),
.Y(n_2528)
);

BUFx6f_ASAP7_75t_L g2529 ( 
.A(n_2435),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2486),
.B(n_2132),
.Y(n_2530)
);

AND2x2_ASAP7_75t_SL g2531 ( 
.A(n_2361),
.B(n_1828),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2462),
.Y(n_2532)
);

AND2x4_ASAP7_75t_L g2533 ( 
.A(n_2421),
.B(n_2133),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2472),
.B(n_2386),
.Y(n_2534)
);

AND2x6_ASAP7_75t_L g2535 ( 
.A(n_2386),
.B(n_1465),
.Y(n_2535)
);

BUFx3_ASAP7_75t_L g2536 ( 
.A(n_2455),
.Y(n_2536)
);

BUFx2_ASAP7_75t_L g2537 ( 
.A(n_2463),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2362),
.Y(n_2538)
);

AND2x6_ASAP7_75t_L g2539 ( 
.A(n_2398),
.B(n_1468),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2364),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2468),
.Y(n_2541)
);

BUFx4f_ASAP7_75t_L g2542 ( 
.A(n_2371),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2399),
.B(n_2447),
.Y(n_2543)
);

CKINVDCx20_ASAP7_75t_R g2544 ( 
.A(n_2358),
.Y(n_2544)
);

BUFx2_ASAP7_75t_L g2545 ( 
.A(n_2379),
.Y(n_2545)
);

AND2x4_ASAP7_75t_L g2546 ( 
.A(n_2426),
.B(n_2147),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2495),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2399),
.Y(n_2548)
);

BUFx2_ASAP7_75t_L g2549 ( 
.A(n_2392),
.Y(n_2549)
);

AND2x2_ASAP7_75t_SL g2550 ( 
.A(n_2382),
.B(n_1831),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_L g2551 ( 
.A(n_2390),
.B(n_1522),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2373),
.B(n_2434),
.Y(n_2552)
);

INVxp67_ASAP7_75t_L g2553 ( 
.A(n_2453),
.Y(n_2553)
);

AND2x2_ASAP7_75t_L g2554 ( 
.A(n_2400),
.B(n_1656),
.Y(n_2554)
);

NOR2xp33_ASAP7_75t_L g2555 ( 
.A(n_2420),
.B(n_1524),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2372),
.Y(n_2556)
);

BUFx10_ASAP7_75t_L g2557 ( 
.A(n_2489),
.Y(n_2557)
);

BUFx6f_ASAP7_75t_L g2558 ( 
.A(n_2441),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_2464),
.B(n_1550),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2487),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2428),
.Y(n_2561)
);

BUFx10_ASAP7_75t_L g2562 ( 
.A(n_2490),
.Y(n_2562)
);

INVx6_ASAP7_75t_L g2563 ( 
.A(n_2456),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2429),
.Y(n_2564)
);

BUFx3_ASAP7_75t_L g2565 ( 
.A(n_2457),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2430),
.Y(n_2566)
);

AND2x6_ASAP7_75t_L g2567 ( 
.A(n_2432),
.B(n_1479),
.Y(n_2567)
);

INVx4_ASAP7_75t_L g2568 ( 
.A(n_2454),
.Y(n_2568)
);

NOR2xp33_ASAP7_75t_L g2569 ( 
.A(n_2436),
.B(n_1552),
.Y(n_2569)
);

INVx4_ASAP7_75t_L g2570 ( 
.A(n_2470),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2439),
.Y(n_2571)
);

INVx6_ASAP7_75t_L g2572 ( 
.A(n_2456),
.Y(n_2572)
);

AOI22xp33_ASAP7_75t_L g2573 ( 
.A1(n_2485),
.A2(n_1938),
.B1(n_1974),
.B2(n_1928),
.Y(n_2573)
);

NOR2xp33_ASAP7_75t_L g2574 ( 
.A(n_2440),
.B(n_1579),
.Y(n_2574)
);

OAI22xp33_ASAP7_75t_L g2575 ( 
.A1(n_2431),
.A2(n_1613),
.B1(n_1694),
.B2(n_1588),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2477),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_SL g2577 ( 
.A(n_2366),
.B(n_1422),
.Y(n_2577)
);

INVx3_ASAP7_75t_L g2578 ( 
.A(n_2456),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2433),
.B(n_1667),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2478),
.Y(n_2580)
);

INVx4_ASAP7_75t_L g2581 ( 
.A(n_2459),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2437),
.B(n_2371),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2437),
.B(n_1423),
.Y(n_2583)
);

INVx3_ASAP7_75t_L g2584 ( 
.A(n_2444),
.Y(n_2584)
);

CKINVDCx20_ASAP7_75t_R g2585 ( 
.A(n_2359),
.Y(n_2585)
);

AND2x4_ASAP7_75t_L g2586 ( 
.A(n_2450),
.B(n_2150),
.Y(n_2586)
);

INVx4_ASAP7_75t_L g2587 ( 
.A(n_2459),
.Y(n_2587)
);

NOR2xp33_ASAP7_75t_L g2588 ( 
.A(n_2480),
.B(n_1754),
.Y(n_2588)
);

INVx4_ASAP7_75t_SL g2589 ( 
.A(n_2401),
.Y(n_2589)
);

NAND2x1p5_ASAP7_75t_L g2590 ( 
.A(n_2450),
.B(n_2153),
.Y(n_2590)
);

NOR2xp33_ASAP7_75t_L g2591 ( 
.A(n_2482),
.B(n_1773),
.Y(n_2591)
);

AO22x2_ASAP7_75t_L g2592 ( 
.A1(n_2414),
.A2(n_2001),
.B1(n_2013),
.B2(n_1812),
.Y(n_2592)
);

INVx4_ASAP7_75t_L g2593 ( 
.A(n_2394),
.Y(n_2593)
);

BUFx3_ASAP7_75t_L g2594 ( 
.A(n_2380),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2391),
.Y(n_2595)
);

HB1xp67_ASAP7_75t_L g2596 ( 
.A(n_2475),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2396),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2402),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2403),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2367),
.B(n_1427),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2369),
.B(n_1428),
.Y(n_2601)
);

NOR2xp33_ASAP7_75t_L g2602 ( 
.A(n_2415),
.B(n_1983),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2408),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2374),
.B(n_2375),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_2370),
.B(n_2031),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2465),
.Y(n_2606)
);

CKINVDCx5p33_ASAP7_75t_R g2607 ( 
.A(n_2491),
.Y(n_2607)
);

NOR2xp33_ASAP7_75t_L g2608 ( 
.A(n_2411),
.B(n_1432),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2442),
.Y(n_2609)
);

OAI22xp5_ASAP7_75t_L g2610 ( 
.A1(n_2424),
.A2(n_1435),
.B1(n_1436),
.B2(n_1433),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2476),
.Y(n_2611)
);

INVx2_ASAP7_75t_SL g2612 ( 
.A(n_2481),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2483),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2467),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2422),
.B(n_1439),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2471),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2406),
.B(n_1442),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2378),
.B(n_1443),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2384),
.Y(n_2619)
);

AOI22xp33_ASAP7_75t_L g2620 ( 
.A1(n_2395),
.A2(n_2384),
.B1(n_2427),
.B2(n_2417),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2387),
.B(n_2385),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_SL g2622 ( 
.A(n_2383),
.B(n_1444),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2425),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_SL g2624 ( 
.A(n_2397),
.B(n_1446),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2397),
.Y(n_2625)
);

NAND2x1p5_ASAP7_75t_L g2626 ( 
.A(n_2416),
.B(n_2155),
.Y(n_2626)
);

INVx4_ASAP7_75t_L g2627 ( 
.A(n_2363),
.Y(n_2627)
);

HB1xp67_ASAP7_75t_L g2628 ( 
.A(n_2377),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2413),
.Y(n_2629)
);

INVx4_ASAP7_75t_L g2630 ( 
.A(n_2493),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_SL g2631 ( 
.A(n_2389),
.B(n_1453),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2496),
.Y(n_2632)
);

NAND3x1_ASAP7_75t_L g2633 ( 
.A(n_2410),
.B(n_1482),
.C(n_1481),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2407),
.Y(n_2634)
);

BUFx6f_ASAP7_75t_L g2635 ( 
.A(n_2409),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2494),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2393),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2360),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2360),
.Y(n_2639)
);

AND2x2_ASAP7_75t_SL g2640 ( 
.A(n_2361),
.B(n_2029),
.Y(n_2640)
);

INVx2_ASAP7_75t_SL g2641 ( 
.A(n_2365),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2381),
.B(n_1761),
.Y(n_2642)
);

INVxp67_ASAP7_75t_SL g2643 ( 
.A(n_2466),
.Y(n_2643)
);

INVx1_ASAP7_75t_SL g2644 ( 
.A(n_2463),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_SL g2645 ( 
.A(n_2448),
.B(n_1455),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2381),
.B(n_1761),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2368),
.Y(n_2647)
);

BUFx6f_ASAP7_75t_SL g2648 ( 
.A(n_2488),
.Y(n_2648)
);

AOI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_2474),
.A2(n_1894),
.B1(n_1912),
.B2(n_1886),
.Y(n_2649)
);

INVx3_ASAP7_75t_L g2650 ( 
.A(n_2412),
.Y(n_2650)
);

BUFx6f_ASAP7_75t_L g2651 ( 
.A(n_2412),
.Y(n_2651)
);

OR2x2_ASAP7_75t_L g2652 ( 
.A(n_2381),
.B(n_2160),
.Y(n_2652)
);

INVx4_ASAP7_75t_L g2653 ( 
.A(n_2405),
.Y(n_2653)
);

NOR2xp33_ASAP7_75t_L g2654 ( 
.A(n_2448),
.B(n_1462),
.Y(n_2654)
);

NOR2xp33_ASAP7_75t_L g2655 ( 
.A(n_2448),
.B(n_1469),
.Y(n_2655)
);

AND2x4_ASAP7_75t_L g2656 ( 
.A(n_2488),
.B(n_2161),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_SL g2657 ( 
.A(n_2448),
.B(n_1472),
.Y(n_2657)
);

BUFx6f_ASAP7_75t_L g2658 ( 
.A(n_2412),
.Y(n_2658)
);

INVx3_ASAP7_75t_L g2659 ( 
.A(n_2412),
.Y(n_2659)
);

AND2x6_ASAP7_75t_L g2660 ( 
.A(n_2438),
.B(n_1484),
.Y(n_2660)
);

BUFx10_ASAP7_75t_L g2661 ( 
.A(n_2356),
.Y(n_2661)
);

NOR2xp33_ASAP7_75t_R g2662 ( 
.A(n_2356),
.B(n_1916),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2404),
.B(n_1473),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2404),
.B(n_1474),
.Y(n_2664)
);

NOR2xp33_ASAP7_75t_SL g2665 ( 
.A(n_2357),
.B(n_1918),
.Y(n_2665)
);

BUFx2_ASAP7_75t_L g2666 ( 
.A(n_2463),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2404),
.B(n_1475),
.Y(n_2667)
);

OR2x2_ASAP7_75t_L g2668 ( 
.A(n_2381),
.B(n_2162),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2404),
.B(n_1476),
.Y(n_2669)
);

AOI22xp33_ASAP7_75t_L g2670 ( 
.A1(n_2386),
.A2(n_2042),
.B1(n_2047),
.B2(n_2040),
.Y(n_2670)
);

BUFx6f_ASAP7_75t_L g2671 ( 
.A(n_2412),
.Y(n_2671)
);

AOI22xp33_ASAP7_75t_L g2672 ( 
.A1(n_2386),
.A2(n_2056),
.B1(n_2050),
.B2(n_1489),
.Y(n_2672)
);

INVx4_ASAP7_75t_L g2673 ( 
.A(n_2405),
.Y(n_2673)
);

NOR2xp33_ASAP7_75t_L g2674 ( 
.A(n_2448),
.B(n_1480),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2360),
.Y(n_2675)
);

CKINVDCx20_ASAP7_75t_R g2676 ( 
.A(n_2358),
.Y(n_2676)
);

BUFx2_ASAP7_75t_L g2677 ( 
.A(n_2463),
.Y(n_2677)
);

BUFx6f_ASAP7_75t_L g2678 ( 
.A(n_2412),
.Y(n_2678)
);

NOR2xp33_ASAP7_75t_L g2679 ( 
.A(n_2602),
.B(n_1952),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2498),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2548),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2518),
.B(n_1851),
.Y(n_2682)
);

NOR2xp33_ASAP7_75t_L g2683 ( 
.A(n_2555),
.B(n_1979),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2511),
.B(n_1485),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2643),
.B(n_1486),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2499),
.B(n_1491),
.Y(n_2686)
);

AOI22xp33_ASAP7_75t_L g2687 ( 
.A1(n_2535),
.A2(n_1493),
.B1(n_1503),
.B2(n_1487),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2541),
.Y(n_2688)
);

NOR2xp33_ASAP7_75t_L g2689 ( 
.A(n_2569),
.B(n_1494),
.Y(n_2689)
);

AOI22xp33_ASAP7_75t_L g2690 ( 
.A1(n_2535),
.A2(n_2539),
.B1(n_2516),
.B2(n_2510),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_SL g2691 ( 
.A(n_2663),
.B(n_1496),
.Y(n_2691)
);

NOR2xp33_ASAP7_75t_L g2692 ( 
.A(n_2605),
.B(n_1497),
.Y(n_2692)
);

AND2x6_ASAP7_75t_SL g2693 ( 
.A(n_2604),
.B(n_1506),
.Y(n_2693)
);

AOI22xp5_ASAP7_75t_L g2694 ( 
.A1(n_2608),
.A2(n_1499),
.B1(n_1500),
.B2(n_1498),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2530),
.B(n_1504),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2534),
.B(n_1505),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2500),
.B(n_1507),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2497),
.B(n_1509),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2642),
.B(n_1511),
.Y(n_2699)
);

NOR2xp33_ASAP7_75t_L g2700 ( 
.A(n_2588),
.B(n_1516),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2646),
.B(n_1518),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2501),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_SL g2703 ( 
.A(n_2664),
.B(n_1521),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2543),
.B(n_1523),
.Y(n_2704)
);

NOR2xp33_ASAP7_75t_L g2705 ( 
.A(n_2591),
.B(n_1526),
.Y(n_2705)
);

NOR2xp33_ASAP7_75t_L g2706 ( 
.A(n_2617),
.B(n_1527),
.Y(n_2706)
);

AND2x6_ASAP7_75t_L g2707 ( 
.A(n_2582),
.B(n_1510),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_SL g2708 ( 
.A(n_2667),
.B(n_1529),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2524),
.B(n_1531),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2654),
.B(n_1532),
.Y(n_2710)
);

NOR2xp33_ASAP7_75t_L g2711 ( 
.A(n_2655),
.B(n_2674),
.Y(n_2711)
);

NOR2xp33_ASAP7_75t_L g2712 ( 
.A(n_2559),
.B(n_1533),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2641),
.B(n_1534),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_SL g2714 ( 
.A(n_2669),
.B(n_1537),
.Y(n_2714)
);

AND2x4_ASAP7_75t_L g2715 ( 
.A(n_2504),
.B(n_2163),
.Y(n_2715)
);

NOR2xp33_ASAP7_75t_L g2716 ( 
.A(n_2574),
.B(n_1538),
.Y(n_2716)
);

INVx2_ASAP7_75t_SL g2717 ( 
.A(n_2572),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2647),
.Y(n_2718)
);

NOR2xp33_ASAP7_75t_L g2719 ( 
.A(n_2553),
.B(n_1553),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_SL g2720 ( 
.A(n_2542),
.B(n_1557),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2554),
.B(n_1920),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2514),
.Y(n_2722)
);

NOR3xp33_ASAP7_75t_L g2723 ( 
.A(n_2631),
.B(n_1566),
.C(n_1565),
.Y(n_2723)
);

AND2x2_ASAP7_75t_L g2724 ( 
.A(n_2579),
.B(n_1920),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2638),
.Y(n_2725)
);

NOR2xp33_ASAP7_75t_L g2726 ( 
.A(n_2644),
.B(n_1568),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2639),
.B(n_1576),
.Y(n_2727)
);

BUFx2_ASAP7_75t_L g2728 ( 
.A(n_2545),
.Y(n_2728)
);

BUFx6f_ASAP7_75t_L g2729 ( 
.A(n_2528),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2675),
.B(n_1580),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2652),
.B(n_1582),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2668),
.B(n_1584),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2573),
.B(n_1590),
.Y(n_2733)
);

AOI22xp5_ASAP7_75t_L g2734 ( 
.A1(n_2539),
.A2(n_1594),
.B1(n_1598),
.B2(n_1593),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2507),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2672),
.B(n_1600),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2508),
.Y(n_2737)
);

INVx2_ASAP7_75t_SL g2738 ( 
.A(n_2656),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2509),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2512),
.B(n_1605),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2540),
.Y(n_2741)
);

A2O1A1Ixp33_ASAP7_75t_L g2742 ( 
.A1(n_2614),
.A2(n_1540),
.B(n_1542),
.C(n_1539),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2546),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2515),
.B(n_1606),
.Y(n_2744)
);

AND2x2_ASAP7_75t_L g2745 ( 
.A(n_2576),
.B(n_2580),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2520),
.B(n_1607),
.Y(n_2746)
);

AOI21xp5_ASAP7_75t_L g2747 ( 
.A1(n_2538),
.A2(n_1545),
.B(n_1543),
.Y(n_2747)
);

NOR2xp33_ASAP7_75t_L g2748 ( 
.A(n_2596),
.B(n_1612),
.Y(n_2748)
);

INVx2_ASAP7_75t_SL g2749 ( 
.A(n_2506),
.Y(n_2749)
);

NOR2xp33_ASAP7_75t_L g2750 ( 
.A(n_2522),
.B(n_1617),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2521),
.B(n_1620),
.Y(n_2751)
);

AND2x2_ASAP7_75t_L g2752 ( 
.A(n_2549),
.B(n_1973),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2525),
.B(n_1623),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2547),
.Y(n_2754)
);

OAI22xp5_ASAP7_75t_L g2755 ( 
.A1(n_2670),
.A2(n_1627),
.B1(n_1628),
.B2(n_1624),
.Y(n_2755)
);

AOI22xp33_ASAP7_75t_L g2756 ( 
.A1(n_2510),
.A2(n_1547),
.B1(n_1549),
.B2(n_1546),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2526),
.B(n_1631),
.Y(n_2757)
);

NOR2xp33_ASAP7_75t_L g2758 ( 
.A(n_2649),
.B(n_1635),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_SL g2759 ( 
.A(n_2600),
.B(n_1637),
.Y(n_2759)
);

O2A1O1Ixp33_ASAP7_75t_L g2760 ( 
.A1(n_2609),
.A2(n_1559),
.B(n_1567),
.C(n_1554),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2532),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2601),
.B(n_2510),
.Y(n_2762)
);

BUFx2_ASAP7_75t_L g2763 ( 
.A(n_2613),
.Y(n_2763)
);

NOR2x1p5_ASAP7_75t_L g2764 ( 
.A(n_2536),
.B(n_1640),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2527),
.Y(n_2765)
);

AOI22xp33_ASAP7_75t_L g2766 ( 
.A1(n_2660),
.A2(n_1572),
.B1(n_1573),
.B2(n_1571),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2533),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_SL g2768 ( 
.A(n_2537),
.B(n_1642),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_SL g2769 ( 
.A(n_2666),
.B(n_1645),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2561),
.B(n_1646),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2564),
.B(n_1652),
.Y(n_2771)
);

AOI22xp5_ASAP7_75t_L g2772 ( 
.A1(n_2519),
.A2(n_1665),
.B1(n_1666),
.B2(n_1664),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2615),
.B(n_1668),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2586),
.Y(n_2774)
);

OAI22x1_ASAP7_75t_R g2775 ( 
.A1(n_2585),
.A2(n_2676),
.B1(n_2544),
.B2(n_2607),
.Y(n_2775)
);

NOR3xp33_ASAP7_75t_L g2776 ( 
.A(n_2503),
.B(n_1670),
.C(n_1669),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_SL g2777 ( 
.A(n_2677),
.B(n_1671),
.Y(n_2777)
);

NOR2xp33_ASAP7_75t_L g2778 ( 
.A(n_2645),
.B(n_1673),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2597),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2599),
.Y(n_2780)
);

AOI22xp5_ASAP7_75t_L g2781 ( 
.A1(n_2657),
.A2(n_1677),
.B1(n_1679),
.B2(n_1676),
.Y(n_2781)
);

INVx2_ASAP7_75t_SL g2782 ( 
.A(n_2529),
.Y(n_2782)
);

OAI22xp5_ASAP7_75t_L g2783 ( 
.A1(n_2603),
.A2(n_1684),
.B1(n_1685),
.B2(n_1681),
.Y(n_2783)
);

NOR3xp33_ASAP7_75t_L g2784 ( 
.A(n_2575),
.B(n_1690),
.C(n_1687),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_SL g2785 ( 
.A(n_2665),
.B(n_1692),
.Y(n_2785)
);

AOI22xp33_ASAP7_75t_L g2786 ( 
.A1(n_2567),
.A2(n_1619),
.B1(n_1625),
.B2(n_1599),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2560),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_2566),
.Y(n_2788)
);

NOR3xp33_ASAP7_75t_L g2789 ( 
.A(n_2612),
.B(n_1709),
.C(n_1706),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_SL g2790 ( 
.A(n_2570),
.B(n_1712),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2571),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2595),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2583),
.B(n_1715),
.Y(n_2793)
);

NOR3xp33_ASAP7_75t_L g2794 ( 
.A(n_2611),
.B(n_1718),
.C(n_1717),
.Y(n_2794)
);

NAND3xp33_ASAP7_75t_L g2795 ( 
.A(n_2610),
.B(n_1721),
.C(n_1720),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2567),
.B(n_1723),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2567),
.B(n_1725),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_SL g2798 ( 
.A(n_2621),
.B(n_1726),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2598),
.Y(n_2799)
);

AND2x4_ASAP7_75t_L g2800 ( 
.A(n_2589),
.B(n_2581),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2577),
.B(n_2523),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2618),
.B(n_1727),
.Y(n_2802)
);

OR2x6_ASAP7_75t_L g2803 ( 
.A(n_2565),
.B(n_1626),
.Y(n_2803)
);

NOR2xp67_ASAP7_75t_L g2804 ( 
.A(n_2505),
.B(n_1728),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_2584),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2513),
.Y(n_2806)
);

AND2x6_ASAP7_75t_SL g2807 ( 
.A(n_2629),
.B(n_1632),
.Y(n_2807)
);

NOR2xp33_ASAP7_75t_L g2808 ( 
.A(n_2626),
.B(n_1732),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_SL g2809 ( 
.A(n_2653),
.B(n_1733),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_SL g2810 ( 
.A(n_2673),
.B(n_1734),
.Y(n_2810)
);

CKINVDCx5p33_ASAP7_75t_R g2811 ( 
.A(n_2662),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2578),
.B(n_1735),
.Y(n_2812)
);

NAND3xp33_ASAP7_75t_L g2813 ( 
.A(n_2620),
.B(n_1741),
.C(n_1740),
.Y(n_2813)
);

NOR2xp33_ASAP7_75t_L g2814 ( 
.A(n_2623),
.B(n_1742),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_SL g2815 ( 
.A(n_2568),
.B(n_1744),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2650),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2659),
.B(n_1745),
.Y(n_2817)
);

NOR2xp33_ASAP7_75t_L g2818 ( 
.A(n_2628),
.B(n_1746),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2558),
.B(n_1747),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2590),
.Y(n_2820)
);

NOR2x1p5_ASAP7_75t_L g2821 ( 
.A(n_2587),
.B(n_1752),
.Y(n_2821)
);

NOR2xp33_ASAP7_75t_L g2822 ( 
.A(n_2606),
.B(n_1756),
.Y(n_2822)
);

INVx8_ASAP7_75t_L g2823 ( 
.A(n_2517),
.Y(n_2823)
);

AOI21xp5_ASAP7_75t_L g2824 ( 
.A1(n_2622),
.A2(n_1634),
.B(n_1633),
.Y(n_2824)
);

OAI22xp33_ASAP7_75t_L g2825 ( 
.A1(n_2619),
.A2(n_1758),
.B1(n_1762),
.B2(n_1757),
.Y(n_2825)
);

AOI22xp33_ASAP7_75t_L g2826 ( 
.A1(n_2592),
.A2(n_2616),
.B1(n_2550),
.B2(n_2531),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_SL g2827 ( 
.A(n_2651),
.B(n_1765),
.Y(n_2827)
);

INVx3_ASAP7_75t_L g2828 ( 
.A(n_2658),
.Y(n_2828)
);

AOI22xp5_ASAP7_75t_L g2829 ( 
.A1(n_2632),
.A2(n_1775),
.B1(n_1776),
.B2(n_1768),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2658),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2671),
.B(n_1777),
.Y(n_2831)
);

A2O1A1Ixp33_ASAP7_75t_L g2832 ( 
.A1(n_2640),
.A2(n_1648),
.B(n_1649),
.C(n_1643),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2671),
.B(n_1778),
.Y(n_2833)
);

OR2x6_ASAP7_75t_L g2834 ( 
.A(n_2635),
.B(n_1659),
.Y(n_2834)
);

NAND2xp33_ASAP7_75t_L g2835 ( 
.A(n_2678),
.B(n_1781),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2627),
.B(n_1782),
.Y(n_2836)
);

AND2x2_ASAP7_75t_L g2837 ( 
.A(n_2594),
.B(n_2630),
.Y(n_2837)
);

AOI22xp33_ASAP7_75t_L g2838 ( 
.A1(n_2624),
.A2(n_1662),
.B1(n_1663),
.B2(n_1660),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2634),
.B(n_1784),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2637),
.B(n_1785),
.Y(n_2840)
);

AOI22xp5_ASAP7_75t_L g2841 ( 
.A1(n_2648),
.A2(n_1789),
.B1(n_1790),
.B2(n_1788),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2636),
.B(n_1792),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2633),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_SL g2844 ( 
.A(n_2502),
.B(n_1793),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2557),
.B(n_1794),
.Y(n_2845)
);

BUFx3_ASAP7_75t_L g2846 ( 
.A(n_2635),
.Y(n_2846)
);

AOI22xp5_ASAP7_75t_L g2847 ( 
.A1(n_2625),
.A2(n_1797),
.B1(n_1798),
.B2(n_1795),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2562),
.B(n_1801),
.Y(n_2848)
);

NOR2xp33_ASAP7_75t_L g2849 ( 
.A(n_2661),
.B(n_1802),
.Y(n_2849)
);

BUFx6f_ASAP7_75t_L g2850 ( 
.A(n_2528),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2556),
.B(n_1804),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2556),
.B(n_1806),
.Y(n_2852)
);

INVx2_ASAP7_75t_SL g2853 ( 
.A(n_2563),
.Y(n_2853)
);

INVx5_ASAP7_75t_L g2854 ( 
.A(n_2535),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_SL g2855 ( 
.A(n_2556),
.B(n_1807),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2556),
.B(n_1808),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_SL g2857 ( 
.A(n_2556),
.B(n_1813),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2548),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2498),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2556),
.B(n_1814),
.Y(n_2860)
);

AOI22xp5_ASAP7_75t_L g2861 ( 
.A1(n_2556),
.A2(n_1819),
.B1(n_1821),
.B2(n_1815),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2498),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2498),
.Y(n_2863)
);

INVx4_ASAP7_75t_L g2864 ( 
.A(n_2581),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2551),
.B(n_1825),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2548),
.Y(n_2866)
);

NOR2xp33_ASAP7_75t_L g2867 ( 
.A(n_2551),
.B(n_1826),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2548),
.Y(n_2868)
);

NOR2xp67_ASAP7_75t_SL g2869 ( 
.A(n_2593),
.B(n_1697),
.Y(n_2869)
);

NOR2xp33_ASAP7_75t_L g2870 ( 
.A(n_2551),
.B(n_1829),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_SL g2871 ( 
.A(n_2556),
.B(n_1832),
.Y(n_2871)
);

INVx4_ASAP7_75t_L g2872 ( 
.A(n_2581),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_SL g2873 ( 
.A(n_2556),
.B(n_1833),
.Y(n_2873)
);

INVx2_ASAP7_75t_SL g2874 ( 
.A(n_2563),
.Y(n_2874)
);

BUFx3_ASAP7_75t_L g2875 ( 
.A(n_2536),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2556),
.B(n_1835),
.Y(n_2876)
);

NOR2xp33_ASAP7_75t_L g2877 ( 
.A(n_2551),
.B(n_1839),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_2548),
.Y(n_2878)
);

NOR2xp33_ASAP7_75t_L g2879 ( 
.A(n_2551),
.B(n_1841),
.Y(n_2879)
);

INVx2_ASAP7_75t_L g2880 ( 
.A(n_2548),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2556),
.B(n_1845),
.Y(n_2881)
);

INVx8_ASAP7_75t_L g2882 ( 
.A(n_2517),
.Y(n_2882)
);

A2O1A1Ixp33_ASAP7_75t_L g2883 ( 
.A1(n_2552),
.A2(n_1702),
.B(n_1703),
.C(n_1700),
.Y(n_2883)
);

INVx4_ASAP7_75t_L g2884 ( 
.A(n_2823),
.Y(n_2884)
);

AO21x1_ASAP7_75t_L g2885 ( 
.A1(n_2711),
.A2(n_1711),
.B(n_1710),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2681),
.Y(n_2886)
);

INVx3_ASAP7_75t_L g2887 ( 
.A(n_2875),
.Y(n_2887)
);

OR2x6_ASAP7_75t_L g2888 ( 
.A(n_2823),
.B(n_1713),
.Y(n_2888)
);

INVx3_ASAP7_75t_L g2889 ( 
.A(n_2846),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_SL g2890 ( 
.A(n_2745),
.B(n_1849),
.Y(n_2890)
);

HB1xp67_ASAP7_75t_L g2891 ( 
.A(n_2763),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2689),
.B(n_1850),
.Y(n_2892)
);

AND2x2_ASAP7_75t_L g2893 ( 
.A(n_2682),
.B(n_1854),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2706),
.B(n_1858),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2865),
.B(n_1859),
.Y(n_2895)
);

NOR2xp33_ASAP7_75t_L g2896 ( 
.A(n_2683),
.B(n_1860),
.Y(n_2896)
);

AOI21xp5_ASAP7_75t_L g2897 ( 
.A1(n_2762),
.A2(n_1731),
.B(n_1729),
.Y(n_2897)
);

NOR2xp33_ASAP7_75t_L g2898 ( 
.A(n_2679),
.B(n_1862),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2867),
.B(n_1863),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2870),
.B(n_1865),
.Y(n_2900)
);

AOI21xp5_ASAP7_75t_L g2901 ( 
.A1(n_2801),
.A2(n_1737),
.B(n_1736),
.Y(n_2901)
);

AOI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2704),
.A2(n_1749),
.B(n_1748),
.Y(n_2902)
);

A2O1A1Ixp33_ASAP7_75t_L g2903 ( 
.A1(n_2877),
.A2(n_1755),
.B(n_1763),
.C(n_1751),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2680),
.Y(n_2904)
);

O2A1O1Ixp5_ASAP7_75t_L g2905 ( 
.A1(n_2879),
.A2(n_1799),
.B(n_1800),
.C(n_1796),
.Y(n_2905)
);

OAI21xp5_ASAP7_75t_L g2906 ( 
.A1(n_2883),
.A2(n_2712),
.B(n_2705),
.Y(n_2906)
);

AO21x1_ASAP7_75t_L g2907 ( 
.A1(n_2700),
.A2(n_2692),
.B(n_2716),
.Y(n_2907)
);

INVx4_ASAP7_75t_L g2908 ( 
.A(n_2882),
.Y(n_2908)
);

NAND2x1p5_ASAP7_75t_L g2909 ( 
.A(n_2864),
.B(n_1805),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2695),
.B(n_1868),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2858),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_SL g2912 ( 
.A(n_2710),
.B(n_1869),
.Y(n_2912)
);

HB1xp67_ASAP7_75t_L g2913 ( 
.A(n_2728),
.Y(n_2913)
);

AOI21xp5_ASAP7_75t_L g2914 ( 
.A1(n_2773),
.A2(n_1818),
.B(n_1817),
.Y(n_2914)
);

AOI21xp5_ASAP7_75t_L g2915 ( 
.A1(n_2793),
.A2(n_1834),
.B(n_1827),
.Y(n_2915)
);

AND2x2_ASAP7_75t_L g2916 ( 
.A(n_2721),
.B(n_1873),
.Y(n_2916)
);

A2O1A1Ixp33_ASAP7_75t_L g2917 ( 
.A1(n_2778),
.A2(n_1843),
.B(n_1853),
.C(n_1837),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2697),
.B(n_1874),
.Y(n_2918)
);

AO21x1_ASAP7_75t_L g2919 ( 
.A1(n_2747),
.A2(n_1856),
.B(n_1855),
.Y(n_2919)
);

AOI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2696),
.A2(n_1866),
.B(n_1864),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_SL g2921 ( 
.A(n_2851),
.B(n_2852),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_SL g2922 ( 
.A(n_2856),
.B(n_1878),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_SL g2923 ( 
.A(n_2860),
.B(n_1880),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2702),
.Y(n_2924)
);

AOI21xp5_ASAP7_75t_L g2925 ( 
.A1(n_2855),
.A2(n_1876),
.B(n_1875),
.Y(n_2925)
);

AOI21xp5_ASAP7_75t_L g2926 ( 
.A1(n_2857),
.A2(n_2873),
.B(n_2871),
.Y(n_2926)
);

AOI21x1_ASAP7_75t_L g2927 ( 
.A1(n_2866),
.A2(n_1885),
.B(n_1881),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2698),
.B(n_1883),
.Y(n_2928)
);

NOR2xp33_ASAP7_75t_L g2929 ( 
.A(n_2719),
.B(n_1884),
.Y(n_2929)
);

AOI21x1_ASAP7_75t_L g2930 ( 
.A1(n_2868),
.A2(n_1900),
.B(n_1899),
.Y(n_2930)
);

BUFx8_ASAP7_75t_L g2931 ( 
.A(n_2800),
.Y(n_2931)
);

NOR3xp33_ASAP7_75t_L g2932 ( 
.A(n_2750),
.B(n_1892),
.C(n_1891),
.Y(n_2932)
);

NOR2xp33_ASAP7_75t_L g2933 ( 
.A(n_2726),
.B(n_1893),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_SL g2934 ( 
.A(n_2876),
.B(n_1896),
.Y(n_2934)
);

AOI21xp5_ASAP7_75t_L g2935 ( 
.A1(n_2802),
.A2(n_1908),
.B(n_1905),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2878),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2722),
.B(n_1897),
.Y(n_2937)
);

AOI21xp5_ASAP7_75t_L g2938 ( 
.A1(n_2880),
.A2(n_1911),
.B(n_1909),
.Y(n_2938)
);

HB1xp67_ASAP7_75t_L g2939 ( 
.A(n_2729),
.Y(n_2939)
);

NOR2xp33_ASAP7_75t_L g2940 ( 
.A(n_2758),
.B(n_1898),
.Y(n_2940)
);

AND2x4_ASAP7_75t_L g2941 ( 
.A(n_2872),
.B(n_1929),
.Y(n_2941)
);

A2O1A1Ixp33_ASAP7_75t_L g2942 ( 
.A1(n_2808),
.A2(n_1947),
.B(n_1948),
.C(n_1946),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2725),
.B(n_1902),
.Y(n_2943)
);

AOI21x1_ASAP7_75t_L g2944 ( 
.A1(n_2741),
.A2(n_1958),
.B(n_1953),
.Y(n_2944)
);

OAI21xp5_ASAP7_75t_L g2945 ( 
.A1(n_2881),
.A2(n_1961),
.B(n_1960),
.Y(n_2945)
);

AOI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_2688),
.A2(n_2854),
.B(n_2703),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2859),
.B(n_1903),
.Y(n_2947)
);

AOI21x1_ASAP7_75t_L g2948 ( 
.A1(n_2737),
.A2(n_1981),
.B(n_1976),
.Y(n_2948)
);

OR2x2_ASAP7_75t_L g2949 ( 
.A(n_2731),
.B(n_2732),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2862),
.B(n_1906),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2863),
.B(n_1910),
.Y(n_2951)
);

AO21x1_ASAP7_75t_L g2952 ( 
.A1(n_2691),
.A2(n_1986),
.B(n_1984),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2718),
.Y(n_2953)
);

AOI21xp33_ASAP7_75t_L g2954 ( 
.A1(n_2686),
.A2(n_1915),
.B(n_1914),
.Y(n_2954)
);

O2A1O1Ixp33_ASAP7_75t_L g2955 ( 
.A1(n_2832),
.A2(n_1991),
.B(n_1992),
.C(n_1988),
.Y(n_2955)
);

AOI21xp5_ASAP7_75t_L g2956 ( 
.A1(n_2854),
.A2(n_2714),
.B(n_2708),
.Y(n_2956)
);

AOI21xp5_ASAP7_75t_L g2957 ( 
.A1(n_2759),
.A2(n_2009),
.B(n_2008),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_L g2958 ( 
.A(n_2709),
.B(n_1919),
.Y(n_2958)
);

AOI21xp5_ASAP7_75t_L g2959 ( 
.A1(n_2690),
.A2(n_2018),
.B(n_2010),
.Y(n_2959)
);

AOI22xp33_ASAP7_75t_L g2960 ( 
.A1(n_2707),
.A2(n_2028),
.B1(n_2030),
.B2(n_2027),
.Y(n_2960)
);

AND2x6_ASAP7_75t_L g2961 ( 
.A(n_2754),
.B(n_2037),
.Y(n_2961)
);

AOI21x1_ASAP7_75t_L g2962 ( 
.A1(n_2739),
.A2(n_2046),
.B(n_2045),
.Y(n_2962)
);

NAND2x1p5_ASAP7_75t_L g2963 ( 
.A(n_2729),
.B(n_330),
.Y(n_2963)
);

OR2x6_ASAP7_75t_SL g2964 ( 
.A(n_2811),
.B(n_1922),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2684),
.B(n_1924),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2685),
.B(n_1926),
.Y(n_2966)
);

O2A1O1Ixp5_ASAP7_75t_L g2967 ( 
.A1(n_2720),
.A2(n_1932),
.B(n_1933),
.C(n_1930),
.Y(n_2967)
);

BUFx4f_ASAP7_75t_L g2968 ( 
.A(n_2850),
.Y(n_2968)
);

A2O1A1Ixp33_ASAP7_75t_L g2969 ( 
.A1(n_2814),
.A2(n_1935),
.B(n_1936),
.C(n_1934),
.Y(n_2969)
);

AOI21xp5_ASAP7_75t_L g2970 ( 
.A1(n_2735),
.A2(n_1940),
.B(n_1939),
.Y(n_2970)
);

OAI21xp5_ASAP7_75t_L g2971 ( 
.A1(n_2736),
.A2(n_2733),
.B(n_2727),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2699),
.B(n_1941),
.Y(n_2972)
);

AOI21xp5_ASAP7_75t_L g2973 ( 
.A1(n_2761),
.A2(n_1944),
.B(n_1942),
.Y(n_2973)
);

AOI21xp5_ASAP7_75t_L g2974 ( 
.A1(n_2740),
.A2(n_1950),
.B(n_1949),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2701),
.B(n_1951),
.Y(n_2975)
);

BUFx6f_ASAP7_75t_L g2976 ( 
.A(n_2782),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2748),
.B(n_1954),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2779),
.B(n_1957),
.Y(n_2978)
);

AOI22xp5_ASAP7_75t_L g2979 ( 
.A1(n_2723),
.A2(n_1965),
.B1(n_1968),
.B2(n_1962),
.Y(n_2979)
);

NAND3xp33_ASAP7_75t_L g2980 ( 
.A(n_2694),
.B(n_1970),
.C(n_1969),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2787),
.Y(n_2981)
);

AOI21xp5_ASAP7_75t_L g2982 ( 
.A1(n_2730),
.A2(n_1972),
.B(n_1971),
.Y(n_2982)
);

OAI22xp5_ASAP7_75t_L g2983 ( 
.A1(n_2780),
.A2(n_1978),
.B1(n_1985),
.B2(n_1975),
.Y(n_2983)
);

OAI22xp33_ASAP7_75t_L g2984 ( 
.A1(n_2861),
.A2(n_1989),
.B1(n_1990),
.B2(n_1987),
.Y(n_2984)
);

AOI21xp5_ASAP7_75t_L g2985 ( 
.A1(n_2744),
.A2(n_1995),
.B(n_1993),
.Y(n_2985)
);

AND2x2_ASAP7_75t_L g2986 ( 
.A(n_2724),
.B(n_1996),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2788),
.Y(n_2987)
);

BUFx2_ASAP7_75t_SL g2988 ( 
.A(n_2837),
.Y(n_2988)
);

AOI21xp5_ASAP7_75t_L g2989 ( 
.A1(n_2746),
.A2(n_1999),
.B(n_1997),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2791),
.Y(n_2990)
);

AOI21xp5_ASAP7_75t_L g2991 ( 
.A1(n_2751),
.A2(n_2004),
.B(n_2003),
.Y(n_2991)
);

NOR2xp33_ASAP7_75t_L g2992 ( 
.A(n_2822),
.B(n_2818),
.Y(n_2992)
);

NOR2xp33_ASAP7_75t_L g2993 ( 
.A(n_2842),
.B(n_2005),
.Y(n_2993)
);

OAI22xp5_ASAP7_75t_L g2994 ( 
.A1(n_2799),
.A2(n_2007),
.B1(n_2011),
.B2(n_2006),
.Y(n_2994)
);

O2A1O1Ixp33_ASAP7_75t_L g2995 ( 
.A1(n_2760),
.A2(n_2016),
.B(n_2017),
.C(n_2014),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2792),
.Y(n_2996)
);

CKINVDCx10_ASAP7_75t_R g2997 ( 
.A(n_2834),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2770),
.B(n_2021),
.Y(n_2998)
);

AO21x1_ASAP7_75t_L g2999 ( 
.A1(n_2785),
.A2(n_332),
.B(n_331),
.Y(n_2999)
);

OAI22xp5_ASAP7_75t_L g3000 ( 
.A1(n_2713),
.A2(n_2023),
.B1(n_2024),
.B2(n_2022),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2771),
.B(n_2025),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2687),
.B(n_2033),
.Y(n_3002)
);

AOI21xp5_ASAP7_75t_L g3003 ( 
.A1(n_2753),
.A2(n_2038),
.B(n_2036),
.Y(n_3003)
);

HB1xp67_ASAP7_75t_L g3004 ( 
.A(n_2828),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_SL g3005 ( 
.A(n_2796),
.B(n_2039),
.Y(n_3005)
);

NOR2xp33_ASAP7_75t_L g3006 ( 
.A(n_2752),
.B(n_2041),
.Y(n_3006)
);

OAI21xp5_ASAP7_75t_L g3007 ( 
.A1(n_2757),
.A2(n_2044),
.B(n_2043),
.Y(n_3007)
);

AO22x1_ASAP7_75t_L g3008 ( 
.A1(n_2843),
.A2(n_2052),
.B1(n_2053),
.B2(n_2051),
.Y(n_3008)
);

NAND3xp33_ASAP7_75t_L g3009 ( 
.A(n_2776),
.B(n_0),
.C(n_1),
.Y(n_3009)
);

NAND2x1p5_ASAP7_75t_L g3010 ( 
.A(n_2749),
.B(n_333),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_SL g3011 ( 
.A(n_2797),
.B(n_2805),
.Y(n_3011)
);

BUFx6f_ASAP7_75t_L g3012 ( 
.A(n_2830),
.Y(n_3012)
);

A2O1A1Ixp33_ASAP7_75t_L g3013 ( 
.A1(n_2795),
.A2(n_3),
.B(n_1),
.C(n_2),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2806),
.Y(n_3014)
);

NOR2xp67_ASAP7_75t_L g3015 ( 
.A(n_2845),
.B(n_2),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_SL g3016 ( 
.A(n_2839),
.B(n_336),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2707),
.B(n_2756),
.Y(n_3017)
);

NOR2xp33_ASAP7_75t_L g3018 ( 
.A(n_2813),
.B(n_339),
.Y(n_3018)
);

A2O1A1Ixp33_ASAP7_75t_L g3019 ( 
.A1(n_2784),
.A2(n_4),
.B(n_2),
.C(n_3),
.Y(n_3019)
);

OAI22xp5_ASAP7_75t_L g3020 ( 
.A1(n_2766),
.A2(n_341),
.B1(n_342),
.B2(n_340),
.Y(n_3020)
);

AOI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2812),
.A2(n_343),
.B(n_340),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2816),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2707),
.B(n_4),
.Y(n_3023)
);

AND2x2_ASAP7_75t_L g3024 ( 
.A(n_2836),
.B(n_344),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2786),
.B(n_4),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2743),
.Y(n_3026)
);

AOI21xp5_ASAP7_75t_L g3027 ( 
.A1(n_2817),
.A2(n_346),
.B(n_345),
.Y(n_3027)
);

BUFx6f_ASAP7_75t_L g3028 ( 
.A(n_2715),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2804),
.B(n_5),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2819),
.B(n_6),
.Y(n_3030)
);

AOI21xp5_ASAP7_75t_L g3031 ( 
.A1(n_2827),
.A2(n_346),
.B(n_345),
.Y(n_3031)
);

AOI22xp5_ASAP7_75t_L g3032 ( 
.A1(n_2794),
.A2(n_349),
.B1(n_350),
.B2(n_348),
.Y(n_3032)
);

NOR2xp33_ASAP7_75t_L g3033 ( 
.A(n_2798),
.B(n_348),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_2831),
.B(n_7),
.Y(n_3034)
);

BUFx6f_ASAP7_75t_L g3035 ( 
.A(n_2717),
.Y(n_3035)
);

AOI21xp5_ASAP7_75t_L g3036 ( 
.A1(n_2738),
.A2(n_352),
.B(n_351),
.Y(n_3036)
);

INVxp67_ASAP7_75t_L g3037 ( 
.A(n_2833),
.Y(n_3037)
);

BUFx8_ASAP7_75t_SL g3038 ( 
.A(n_2834),
.Y(n_3038)
);

OAI21x1_ASAP7_75t_L g3039 ( 
.A1(n_2820),
.A2(n_353),
.B(n_351),
.Y(n_3039)
);

OAI22xp5_ASAP7_75t_L g3040 ( 
.A1(n_2826),
.A2(n_354),
.B1(n_355),
.B2(n_353),
.Y(n_3040)
);

O2A1O1Ixp33_ASAP7_75t_L g3041 ( 
.A1(n_2742),
.A2(n_355),
.B(n_356),
.C(n_354),
.Y(n_3041)
);

AOI22x1_ASAP7_75t_L g3042 ( 
.A1(n_2824),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_3042)
);

OAI21xp33_ASAP7_75t_L g3043 ( 
.A1(n_2772),
.A2(n_8),
.B(n_9),
.Y(n_3043)
);

AOI21xp5_ASAP7_75t_L g3044 ( 
.A1(n_2765),
.A2(n_358),
.B(n_357),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2869),
.B(n_9),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_SL g3046 ( 
.A(n_2840),
.B(n_2789),
.Y(n_3046)
);

AOI21xp5_ASAP7_75t_L g3047 ( 
.A1(n_2767),
.A2(n_2769),
.B(n_2768),
.Y(n_3047)
);

AOI21xp5_ASAP7_75t_L g3048 ( 
.A1(n_2777),
.A2(n_2774),
.B(n_2790),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2849),
.B(n_10),
.Y(n_3049)
);

NOR2x1p5_ASAP7_75t_L g3050 ( 
.A(n_2848),
.B(n_2775),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2734),
.B(n_10),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2904),
.Y(n_3052)
);

NOR2xp33_ASAP7_75t_R g3053 ( 
.A(n_2889),
.B(n_2853),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2924),
.Y(n_3054)
);

BUFx6f_ASAP7_75t_L g3055 ( 
.A(n_3028),
.Y(n_3055)
);

OR2x6_ASAP7_75t_L g3056 ( 
.A(n_2988),
.B(n_2874),
.Y(n_3056)
);

A2O1A1Ixp33_ASAP7_75t_L g3057 ( 
.A1(n_2940),
.A2(n_2781),
.B(n_2838),
.C(n_2847),
.Y(n_3057)
);

AOI21xp33_ASAP7_75t_L g3058 ( 
.A1(n_2896),
.A2(n_2755),
.B(n_2825),
.Y(n_3058)
);

NOR2xp33_ASAP7_75t_L g3059 ( 
.A(n_2898),
.B(n_2809),
.Y(n_3059)
);

A2O1A1Ixp33_ASAP7_75t_L g3060 ( 
.A1(n_2929),
.A2(n_2829),
.B(n_2815),
.C(n_2810),
.Y(n_3060)
);

AOI21xp5_ASAP7_75t_L g3061 ( 
.A1(n_2921),
.A2(n_2835),
.B(n_2844),
.Y(n_3061)
);

A2O1A1Ixp33_ASAP7_75t_L g3062 ( 
.A1(n_2933),
.A2(n_2821),
.B(n_2764),
.C(n_2841),
.Y(n_3062)
);

O2A1O1Ixp33_ASAP7_75t_L g3063 ( 
.A1(n_3049),
.A2(n_2783),
.B(n_2803),
.C(n_2693),
.Y(n_3063)
);

HB1xp67_ASAP7_75t_L g3064 ( 
.A(n_2891),
.Y(n_3064)
);

INVx5_ASAP7_75t_L g3065 ( 
.A(n_3038),
.Y(n_3065)
);

CKINVDCx20_ASAP7_75t_R g3066 ( 
.A(n_2931),
.Y(n_3066)
);

OR2x6_ASAP7_75t_L g3067 ( 
.A(n_2884),
.B(n_2807),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2949),
.B(n_11),
.Y(n_3068)
);

OAI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_2971),
.A2(n_12),
.B(n_14),
.Y(n_3069)
);

CKINVDCx5p33_ASAP7_75t_R g3070 ( 
.A(n_2997),
.Y(n_3070)
);

NOR2xp33_ASAP7_75t_L g3071 ( 
.A(n_2892),
.B(n_360),
.Y(n_3071)
);

AOI22xp33_ASAP7_75t_L g3072 ( 
.A1(n_2907),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2895),
.B(n_16),
.Y(n_3073)
);

INVxp67_ASAP7_75t_L g3074 ( 
.A(n_2913),
.Y(n_3074)
);

AOI21x1_ASAP7_75t_L g3075 ( 
.A1(n_2926),
.A2(n_362),
.B(n_361),
.Y(n_3075)
);

AOI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_3046),
.A2(n_364),
.B(n_363),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_2899),
.B(n_17),
.Y(n_3077)
);

NOR2xp33_ASAP7_75t_L g3078 ( 
.A(n_2900),
.B(n_364),
.Y(n_3078)
);

INVx3_ASAP7_75t_L g3079 ( 
.A(n_2908),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2894),
.B(n_17),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2993),
.B(n_18),
.Y(n_3081)
);

BUFx2_ASAP7_75t_L g3082 ( 
.A(n_2939),
.Y(n_3082)
);

AOI22xp5_ASAP7_75t_L g3083 ( 
.A1(n_2932),
.A2(n_367),
.B1(n_368),
.B2(n_366),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_SL g3084 ( 
.A(n_3037),
.B(n_3006),
.Y(n_3084)
);

INVx4_ASAP7_75t_L g3085 ( 
.A(n_2976),
.Y(n_3085)
);

AND2x4_ASAP7_75t_L g3086 ( 
.A(n_3028),
.B(n_366),
.Y(n_3086)
);

INVx5_ASAP7_75t_L g3087 ( 
.A(n_3035),
.Y(n_3087)
);

AND2x2_ASAP7_75t_L g3088 ( 
.A(n_2893),
.B(n_369),
.Y(n_3088)
);

OAI21x1_ASAP7_75t_L g3089 ( 
.A1(n_2927),
.A2(n_18),
.B(n_19),
.Y(n_3089)
);

OAI22x1_ASAP7_75t_L g3090 ( 
.A1(n_3042),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_3090)
);

AO21x2_ASAP7_75t_L g3091 ( 
.A1(n_2956),
.A2(n_21),
.B(n_22),
.Y(n_3091)
);

BUFx12f_ASAP7_75t_L g3092 ( 
.A(n_2888),
.Y(n_3092)
);

AOI21xp5_ASAP7_75t_L g3093 ( 
.A1(n_3011),
.A2(n_372),
.B(n_370),
.Y(n_3093)
);

AO32x1_ASAP7_75t_L g3094 ( 
.A1(n_3040),
.A2(n_24),
.A3(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_3094)
);

AOI21xp5_ASAP7_75t_L g3095 ( 
.A1(n_2946),
.A2(n_374),
.B(n_373),
.Y(n_3095)
);

BUFx6f_ASAP7_75t_L g3096 ( 
.A(n_2976),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2996),
.Y(n_3097)
);

BUFx3_ASAP7_75t_L g3098 ( 
.A(n_2976),
.Y(n_3098)
);

OR2x6_ASAP7_75t_L g3099 ( 
.A(n_2888),
.B(n_374),
.Y(n_3099)
);

INVx3_ASAP7_75t_L g3100 ( 
.A(n_3012),
.Y(n_3100)
);

NOR2xp33_ASAP7_75t_L g3101 ( 
.A(n_2977),
.B(n_375),
.Y(n_3101)
);

INVxp67_ASAP7_75t_L g3102 ( 
.A(n_3004),
.Y(n_3102)
);

INVx8_ASAP7_75t_L g3103 ( 
.A(n_3012),
.Y(n_3103)
);

O2A1O1Ixp33_ASAP7_75t_SL g3104 ( 
.A1(n_3013),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2910),
.B(n_24),
.Y(n_3105)
);

OAI21xp5_ASAP7_75t_L g3106 ( 
.A1(n_2945),
.A2(n_26),
.B(n_27),
.Y(n_3106)
);

AOI21xp5_ASAP7_75t_L g3107 ( 
.A1(n_3048),
.A2(n_377),
.B(n_376),
.Y(n_3107)
);

OAI22xp5_ASAP7_75t_SL g3108 ( 
.A1(n_3033),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_3108)
);

OAI21x1_ASAP7_75t_L g3109 ( 
.A1(n_2930),
.A2(n_27),
.B(n_29),
.Y(n_3109)
);

BUFx6f_ASAP7_75t_L g3110 ( 
.A(n_3012),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_2953),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_2981),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2918),
.B(n_29),
.Y(n_3113)
);

AOI21xp5_ASAP7_75t_L g3114 ( 
.A1(n_3047),
.A2(n_379),
.B(n_378),
.Y(n_3114)
);

AOI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_2928),
.A2(n_380),
.B(n_379),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2958),
.B(n_30),
.Y(n_3116)
);

OAI21x1_ASAP7_75t_L g3117 ( 
.A1(n_2948),
.A2(n_31),
.B(n_32),
.Y(n_3117)
);

INVx2_ASAP7_75t_L g3118 ( 
.A(n_2987),
.Y(n_3118)
);

OAI22xp5_ASAP7_75t_L g3119 ( 
.A1(n_2972),
.A2(n_384),
.B1(n_385),
.B2(n_381),
.Y(n_3119)
);

INVx2_ASAP7_75t_SL g3120 ( 
.A(n_2941),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2965),
.B(n_31),
.Y(n_3121)
);

OAI21xp33_ASAP7_75t_SL g3122 ( 
.A1(n_3051),
.A2(n_3016),
.B(n_3030),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_2966),
.B(n_33),
.Y(n_3123)
);

NOR3xp33_ASAP7_75t_SL g3124 ( 
.A(n_3009),
.B(n_33),
.C(n_34),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2990),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2886),
.Y(n_3126)
);

OAI22xp5_ASAP7_75t_L g3127 ( 
.A1(n_2975),
.A2(n_387),
.B1(n_388),
.B2(n_386),
.Y(n_3127)
);

O2A1O1Ixp33_ASAP7_75t_L g3128 ( 
.A1(n_3019),
.A2(n_387),
.B(n_389),
.C(n_386),
.Y(n_3128)
);

NOR3xp33_ASAP7_75t_SL g3129 ( 
.A(n_2984),
.B(n_34),
.C(n_35),
.Y(n_3129)
);

OAI22xp5_ASAP7_75t_L g3130 ( 
.A1(n_2998),
.A2(n_392),
.B1(n_393),
.B2(n_390),
.Y(n_3130)
);

AOI21xp5_ASAP7_75t_L g3131 ( 
.A1(n_3005),
.A2(n_2923),
.B(n_2922),
.Y(n_3131)
);

OAI22xp5_ASAP7_75t_L g3132 ( 
.A1(n_3001),
.A2(n_395),
.B1(n_396),
.B2(n_394),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2911),
.Y(n_3133)
);

CKINVDCx11_ASAP7_75t_R g3134 ( 
.A(n_2964),
.Y(n_3134)
);

BUFx3_ASAP7_75t_L g3135 ( 
.A(n_3026),
.Y(n_3135)
);

NOR2xp33_ASAP7_75t_R g3136 ( 
.A(n_2962),
.B(n_398),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_SL g3137 ( 
.A(n_3024),
.B(n_399),
.Y(n_3137)
);

AOI22xp33_ASAP7_75t_L g3138 ( 
.A1(n_3018),
.A2(n_3043),
.B1(n_2980),
.B2(n_2954),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2936),
.Y(n_3139)
);

AOI22xp5_ASAP7_75t_L g3140 ( 
.A1(n_3050),
.A2(n_401),
.B1(n_402),
.B2(n_400),
.Y(n_3140)
);

O2A1O1Ixp33_ASAP7_75t_L g3141 ( 
.A1(n_2942),
.A2(n_2903),
.B(n_2969),
.C(n_2917),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_3014),
.Y(n_3142)
);

OAI22xp5_ASAP7_75t_L g3143 ( 
.A1(n_3022),
.A2(n_403),
.B1(n_404),
.B2(n_401),
.Y(n_3143)
);

AOI21xp5_ASAP7_75t_L g3144 ( 
.A1(n_2934),
.A2(n_406),
.B(n_405),
.Y(n_3144)
);

AOI21xp5_ASAP7_75t_L g3145 ( 
.A1(n_2912),
.A2(n_408),
.B(n_407),
.Y(n_3145)
);

A2O1A1Ixp33_ASAP7_75t_L g3146 ( 
.A1(n_2995),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_3146)
);

O2A1O1Ixp33_ASAP7_75t_SL g3147 ( 
.A1(n_3017),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_3147)
);

NOR2xp33_ASAP7_75t_L g3148 ( 
.A(n_2986),
.B(n_408),
.Y(n_3148)
);

O2A1O1Ixp33_ASAP7_75t_L g3149 ( 
.A1(n_3034),
.A2(n_410),
.B(n_411),
.C(n_409),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_2944),
.Y(n_3150)
);

AND2x6_ASAP7_75t_L g3151 ( 
.A(n_3032),
.B(n_40),
.Y(n_3151)
);

OAI21xp5_ASAP7_75t_L g3152 ( 
.A1(n_2967),
.A2(n_41),
.B(n_42),
.Y(n_3152)
);

A2O1A1Ixp33_ASAP7_75t_L g3153 ( 
.A1(n_2905),
.A2(n_44),
.B(n_41),
.C(n_43),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_3025),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_SL g3155 ( 
.A(n_2916),
.B(n_409),
.Y(n_3155)
);

A2O1A1Ixp33_ASAP7_75t_L g3156 ( 
.A1(n_3031),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2937),
.Y(n_3157)
);

CKINVDCx5p33_ASAP7_75t_R g3158 ( 
.A(n_3008),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2943),
.B(n_44),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2947),
.B(n_45),
.Y(n_3160)
);

CKINVDCx5p33_ASAP7_75t_R g3161 ( 
.A(n_2890),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2950),
.B(n_45),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_3007),
.B(n_412),
.Y(n_3163)
);

A2O1A1Ixp33_ASAP7_75t_L g3164 ( 
.A1(n_2897),
.A2(n_48),
.B(n_46),
.C(n_47),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_2952),
.B(n_413),
.Y(n_3165)
);

NOR2xp67_ASAP7_75t_SL g3166 ( 
.A(n_3045),
.B(n_46),
.Y(n_3166)
);

CKINVDCx5p33_ASAP7_75t_R g3167 ( 
.A(n_2994),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2951),
.B(n_46),
.Y(n_3168)
);

INVx4_ASAP7_75t_L g3169 ( 
.A(n_2961),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_SL g3170 ( 
.A(n_3015),
.B(n_414),
.Y(n_3170)
);

BUFx3_ASAP7_75t_L g3171 ( 
.A(n_2909),
.Y(n_3171)
);

AOI22x1_ASAP7_75t_L g3172 ( 
.A1(n_2915),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_3172)
);

BUFx3_ASAP7_75t_L g3173 ( 
.A(n_3010),
.Y(n_3173)
);

AND2x6_ASAP7_75t_L g3174 ( 
.A(n_3023),
.B(n_47),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_SL g3175 ( 
.A(n_2979),
.B(n_3029),
.Y(n_3175)
);

INVx2_ASAP7_75t_SL g3176 ( 
.A(n_2963),
.Y(n_3176)
);

O2A1O1Ixp33_ASAP7_75t_L g3177 ( 
.A1(n_3020),
.A2(n_416),
.B(n_417),
.C(n_415),
.Y(n_3177)
);

NOR3xp33_ASAP7_75t_SL g3178 ( 
.A(n_3000),
.B(n_51),
.C(n_52),
.Y(n_3178)
);

OAI22xp5_ASAP7_75t_L g3179 ( 
.A1(n_2978),
.A2(n_418),
.B1(n_419),
.B2(n_416),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_2901),
.B(n_51),
.Y(n_3180)
);

AND2x2_ASAP7_75t_L g3181 ( 
.A(n_3002),
.B(n_420),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_SL g3182 ( 
.A(n_2982),
.B(n_421),
.Y(n_3182)
);

OAI21x1_ASAP7_75t_L g3183 ( 
.A1(n_3039),
.A2(n_52),
.B(n_53),
.Y(n_3183)
);

O2A1O1Ixp33_ASAP7_75t_L g3184 ( 
.A1(n_3041),
.A2(n_423),
.B(n_424),
.C(n_422),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_2920),
.B(n_53),
.Y(n_3185)
);

INVx2_ASAP7_75t_SL g3186 ( 
.A(n_2961),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2919),
.Y(n_3187)
);

NOR2xp33_ASAP7_75t_SL g3188 ( 
.A(n_3044),
.B(n_53),
.Y(n_3188)
);

OR2x2_ASAP7_75t_L g3189 ( 
.A(n_2983),
.B(n_54),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_2960),
.B(n_425),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_SL g3191 ( 
.A(n_2991),
.B(n_427),
.Y(n_3191)
);

AOI21xp5_ASAP7_75t_L g3192 ( 
.A1(n_2902),
.A2(n_431),
.B(n_428),
.Y(n_3192)
);

BUFx12f_ASAP7_75t_L g3193 ( 
.A(n_2999),
.Y(n_3193)
);

AOI21xp5_ASAP7_75t_L g3194 ( 
.A1(n_2935),
.A2(n_432),
.B(n_428),
.Y(n_3194)
);

AND2x2_ASAP7_75t_L g3195 ( 
.A(n_2885),
.B(n_432),
.Y(n_3195)
);

HB1xp67_ASAP7_75t_L g3196 ( 
.A(n_2938),
.Y(n_3196)
);

A2O1A1Ixp33_ASAP7_75t_L g3197 ( 
.A1(n_3021),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_3197)
);

A2O1A1Ixp33_ASAP7_75t_L g3198 ( 
.A1(n_3027),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_3198)
);

CKINVDCx5p33_ASAP7_75t_R g3199 ( 
.A(n_2914),
.Y(n_3199)
);

BUFx12f_ASAP7_75t_SL g3200 ( 
.A(n_2959),
.Y(n_3200)
);

AOI21xp5_ASAP7_75t_L g3201 ( 
.A1(n_2973),
.A2(n_434),
.B(n_433),
.Y(n_3201)
);

NOR2xp33_ASAP7_75t_L g3202 ( 
.A(n_3003),
.B(n_435),
.Y(n_3202)
);

OAI22xp5_ASAP7_75t_L g3203 ( 
.A1(n_2974),
.A2(n_436),
.B1(n_437),
.B2(n_435),
.Y(n_3203)
);

INVx3_ASAP7_75t_L g3204 ( 
.A(n_3036),
.Y(n_3204)
);

BUFx10_ASAP7_75t_L g3205 ( 
.A(n_2985),
.Y(n_3205)
);

OR2x2_ASAP7_75t_L g3206 ( 
.A(n_2989),
.B(n_57),
.Y(n_3206)
);

OR2x6_ASAP7_75t_L g3207 ( 
.A(n_2955),
.B(n_437),
.Y(n_3207)
);

BUFx6f_ASAP7_75t_L g3208 ( 
.A(n_2925),
.Y(n_3208)
);

NOR2xp33_ASAP7_75t_L g3209 ( 
.A(n_2970),
.B(n_438),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_SL g3210 ( 
.A(n_2957),
.B(n_439),
.Y(n_3210)
);

INVx1_ASAP7_75t_SL g3211 ( 
.A(n_2891),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_SL g3212 ( 
.A(n_2992),
.B(n_441),
.Y(n_3212)
);

OAI21xp5_ASAP7_75t_L g3213 ( 
.A1(n_2906),
.A2(n_59),
.B(n_60),
.Y(n_3213)
);

BUFx6f_ASAP7_75t_L g3214 ( 
.A(n_2968),
.Y(n_3214)
);

NAND2x1p5_ASAP7_75t_L g3215 ( 
.A(n_2887),
.B(n_442),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2904),
.Y(n_3216)
);

NAND2xp33_ASAP7_75t_L g3217 ( 
.A(n_2906),
.B(n_62),
.Y(n_3217)
);

NOR2x1_ASAP7_75t_L g3218 ( 
.A(n_2887),
.B(n_443),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_3157),
.B(n_63),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_3154),
.B(n_64),
.Y(n_3220)
);

AOI21xp33_ASAP7_75t_L g3221 ( 
.A1(n_3059),
.A2(n_65),
.B(n_66),
.Y(n_3221)
);

INVx3_ASAP7_75t_L g3222 ( 
.A(n_3087),
.Y(n_3222)
);

CKINVDCx20_ASAP7_75t_R g3223 ( 
.A(n_3066),
.Y(n_3223)
);

AOI21xp5_ASAP7_75t_L g3224 ( 
.A1(n_3217),
.A2(n_446),
.B(n_445),
.Y(n_3224)
);

INVx3_ASAP7_75t_L g3225 ( 
.A(n_3087),
.Y(n_3225)
);

AND2x4_ASAP7_75t_L g3226 ( 
.A(n_3098),
.B(n_449),
.Y(n_3226)
);

BUFx2_ASAP7_75t_SL g3227 ( 
.A(n_3214),
.Y(n_3227)
);

OAI21xp5_ASAP7_75t_L g3228 ( 
.A1(n_3138),
.A2(n_67),
.B(n_68),
.Y(n_3228)
);

NOR2xp67_ASAP7_75t_L g3229 ( 
.A(n_3074),
.B(n_69),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_3084),
.B(n_69),
.Y(n_3230)
);

AO22x2_ASAP7_75t_L g3231 ( 
.A1(n_3213),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_3068),
.B(n_70),
.Y(n_3232)
);

INVx1_ASAP7_75t_SL g3233 ( 
.A(n_3211),
.Y(n_3233)
);

NOR2xp33_ASAP7_75t_SL g3234 ( 
.A(n_3070),
.B(n_73),
.Y(n_3234)
);

OAI21xp5_ASAP7_75t_L g3235 ( 
.A1(n_3058),
.A2(n_74),
.B(n_75),
.Y(n_3235)
);

INVxp67_ASAP7_75t_SL g3236 ( 
.A(n_3064),
.Y(n_3236)
);

BUFx6f_ASAP7_75t_L g3237 ( 
.A(n_3096),
.Y(n_3237)
);

INVx5_ASAP7_75t_L g3238 ( 
.A(n_3103),
.Y(n_3238)
);

AND2x4_ASAP7_75t_SL g3239 ( 
.A(n_3085),
.B(n_450),
.Y(n_3239)
);

AO32x2_ASAP7_75t_L g3240 ( 
.A1(n_3108),
.A2(n_77),
.A3(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_3240)
);

OAI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_3057),
.A2(n_3122),
.B(n_3081),
.Y(n_3241)
);

BUFx12f_ASAP7_75t_L g3242 ( 
.A(n_3065),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_3071),
.B(n_78),
.Y(n_3243)
);

AOI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_3060),
.A2(n_453),
.B(n_452),
.Y(n_3244)
);

OAI21x1_ASAP7_75t_L g3245 ( 
.A1(n_3183),
.A2(n_78),
.B(n_79),
.Y(n_3245)
);

INVx2_ASAP7_75t_SL g3246 ( 
.A(n_3053),
.Y(n_3246)
);

OAI22xp5_ASAP7_75t_L g3247 ( 
.A1(n_3167),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_3078),
.B(n_80),
.Y(n_3248)
);

AO31x2_ASAP7_75t_L g3249 ( 
.A1(n_3150),
.A2(n_82),
.A3(n_80),
.B(n_81),
.Y(n_3249)
);

INVx1_ASAP7_75t_SL g3250 ( 
.A(n_3082),
.Y(n_3250)
);

AND2x4_ASAP7_75t_L g3251 ( 
.A(n_3120),
.B(n_452),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_3101),
.B(n_82),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3073),
.B(n_3077),
.Y(n_3253)
);

OAI21x1_ASAP7_75t_L g3254 ( 
.A1(n_3075),
.A2(n_84),
.B(n_85),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_3080),
.B(n_86),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_3116),
.B(n_86),
.Y(n_3256)
);

A2O1A1Ixp33_ASAP7_75t_L g3257 ( 
.A1(n_3141),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_3257)
);

AOI21xp5_ASAP7_75t_L g3258 ( 
.A1(n_3131),
.A2(n_456),
.B(n_455),
.Y(n_3258)
);

INVx2_ASAP7_75t_SL g3259 ( 
.A(n_3055),
.Y(n_3259)
);

AO31x2_ASAP7_75t_L g3260 ( 
.A1(n_3187),
.A2(n_91),
.A3(n_87),
.B(n_89),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3052),
.Y(n_3261)
);

OAI21xp5_ASAP7_75t_L g3262 ( 
.A1(n_3175),
.A2(n_3069),
.B(n_3106),
.Y(n_3262)
);

AOI21xp5_ASAP7_75t_L g3263 ( 
.A1(n_3061),
.A2(n_458),
.B(n_457),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3054),
.Y(n_3264)
);

OAI22xp5_ASAP7_75t_L g3265 ( 
.A1(n_3199),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_3265)
);

OAI21x1_ASAP7_75t_L g3266 ( 
.A1(n_3089),
.A2(n_92),
.B(n_93),
.Y(n_3266)
);

AO31x2_ASAP7_75t_L g3267 ( 
.A1(n_3090),
.A2(n_3153),
.A3(n_3107),
.B(n_3114),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3105),
.B(n_3113),
.Y(n_3268)
);

OAI22xp5_ASAP7_75t_L g3269 ( 
.A1(n_3161),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_3269)
);

INVx2_ASAP7_75t_SL g3270 ( 
.A(n_3055),
.Y(n_3270)
);

AO21x2_ASAP7_75t_L g3271 ( 
.A1(n_3152),
.A2(n_94),
.B(n_95),
.Y(n_3271)
);

A2O1A1Ixp33_ASAP7_75t_L g3272 ( 
.A1(n_3202),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_3272)
);

OAI21x1_ASAP7_75t_L g3273 ( 
.A1(n_3109),
.A2(n_96),
.B(n_97),
.Y(n_3273)
);

INVx6_ASAP7_75t_SL g3274 ( 
.A(n_3067),
.Y(n_3274)
);

BUFx4_ASAP7_75t_SL g3275 ( 
.A(n_3099),
.Y(n_3275)
);

OAI21x1_ASAP7_75t_L g3276 ( 
.A1(n_3117),
.A2(n_99),
.B(n_100),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_3121),
.B(n_99),
.Y(n_3277)
);

NAND2x1_ASAP7_75t_L g3278 ( 
.A(n_3204),
.B(n_457),
.Y(n_3278)
);

OAI21x1_ASAP7_75t_L g3279 ( 
.A1(n_3095),
.A2(n_99),
.B(n_100),
.Y(n_3279)
);

A2O1A1Ixp33_ASAP7_75t_L g3280 ( 
.A1(n_3163),
.A2(n_3063),
.B(n_3209),
.C(n_3062),
.Y(n_3280)
);

AOI21xp5_ASAP7_75t_L g3281 ( 
.A1(n_3196),
.A2(n_459),
.B(n_458),
.Y(n_3281)
);

NOR2xp67_ASAP7_75t_L g3282 ( 
.A(n_3079),
.B(n_101),
.Y(n_3282)
);

NOR2x1_ASAP7_75t_SL g3283 ( 
.A(n_3193),
.B(n_460),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3123),
.B(n_102),
.Y(n_3284)
);

NAND3xp33_ASAP7_75t_L g3285 ( 
.A(n_3129),
.B(n_102),
.C(n_103),
.Y(n_3285)
);

NOR2xp67_ASAP7_75t_SL g3286 ( 
.A(n_3092),
.B(n_102),
.Y(n_3286)
);

A2O1A1Ixp33_ASAP7_75t_L g3287 ( 
.A1(n_3148),
.A2(n_3177),
.B(n_3145),
.C(n_3128),
.Y(n_3287)
);

A2O1A1Ixp33_ASAP7_75t_L g3288 ( 
.A1(n_3115),
.A2(n_106),
.B(n_104),
.C(n_105),
.Y(n_3288)
);

AO21x1_ASAP7_75t_L g3289 ( 
.A1(n_3184),
.A2(n_465),
.B(n_464),
.Y(n_3289)
);

OAI21xp5_ASAP7_75t_L g3290 ( 
.A1(n_3076),
.A2(n_105),
.B(n_106),
.Y(n_3290)
);

AND2x2_ASAP7_75t_L g3291 ( 
.A(n_3088),
.B(n_107),
.Y(n_3291)
);

AND2x2_ASAP7_75t_L g3292 ( 
.A(n_3181),
.B(n_107),
.Y(n_3292)
);

AND2x4_ASAP7_75t_L g3293 ( 
.A(n_3056),
.B(n_466),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3159),
.B(n_108),
.Y(n_3294)
);

AOI21xp5_ASAP7_75t_L g3295 ( 
.A1(n_3182),
.A2(n_468),
.B(n_467),
.Y(n_3295)
);

OAI21x1_ASAP7_75t_L g3296 ( 
.A1(n_3191),
.A2(n_109),
.B(n_110),
.Y(n_3296)
);

AND2x2_ASAP7_75t_L g3297 ( 
.A(n_3178),
.B(n_3190),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_3160),
.B(n_109),
.Y(n_3298)
);

AOI21xp5_ASAP7_75t_L g3299 ( 
.A1(n_3188),
.A2(n_468),
.B(n_467),
.Y(n_3299)
);

NOR2xp33_ASAP7_75t_SL g3300 ( 
.A(n_3169),
.B(n_110),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_3162),
.B(n_3168),
.Y(n_3301)
);

OAI22xp5_ASAP7_75t_L g3302 ( 
.A1(n_3135),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_3302)
);

AO31x2_ASAP7_75t_L g3303 ( 
.A1(n_3156),
.A2(n_3197),
.A3(n_3198),
.B(n_3146),
.Y(n_3303)
);

AOI21xp5_ASAP7_75t_L g3304 ( 
.A1(n_3208),
.A2(n_470),
.B(n_469),
.Y(n_3304)
);

CKINVDCx20_ASAP7_75t_R g3305 ( 
.A(n_3134),
.Y(n_3305)
);

OAI21x1_ASAP7_75t_L g3306 ( 
.A1(n_3201),
.A2(n_114),
.B(n_115),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3151),
.B(n_116),
.Y(n_3307)
);

AO31x2_ASAP7_75t_L g3308 ( 
.A1(n_3164),
.A2(n_119),
.A3(n_117),
.B(n_118),
.Y(n_3308)
);

BUFx3_ASAP7_75t_L g3309 ( 
.A(n_3056),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_SL g3310 ( 
.A(n_3158),
.B(n_471),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3111),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_3216),
.Y(n_3312)
);

AOI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_3208),
.A2(n_473),
.B(n_472),
.Y(n_3313)
);

OA21x2_ASAP7_75t_L g3314 ( 
.A1(n_3093),
.A2(n_120),
.B(n_121),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_L g3315 ( 
.A(n_3212),
.B(n_120),
.Y(n_3315)
);

NOR2xp33_ASAP7_75t_L g3316 ( 
.A(n_3102),
.B(n_473),
.Y(n_3316)
);

NOR2xp67_ASAP7_75t_L g3317 ( 
.A(n_3142),
.B(n_121),
.Y(n_3317)
);

AOI21xp5_ASAP7_75t_L g3318 ( 
.A1(n_3210),
.A2(n_3180),
.B(n_3207),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3097),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_3112),
.B(n_122),
.Y(n_3320)
);

AND2x2_ASAP7_75t_L g3321 ( 
.A(n_3195),
.B(n_3124),
.Y(n_3321)
);

OAI22xp5_ASAP7_75t_L g3322 ( 
.A1(n_3140),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_3322)
);

OAI22x1_ASAP7_75t_L g3323 ( 
.A1(n_3083),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_3323)
);

BUFx6f_ASAP7_75t_L g3324 ( 
.A(n_3110),
.Y(n_3324)
);

AOI22xp33_ASAP7_75t_L g3325 ( 
.A1(n_3207),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_3325)
);

AOI211x1_ASAP7_75t_L g3326 ( 
.A1(n_3137),
.A2(n_127),
.B(n_125),
.C(n_126),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3125),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3118),
.B(n_127),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3126),
.Y(n_3329)
);

BUFx6f_ASAP7_75t_L g3330 ( 
.A(n_3110),
.Y(n_3330)
);

CKINVDCx11_ASAP7_75t_R g3331 ( 
.A(n_3099),
.Y(n_3331)
);

BUFx4_ASAP7_75t_SL g3332 ( 
.A(n_3173),
.Y(n_3332)
);

OR2x6_ASAP7_75t_L g3333 ( 
.A(n_3176),
.B(n_475),
.Y(n_3333)
);

AO31x2_ASAP7_75t_L g3334 ( 
.A1(n_3203),
.A2(n_131),
.A3(n_129),
.B(n_130),
.Y(n_3334)
);

INVx3_ASAP7_75t_L g3335 ( 
.A(n_3100),
.Y(n_3335)
);

AOI211x1_ASAP7_75t_L g3336 ( 
.A1(n_3155),
.A2(n_131),
.B(n_129),
.C(n_130),
.Y(n_3336)
);

BUFx6f_ASAP7_75t_L g3337 ( 
.A(n_3171),
.Y(n_3337)
);

OAI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_3072),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_3338)
);

AOI21xp33_ASAP7_75t_L g3339 ( 
.A1(n_3206),
.A2(n_134),
.B(n_135),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3133),
.Y(n_3340)
);

AOI21xp5_ASAP7_75t_L g3341 ( 
.A1(n_3192),
.A2(n_3194),
.B(n_3094),
.Y(n_3341)
);

BUFx2_ASAP7_75t_L g3342 ( 
.A(n_3139),
.Y(n_3342)
);

OAI21x1_ASAP7_75t_L g3343 ( 
.A1(n_3144),
.A2(n_136),
.B(n_137),
.Y(n_3343)
);

AOI21xp5_ASAP7_75t_L g3344 ( 
.A1(n_3094),
.A2(n_476),
.B(n_475),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_3091),
.Y(n_3345)
);

OAI22xp5_ASAP7_75t_L g3346 ( 
.A1(n_3189),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_3346)
);

OA21x2_ASAP7_75t_L g3347 ( 
.A1(n_3165),
.A2(n_140),
.B(n_141),
.Y(n_3347)
);

NAND2x1p5_ASAP7_75t_L g3348 ( 
.A(n_3086),
.B(n_477),
.Y(n_3348)
);

OA21x2_ASAP7_75t_L g3349 ( 
.A1(n_3241),
.A2(n_3172),
.B(n_3185),
.Y(n_3349)
);

NOR2x1_ASAP7_75t_SL g3350 ( 
.A(n_3271),
.B(n_3345),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3261),
.Y(n_3351)
);

AND2x4_ASAP7_75t_L g3352 ( 
.A(n_3309),
.B(n_3186),
.Y(n_3352)
);

OAI21xp5_ASAP7_75t_L g3353 ( 
.A1(n_3244),
.A2(n_3149),
.B(n_3127),
.Y(n_3353)
);

NOR2xp67_ASAP7_75t_L g3354 ( 
.A(n_3246),
.B(n_3170),
.Y(n_3354)
);

HB1xp67_ASAP7_75t_L g3355 ( 
.A(n_3236),
.Y(n_3355)
);

NOR2xp33_ASAP7_75t_L g3356 ( 
.A(n_3233),
.B(n_3215),
.Y(n_3356)
);

AND2x2_ASAP7_75t_L g3357 ( 
.A(n_3321),
.B(n_3218),
.Y(n_3357)
);

O2A1O1Ixp33_ASAP7_75t_L g3358 ( 
.A1(n_3280),
.A2(n_3130),
.B(n_3132),
.C(n_3119),
.Y(n_3358)
);

OR2x6_ASAP7_75t_L g3359 ( 
.A(n_3242),
.B(n_3143),
.Y(n_3359)
);

NAND3xp33_ASAP7_75t_L g3360 ( 
.A(n_3287),
.B(n_3166),
.C(n_3179),
.Y(n_3360)
);

OAI21x1_ASAP7_75t_L g3361 ( 
.A1(n_3254),
.A2(n_3205),
.B(n_3200),
.Y(n_3361)
);

O2A1O1Ixp5_ASAP7_75t_L g3362 ( 
.A1(n_3262),
.A2(n_3104),
.B(n_3147),
.C(n_3136),
.Y(n_3362)
);

OAI21x1_ASAP7_75t_L g3363 ( 
.A1(n_3341),
.A2(n_3276),
.B(n_3245),
.Y(n_3363)
);

AND2x4_ASAP7_75t_L g3364 ( 
.A(n_3250),
.B(n_3174),
.Y(n_3364)
);

OAI21x1_ASAP7_75t_L g3365 ( 
.A1(n_3266),
.A2(n_3174),
.B(n_142),
.Y(n_3365)
);

OAI21x1_ASAP7_75t_L g3366 ( 
.A1(n_3273),
.A2(n_143),
.B(n_144),
.Y(n_3366)
);

BUFx2_ASAP7_75t_R g3367 ( 
.A(n_3227),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3264),
.Y(n_3368)
);

A2O1A1Ixp33_ASAP7_75t_L g3369 ( 
.A1(n_3224),
.A2(n_479),
.B(n_480),
.C(n_478),
.Y(n_3369)
);

AOI21x1_ASAP7_75t_L g3370 ( 
.A1(n_3318),
.A2(n_144),
.B(n_145),
.Y(n_3370)
);

HB1xp67_ASAP7_75t_L g3371 ( 
.A(n_3342),
.Y(n_3371)
);

NOR2xp67_ASAP7_75t_L g3372 ( 
.A(n_3238),
.B(n_146),
.Y(n_3372)
);

OAI21x1_ASAP7_75t_L g3373 ( 
.A1(n_3306),
.A2(n_147),
.B(n_148),
.Y(n_3373)
);

OAI21x1_ASAP7_75t_L g3374 ( 
.A1(n_3279),
.A2(n_147),
.B(n_148),
.Y(n_3374)
);

AO31x2_ASAP7_75t_L g3375 ( 
.A1(n_3289),
.A2(n_150),
.A3(n_148),
.B(n_149),
.Y(n_3375)
);

INVx2_ASAP7_75t_SL g3376 ( 
.A(n_3332),
.Y(n_3376)
);

CKINVDCx5p33_ASAP7_75t_R g3377 ( 
.A(n_3223),
.Y(n_3377)
);

INVx2_ASAP7_75t_L g3378 ( 
.A(n_3311),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3268),
.B(n_3301),
.Y(n_3379)
);

OAI21x1_ASAP7_75t_L g3380 ( 
.A1(n_3263),
.A2(n_151),
.B(n_152),
.Y(n_3380)
);

AO21x2_ASAP7_75t_L g3381 ( 
.A1(n_3235),
.A2(n_153),
.B(n_154),
.Y(n_3381)
);

AOI21x1_ASAP7_75t_L g3382 ( 
.A1(n_3278),
.A2(n_154),
.B(n_155),
.Y(n_3382)
);

AOI22xp33_ASAP7_75t_L g3383 ( 
.A1(n_3228),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_3383)
);

OAI21xp5_ASAP7_75t_L g3384 ( 
.A1(n_3290),
.A2(n_156),
.B(n_157),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3253),
.B(n_3297),
.Y(n_3385)
);

OA21x2_ASAP7_75t_L g3386 ( 
.A1(n_3258),
.A2(n_3281),
.B(n_3257),
.Y(n_3386)
);

OAI22xp5_ASAP7_75t_L g3387 ( 
.A1(n_3285),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_3387)
);

O2A1O1Ixp33_ASAP7_75t_L g3388 ( 
.A1(n_3272),
.A2(n_165),
.B(n_163),
.C(n_164),
.Y(n_3388)
);

AOI22xp33_ASAP7_75t_SL g3389 ( 
.A1(n_3231),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_3389)
);

AOI221x1_ASAP7_75t_L g3390 ( 
.A1(n_3323),
.A2(n_484),
.B1(n_485),
.B2(n_483),
.C(n_482),
.Y(n_3390)
);

AND2x2_ASAP7_75t_L g3391 ( 
.A(n_3292),
.B(n_482),
.Y(n_3391)
);

OAI21x1_ASAP7_75t_L g3392 ( 
.A1(n_3343),
.A2(n_167),
.B(n_168),
.Y(n_3392)
);

OAI21x1_ASAP7_75t_L g3393 ( 
.A1(n_3296),
.A2(n_168),
.B(n_169),
.Y(n_3393)
);

OAI21x1_ASAP7_75t_L g3394 ( 
.A1(n_3319),
.A2(n_169),
.B(n_170),
.Y(n_3394)
);

OAI21x1_ASAP7_75t_L g3395 ( 
.A1(n_3312),
.A2(n_169),
.B(n_170),
.Y(n_3395)
);

OAI21x1_ASAP7_75t_L g3396 ( 
.A1(n_3304),
.A2(n_172),
.B(n_173),
.Y(n_3396)
);

AOI21xp5_ASAP7_75t_L g3397 ( 
.A1(n_3299),
.A2(n_488),
.B(n_487),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3327),
.Y(n_3398)
);

OAI21x1_ASAP7_75t_L g3399 ( 
.A1(n_3313),
.A2(n_174),
.B(n_175),
.Y(n_3399)
);

OAI21xp5_ASAP7_75t_L g3400 ( 
.A1(n_3295),
.A2(n_174),
.B(n_175),
.Y(n_3400)
);

AOI21xp5_ASAP7_75t_L g3401 ( 
.A1(n_3300),
.A2(n_491),
.B(n_490),
.Y(n_3401)
);

OAI21x1_ASAP7_75t_L g3402 ( 
.A1(n_3329),
.A2(n_176),
.B(n_178),
.Y(n_3402)
);

BUFx2_ASAP7_75t_SL g3403 ( 
.A(n_3222),
.Y(n_3403)
);

CKINVDCx16_ASAP7_75t_R g3404 ( 
.A(n_3305),
.Y(n_3404)
);

INVx2_ASAP7_75t_L g3405 ( 
.A(n_3340),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3232),
.B(n_492),
.Y(n_3406)
);

OAI22xp5_ASAP7_75t_L g3407 ( 
.A1(n_3243),
.A2(n_182),
.B1(n_179),
.B2(n_180),
.Y(n_3407)
);

OAI21xp5_ASAP7_75t_L g3408 ( 
.A1(n_3288),
.A2(n_179),
.B(n_180),
.Y(n_3408)
);

OAI21x1_ASAP7_75t_L g3409 ( 
.A1(n_3314),
.A2(n_183),
.B(n_184),
.Y(n_3409)
);

INVx2_ASAP7_75t_L g3410 ( 
.A(n_3335),
.Y(n_3410)
);

AOI21xp33_ASAP7_75t_L g3411 ( 
.A1(n_3248),
.A2(n_186),
.B(n_187),
.Y(n_3411)
);

OAI221xp5_ASAP7_75t_L g3412 ( 
.A1(n_3252),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.C(n_189),
.Y(n_3412)
);

OAI21x1_ASAP7_75t_L g3413 ( 
.A1(n_3320),
.A2(n_189),
.B(n_190),
.Y(n_3413)
);

OAI22xp5_ASAP7_75t_L g3414 ( 
.A1(n_3325),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_3414)
);

NOR2x1_ASAP7_75t_SL g3415 ( 
.A(n_3333),
.B(n_495),
.Y(n_3415)
);

INVx3_ASAP7_75t_L g3416 ( 
.A(n_3337),
.Y(n_3416)
);

AO31x2_ASAP7_75t_L g3417 ( 
.A1(n_3344),
.A2(n_193),
.A3(n_191),
.B(n_192),
.Y(n_3417)
);

OAI21x1_ASAP7_75t_L g3418 ( 
.A1(n_3328),
.A2(n_194),
.B(n_195),
.Y(n_3418)
);

OA21x2_ASAP7_75t_L g3419 ( 
.A1(n_3339),
.A2(n_196),
.B(n_197),
.Y(n_3419)
);

NAND3xp33_ASAP7_75t_L g3420 ( 
.A(n_3221),
.B(n_196),
.C(n_197),
.Y(n_3420)
);

AOI21x1_ASAP7_75t_L g3421 ( 
.A1(n_3255),
.A2(n_196),
.B(n_198),
.Y(n_3421)
);

BUFx6f_ASAP7_75t_L g3422 ( 
.A(n_3237),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_3220),
.B(n_497),
.Y(n_3423)
);

AOI22xp5_ASAP7_75t_L g3424 ( 
.A1(n_3322),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_3424)
);

AO31x2_ASAP7_75t_L g3425 ( 
.A1(n_3338),
.A2(n_200),
.A3(n_198),
.B(n_199),
.Y(n_3425)
);

OAI21xp5_ASAP7_75t_L g3426 ( 
.A1(n_3256),
.A2(n_199),
.B(n_200),
.Y(n_3426)
);

OAI22xp5_ASAP7_75t_L g3427 ( 
.A1(n_3307),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3249),
.Y(n_3428)
);

OAI21x1_ASAP7_75t_L g3429 ( 
.A1(n_3347),
.A2(n_203),
.B(n_204),
.Y(n_3429)
);

OAI21x1_ASAP7_75t_L g3430 ( 
.A1(n_3363),
.A2(n_3219),
.B(n_3317),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3351),
.Y(n_3431)
);

OAI21x1_ASAP7_75t_L g3432 ( 
.A1(n_3361),
.A2(n_3230),
.B(n_3294),
.Y(n_3432)
);

OA21x2_ASAP7_75t_L g3433 ( 
.A1(n_3409),
.A2(n_3298),
.B(n_3284),
.Y(n_3433)
);

AO31x2_ASAP7_75t_L g3434 ( 
.A1(n_3350),
.A2(n_3283),
.A3(n_3265),
.B(n_3346),
.Y(n_3434)
);

INVx2_ASAP7_75t_L g3435 ( 
.A(n_3405),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3368),
.Y(n_3436)
);

OAI21xp5_ASAP7_75t_L g3437 ( 
.A1(n_3360),
.A2(n_3277),
.B(n_3315),
.Y(n_3437)
);

AOI21xp5_ASAP7_75t_L g3438 ( 
.A1(n_3353),
.A2(n_3358),
.B(n_3384),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_3379),
.B(n_3336),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3355),
.B(n_3385),
.Y(n_3440)
);

INVx3_ASAP7_75t_L g3441 ( 
.A(n_3422),
.Y(n_3441)
);

OA21x2_ASAP7_75t_L g3442 ( 
.A1(n_3365),
.A2(n_3310),
.B(n_3282),
.Y(n_3442)
);

AOI21xp5_ASAP7_75t_L g3443 ( 
.A1(n_3386),
.A2(n_3302),
.B(n_3247),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3371),
.B(n_3326),
.Y(n_3444)
);

AO21x2_ASAP7_75t_L g3445 ( 
.A1(n_3428),
.A2(n_3229),
.B(n_3269),
.Y(n_3445)
);

CKINVDCx8_ASAP7_75t_R g3446 ( 
.A(n_3377),
.Y(n_3446)
);

AOI21xp5_ASAP7_75t_SL g3447 ( 
.A1(n_3369),
.A2(n_3293),
.B(n_3333),
.Y(n_3447)
);

OAI21x1_ASAP7_75t_L g3448 ( 
.A1(n_3373),
.A2(n_3267),
.B(n_3225),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_3398),
.Y(n_3449)
);

OA21x2_ASAP7_75t_L g3450 ( 
.A1(n_3366),
.A2(n_3316),
.B(n_3291),
.Y(n_3450)
);

AND2x2_ASAP7_75t_L g3451 ( 
.A(n_3357),
.B(n_3226),
.Y(n_3451)
);

AOI22xp33_ASAP7_75t_L g3452 ( 
.A1(n_3408),
.A2(n_3331),
.B1(n_3286),
.B2(n_3234),
.Y(n_3452)
);

OAI21x1_ASAP7_75t_L g3453 ( 
.A1(n_3374),
.A2(n_3267),
.B(n_3348),
.Y(n_3453)
);

AOI21xp5_ASAP7_75t_L g3454 ( 
.A1(n_3349),
.A2(n_3303),
.B(n_3239),
.Y(n_3454)
);

BUFx10_ASAP7_75t_L g3455 ( 
.A(n_3376),
.Y(n_3455)
);

OA21x2_ASAP7_75t_L g3456 ( 
.A1(n_3394),
.A2(n_3260),
.B(n_3251),
.Y(n_3456)
);

OAI21x1_ASAP7_75t_L g3457 ( 
.A1(n_3392),
.A2(n_3308),
.B(n_3303),
.Y(n_3457)
);

AOI21xp33_ASAP7_75t_L g3458 ( 
.A1(n_3400),
.A2(n_3270),
.B(n_3259),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3378),
.Y(n_3459)
);

OR2x6_ASAP7_75t_L g3460 ( 
.A(n_3403),
.B(n_3324),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_3410),
.Y(n_3461)
);

OA21x2_ASAP7_75t_L g3462 ( 
.A1(n_3395),
.A2(n_3334),
.B(n_3240),
.Y(n_3462)
);

AOI32xp33_ASAP7_75t_L g3463 ( 
.A1(n_3389),
.A2(n_3240),
.A3(n_3275),
.B1(n_206),
.B2(n_204),
.Y(n_3463)
);

INVx2_ASAP7_75t_L g3464 ( 
.A(n_3402),
.Y(n_3464)
);

OAI21x1_ASAP7_75t_L g3465 ( 
.A1(n_3380),
.A2(n_3334),
.B(n_3274),
.Y(n_3465)
);

AO21x2_ASAP7_75t_L g3466 ( 
.A1(n_3370),
.A2(n_3330),
.B(n_205),
.Y(n_3466)
);

AOI21xp5_ASAP7_75t_L g3467 ( 
.A1(n_3362),
.A2(n_3330),
.B(n_205),
.Y(n_3467)
);

AND2x2_ASAP7_75t_L g3468 ( 
.A(n_3364),
.B(n_498),
.Y(n_3468)
);

CKINVDCx11_ASAP7_75t_R g3469 ( 
.A(n_3404),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3423),
.B(n_499),
.Y(n_3470)
);

OAI221xp5_ASAP7_75t_L g3471 ( 
.A1(n_3426),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.C(n_209),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3375),
.Y(n_3472)
);

AO21x2_ASAP7_75t_L g3473 ( 
.A1(n_3382),
.A2(n_207),
.B(n_208),
.Y(n_3473)
);

AND2x4_ASAP7_75t_L g3474 ( 
.A(n_3352),
.B(n_500),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3429),
.Y(n_3475)
);

OAI21x1_ASAP7_75t_L g3476 ( 
.A1(n_3396),
.A2(n_3399),
.B(n_3393),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_3413),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3375),
.Y(n_3478)
);

OAI21x1_ASAP7_75t_L g3479 ( 
.A1(n_3418),
.A2(n_209),
.B(n_210),
.Y(n_3479)
);

OAI21x1_ASAP7_75t_L g3480 ( 
.A1(n_3397),
.A2(n_210),
.B(n_211),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3421),
.Y(n_3481)
);

OA21x2_ASAP7_75t_L g3482 ( 
.A1(n_3390),
.A2(n_212),
.B(n_214),
.Y(n_3482)
);

HB1xp67_ASAP7_75t_L g3483 ( 
.A(n_3417),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3406),
.B(n_3356),
.Y(n_3484)
);

INVx4_ASAP7_75t_L g3485 ( 
.A(n_3416),
.Y(n_3485)
);

OAI22xp5_ASAP7_75t_L g3486 ( 
.A1(n_3383),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.Y(n_3486)
);

OAI21x1_ASAP7_75t_L g3487 ( 
.A1(n_3388),
.A2(n_217),
.B(n_218),
.Y(n_3487)
);

AO31x2_ASAP7_75t_L g3488 ( 
.A1(n_3387),
.A2(n_221),
.A3(n_219),
.B(n_220),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_3381),
.B(n_504),
.Y(n_3489)
);

AND2x2_ASAP7_75t_L g3490 ( 
.A(n_3391),
.B(n_506),
.Y(n_3490)
);

AO21x2_ASAP7_75t_L g3491 ( 
.A1(n_3420),
.A2(n_219),
.B(n_220),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3419),
.Y(n_3492)
);

AOI211xp5_ASAP7_75t_L g3493 ( 
.A1(n_3412),
.A2(n_224),
.B(n_222),
.C(n_223),
.Y(n_3493)
);

BUFx2_ASAP7_75t_L g3494 ( 
.A(n_3359),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3411),
.B(n_508),
.Y(n_3495)
);

AOI21xp5_ASAP7_75t_L g3496 ( 
.A1(n_3401),
.A2(n_222),
.B(n_223),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3354),
.B(n_3407),
.Y(n_3497)
);

INVx2_ASAP7_75t_L g3498 ( 
.A(n_3425),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3427),
.B(n_509),
.Y(n_3499)
);

BUFx6f_ASAP7_75t_L g3500 ( 
.A(n_3367),
.Y(n_3500)
);

AND2x4_ASAP7_75t_L g3501 ( 
.A(n_3372),
.B(n_510),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3431),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3436),
.Y(n_3503)
);

BUFx2_ASAP7_75t_L g3504 ( 
.A(n_3494),
.Y(n_3504)
);

AO21x2_ASAP7_75t_L g3505 ( 
.A1(n_3492),
.A2(n_3415),
.B(n_3424),
.Y(n_3505)
);

OR2x6_ASAP7_75t_L g3506 ( 
.A(n_3454),
.B(n_3414),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3449),
.Y(n_3507)
);

AND2x2_ASAP7_75t_L g3508 ( 
.A(n_3451),
.B(n_512),
.Y(n_3508)
);

INVx2_ASAP7_75t_L g3509 ( 
.A(n_3435),
.Y(n_3509)
);

OA21x2_ASAP7_75t_L g3510 ( 
.A1(n_3430),
.A2(n_515),
.B(n_514),
.Y(n_3510)
);

AO31x2_ASAP7_75t_L g3511 ( 
.A1(n_3498),
.A2(n_227),
.A3(n_225),
.B(n_226),
.Y(n_3511)
);

AO21x1_ASAP7_75t_SL g3512 ( 
.A1(n_3472),
.A2(n_226),
.B(n_227),
.Y(n_3512)
);

OR2x6_ASAP7_75t_L g3513 ( 
.A(n_3447),
.B(n_517),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3459),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3483),
.Y(n_3515)
);

OA21x2_ASAP7_75t_L g3516 ( 
.A1(n_3432),
.A2(n_3481),
.B(n_3465),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3461),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3475),
.Y(n_3518)
);

INVx2_ASAP7_75t_L g3519 ( 
.A(n_3464),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_3477),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_3448),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3478),
.Y(n_3522)
);

AO21x2_ASAP7_75t_L g3523 ( 
.A1(n_3438),
.A2(n_226),
.B(n_227),
.Y(n_3523)
);

BUFx6f_ASAP7_75t_L g3524 ( 
.A(n_3469),
.Y(n_3524)
);

HB1xp67_ASAP7_75t_L g3525 ( 
.A(n_3457),
.Y(n_3525)
);

INVx3_ASAP7_75t_L g3526 ( 
.A(n_3485),
.Y(n_3526)
);

INVx2_ASAP7_75t_SL g3527 ( 
.A(n_3455),
.Y(n_3527)
);

INVxp67_ASAP7_75t_L g3528 ( 
.A(n_3484),
.Y(n_3528)
);

HB1xp67_ASAP7_75t_L g3529 ( 
.A(n_3450),
.Y(n_3529)
);

BUFx3_ASAP7_75t_L g3530 ( 
.A(n_3446),
.Y(n_3530)
);

OAI21x1_ASAP7_75t_L g3531 ( 
.A1(n_3476),
.A2(n_228),
.B(n_229),
.Y(n_3531)
);

BUFx3_ASAP7_75t_L g3532 ( 
.A(n_3441),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_3444),
.B(n_518),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3456),
.Y(n_3534)
);

INVx4_ASAP7_75t_L g3535 ( 
.A(n_3500),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_3453),
.Y(n_3536)
);

INVx2_ASAP7_75t_L g3537 ( 
.A(n_3433),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3462),
.Y(n_3538)
);

BUFx4f_ASAP7_75t_L g3539 ( 
.A(n_3460),
.Y(n_3539)
);

AND2x2_ASAP7_75t_L g3540 ( 
.A(n_3468),
.B(n_519),
.Y(n_3540)
);

AND2x4_ASAP7_75t_SL g3541 ( 
.A(n_3474),
.B(n_519),
.Y(n_3541)
);

AND2x2_ASAP7_75t_L g3542 ( 
.A(n_3490),
.B(n_520),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3489),
.Y(n_3543)
);

OAI21xp5_ASAP7_75t_L g3544 ( 
.A1(n_3496),
.A2(n_228),
.B(n_229),
.Y(n_3544)
);

AOI22xp33_ASAP7_75t_SL g3545 ( 
.A1(n_3471),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3479),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3473),
.Y(n_3547)
);

BUFx2_ASAP7_75t_L g3548 ( 
.A(n_3442),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3466),
.Y(n_3549)
);

HB1xp67_ASAP7_75t_L g3550 ( 
.A(n_3434),
.Y(n_3550)
);

OAI21x1_ASAP7_75t_L g3551 ( 
.A1(n_3443),
.A2(n_230),
.B(n_232),
.Y(n_3551)
);

INVx2_ASAP7_75t_L g3552 ( 
.A(n_3434),
.Y(n_3552)
);

BUFx2_ASAP7_75t_SL g3553 ( 
.A(n_3501),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3480),
.Y(n_3554)
);

OA21x2_ASAP7_75t_L g3555 ( 
.A1(n_3437),
.A2(n_522),
.B(n_521),
.Y(n_3555)
);

INVxp67_ASAP7_75t_SL g3556 ( 
.A(n_3439),
.Y(n_3556)
);

INVx2_ASAP7_75t_L g3557 ( 
.A(n_3445),
.Y(n_3557)
);

INVx2_ASAP7_75t_L g3558 ( 
.A(n_3497),
.Y(n_3558)
);

OAI21x1_ASAP7_75t_L g3559 ( 
.A1(n_3467),
.A2(n_232),
.B(n_233),
.Y(n_3559)
);

AND2x2_ASAP7_75t_L g3560 ( 
.A(n_3470),
.B(n_522),
.Y(n_3560)
);

BUFx3_ASAP7_75t_L g3561 ( 
.A(n_3495),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_3491),
.Y(n_3562)
);

INVx1_ASAP7_75t_SL g3563 ( 
.A(n_3499),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3482),
.Y(n_3564)
);

OA21x2_ASAP7_75t_L g3565 ( 
.A1(n_3458),
.A2(n_524),
.B(n_523),
.Y(n_3565)
);

INVx3_ASAP7_75t_L g3566 ( 
.A(n_3488),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3488),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3487),
.Y(n_3568)
);

BUFx3_ASAP7_75t_L g3569 ( 
.A(n_3486),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3493),
.Y(n_3570)
);

AND2x4_ASAP7_75t_L g3571 ( 
.A(n_3452),
.B(n_525),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3463),
.Y(n_3572)
);

AND2x2_ASAP7_75t_L g3573 ( 
.A(n_3440),
.B(n_526),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3431),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_3449),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_SL g3576 ( 
.A(n_3438),
.B(n_526),
.Y(n_3576)
);

AND2x2_ASAP7_75t_L g3577 ( 
.A(n_3440),
.B(n_528),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3431),
.Y(n_3578)
);

INVxp67_ASAP7_75t_L g3579 ( 
.A(n_3440),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3556),
.B(n_529),
.Y(n_3580)
);

AND2x2_ASAP7_75t_L g3581 ( 
.A(n_3504),
.B(n_235),
.Y(n_3581)
);

AND2x2_ASAP7_75t_L g3582 ( 
.A(n_3579),
.B(n_236),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_3502),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3503),
.Y(n_3584)
);

OR2x6_ASAP7_75t_L g3585 ( 
.A(n_3524),
.B(n_532),
.Y(n_3585)
);

AOI221xp5_ASAP7_75t_L g3586 ( 
.A1(n_3576),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.C(n_240),
.Y(n_3586)
);

CKINVDCx20_ASAP7_75t_R g3587 ( 
.A(n_3530),
.Y(n_3587)
);

OAI211xp5_ASAP7_75t_SL g3588 ( 
.A1(n_3543),
.A2(n_241),
.B(n_238),
.C(n_239),
.Y(n_3588)
);

OAI21x1_ASAP7_75t_SL g3589 ( 
.A1(n_3562),
.A2(n_241),
.B(n_242),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_3578),
.Y(n_3590)
);

AOI22xp33_ASAP7_75t_L g3591 ( 
.A1(n_3569),
.A2(n_535),
.B1(n_536),
.B2(n_534),
.Y(n_3591)
);

AOI222xp33_ASAP7_75t_L g3592 ( 
.A1(n_3544),
.A2(n_244),
.B1(n_246),
.B2(n_242),
.C1(n_243),
.C2(n_245),
.Y(n_3592)
);

A2O1A1Ixp33_ASAP7_75t_L g3593 ( 
.A1(n_3545),
.A2(n_536),
.B(n_537),
.C(n_535),
.Y(n_3593)
);

BUFx2_ASAP7_75t_L g3594 ( 
.A(n_3524),
.Y(n_3594)
);

OA21x2_ASAP7_75t_L g3595 ( 
.A1(n_3548),
.A2(n_243),
.B(n_244),
.Y(n_3595)
);

OAI22xp5_ASAP7_75t_L g3596 ( 
.A1(n_3539),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.Y(n_3596)
);

AND2x2_ASAP7_75t_L g3597 ( 
.A(n_3558),
.B(n_246),
.Y(n_3597)
);

INVx4_ASAP7_75t_L g3598 ( 
.A(n_3535),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3574),
.Y(n_3599)
);

AOI221xp5_ASAP7_75t_L g3600 ( 
.A1(n_3567),
.A2(n_3533),
.B1(n_3566),
.B2(n_3563),
.C(n_3549),
.Y(n_3600)
);

AOI22xp33_ASAP7_75t_L g3601 ( 
.A1(n_3506),
.A2(n_542),
.B1(n_543),
.B2(n_541),
.Y(n_3601)
);

AOI22xp33_ASAP7_75t_L g3602 ( 
.A1(n_3506),
.A2(n_547),
.B1(n_548),
.B2(n_544),
.Y(n_3602)
);

OAI21x1_ASAP7_75t_L g3603 ( 
.A1(n_3557),
.A2(n_248),
.B(n_249),
.Y(n_3603)
);

NOR2xp33_ASAP7_75t_L g3604 ( 
.A(n_3528),
.B(n_549),
.Y(n_3604)
);

OAI22xp33_ASAP7_75t_L g3605 ( 
.A1(n_3555),
.A2(n_551),
.B1(n_552),
.B2(n_550),
.Y(n_3605)
);

OAI21x1_ASAP7_75t_L g3606 ( 
.A1(n_3534),
.A2(n_251),
.B(n_252),
.Y(n_3606)
);

AOI22xp33_ASAP7_75t_L g3607 ( 
.A1(n_3561),
.A2(n_554),
.B1(n_555),
.B2(n_552),
.Y(n_3607)
);

AOI22xp33_ASAP7_75t_SL g3608 ( 
.A1(n_3571),
.A2(n_556),
.B1(n_557),
.B2(n_555),
.Y(n_3608)
);

INVx2_ASAP7_75t_L g3609 ( 
.A(n_3575),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_SL g3610 ( 
.A(n_3526),
.B(n_556),
.Y(n_3610)
);

OAI21xp5_ASAP7_75t_L g3611 ( 
.A1(n_3551),
.A2(n_560),
.B(n_558),
.Y(n_3611)
);

AOI221xp5_ASAP7_75t_L g3612 ( 
.A1(n_3564),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.C(n_256),
.Y(n_3612)
);

INVx2_ASAP7_75t_L g3613 ( 
.A(n_3517),
.Y(n_3613)
);

AND2x2_ASAP7_75t_L g3614 ( 
.A(n_3507),
.B(n_3514),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3522),
.Y(n_3615)
);

OA21x2_ASAP7_75t_L g3616 ( 
.A1(n_3538),
.A2(n_256),
.B(n_258),
.Y(n_3616)
);

AOI22xp33_ASAP7_75t_L g3617 ( 
.A1(n_3505),
.A2(n_561),
.B1(n_562),
.B2(n_560),
.Y(n_3617)
);

AOI21xp33_ASAP7_75t_L g3618 ( 
.A1(n_3554),
.A2(n_3568),
.B(n_3546),
.Y(n_3618)
);

AOI22xp33_ASAP7_75t_L g3619 ( 
.A1(n_3523),
.A2(n_565),
.B1(n_567),
.B2(n_563),
.Y(n_3619)
);

OAI21x1_ASAP7_75t_L g3620 ( 
.A1(n_3552),
.A2(n_259),
.B(n_261),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3515),
.Y(n_3621)
);

INVx2_ASAP7_75t_L g3622 ( 
.A(n_3509),
.Y(n_3622)
);

AOI221xp5_ASAP7_75t_L g3623 ( 
.A1(n_3547),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.C(n_265),
.Y(n_3623)
);

AOI22xp33_ASAP7_75t_L g3624 ( 
.A1(n_3553),
.A2(n_570),
.B1(n_571),
.B2(n_569),
.Y(n_3624)
);

OAI21x1_ASAP7_75t_L g3625 ( 
.A1(n_3521),
.A2(n_262),
.B(n_263),
.Y(n_3625)
);

AOI22xp33_ASAP7_75t_SL g3626 ( 
.A1(n_3510),
.A2(n_572),
.B1(n_573),
.B2(n_570),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3529),
.Y(n_3627)
);

AOI33xp33_ASAP7_75t_L g3628 ( 
.A1(n_3560),
.A2(n_267),
.A3(n_269),
.B1(n_265),
.B2(n_266),
.B3(n_268),
.Y(n_3628)
);

BUFx6f_ASAP7_75t_SL g3629 ( 
.A(n_3527),
.Y(n_3629)
);

AND2x2_ASAP7_75t_L g3630 ( 
.A(n_3532),
.B(n_266),
.Y(n_3630)
);

NAND2x1p5_ASAP7_75t_L g3631 ( 
.A(n_3516),
.B(n_578),
.Y(n_3631)
);

AOI22xp33_ASAP7_75t_L g3632 ( 
.A1(n_3565),
.A2(n_580),
.B1(n_581),
.B2(n_579),
.Y(n_3632)
);

AOI21xp5_ASAP7_75t_L g3633 ( 
.A1(n_3537),
.A2(n_267),
.B(n_268),
.Y(n_3633)
);

AOI22x1_ASAP7_75t_L g3634 ( 
.A1(n_3550),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_3634)
);

HB1xp67_ASAP7_75t_L g3635 ( 
.A(n_3520),
.Y(n_3635)
);

HB1xp67_ASAP7_75t_L g3636 ( 
.A(n_3518),
.Y(n_3636)
);

INVx2_ASAP7_75t_L g3637 ( 
.A(n_3519),
.Y(n_3637)
);

OAI21x1_ASAP7_75t_L g3638 ( 
.A1(n_3536),
.A2(n_270),
.B(n_272),
.Y(n_3638)
);

AOI22xp33_ASAP7_75t_L g3639 ( 
.A1(n_3573),
.A2(n_587),
.B1(n_589),
.B2(n_586),
.Y(n_3639)
);

AOI22xp33_ASAP7_75t_L g3640 ( 
.A1(n_3577),
.A2(n_590),
.B1(n_591),
.B2(n_589),
.Y(n_3640)
);

OAI22xp5_ASAP7_75t_L g3641 ( 
.A1(n_3541),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_3641)
);

INVx4_ASAP7_75t_SL g3642 ( 
.A(n_3511),
.Y(n_3642)
);

OA21x2_ASAP7_75t_L g3643 ( 
.A1(n_3531),
.A2(n_276),
.B(n_278),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3525),
.Y(n_3644)
);

AOI22xp33_ASAP7_75t_L g3645 ( 
.A1(n_3559),
.A2(n_593),
.B1(n_595),
.B2(n_592),
.Y(n_3645)
);

AND2x2_ASAP7_75t_L g3646 ( 
.A(n_3508),
.B(n_278),
.Y(n_3646)
);

AOI221xp5_ASAP7_75t_L g3647 ( 
.A1(n_3542),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.C(n_283),
.Y(n_3647)
);

AOI22xp5_ASAP7_75t_L g3648 ( 
.A1(n_3540),
.A2(n_597),
.B1(n_598),
.B2(n_596),
.Y(n_3648)
);

OAI22xp33_ASAP7_75t_L g3649 ( 
.A1(n_3512),
.A2(n_598),
.B1(n_599),
.B2(n_597),
.Y(n_3649)
);

AOI221xp5_ASAP7_75t_L g3650 ( 
.A1(n_3570),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.C(n_284),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3502),
.Y(n_3651)
);

AOI211xp5_ASAP7_75t_L g3652 ( 
.A1(n_3570),
.A2(n_286),
.B(n_284),
.C(n_285),
.Y(n_3652)
);

INVx3_ASAP7_75t_SL g3653 ( 
.A(n_3524),
.Y(n_3653)
);

OAI22xp33_ASAP7_75t_L g3654 ( 
.A1(n_3513),
.A2(n_601),
.B1(n_603),
.B2(n_600),
.Y(n_3654)
);

BUFx2_ASAP7_75t_L g3655 ( 
.A(n_3504),
.Y(n_3655)
);

BUFx6f_ASAP7_75t_L g3656 ( 
.A(n_3524),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3504),
.B(n_287),
.Y(n_3657)
);

AOI22xp33_ASAP7_75t_L g3658 ( 
.A1(n_3572),
.A2(n_605),
.B1(n_606),
.B2(n_603),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3502),
.Y(n_3659)
);

BUFx12f_ASAP7_75t_L g3660 ( 
.A(n_3524),
.Y(n_3660)
);

AOI22xp33_ASAP7_75t_L g3661 ( 
.A1(n_3572),
.A2(n_606),
.B1(n_607),
.B2(n_605),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3615),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3600),
.B(n_607),
.Y(n_3663)
);

INVx2_ASAP7_75t_L g3664 ( 
.A(n_3644),
.Y(n_3664)
);

OR2x2_ASAP7_75t_L g3665 ( 
.A(n_3613),
.B(n_288),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3637),
.Y(n_3666)
);

AND2x2_ASAP7_75t_L g3667 ( 
.A(n_3635),
.B(n_288),
.Y(n_3667)
);

INVx1_ASAP7_75t_L g3668 ( 
.A(n_3621),
.Y(n_3668)
);

AND2x2_ASAP7_75t_L g3669 ( 
.A(n_3636),
.B(n_289),
.Y(n_3669)
);

INVx1_ASAP7_75t_SL g3670 ( 
.A(n_3653),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3583),
.Y(n_3671)
);

OR2x2_ASAP7_75t_L g3672 ( 
.A(n_3622),
.B(n_289),
.Y(n_3672)
);

INVx2_ASAP7_75t_L g3673 ( 
.A(n_3590),
.Y(n_3673)
);

INVx4_ASAP7_75t_L g3674 ( 
.A(n_3656),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_3614),
.B(n_608),
.Y(n_3675)
);

INVxp67_ASAP7_75t_SL g3676 ( 
.A(n_3631),
.Y(n_3676)
);

BUFx2_ASAP7_75t_L g3677 ( 
.A(n_3594),
.Y(n_3677)
);

AOI22xp33_ASAP7_75t_SL g3678 ( 
.A1(n_3634),
.A2(n_610),
.B1(n_611),
.B2(n_609),
.Y(n_3678)
);

AND2x2_ASAP7_75t_L g3679 ( 
.A(n_3609),
.B(n_290),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_L g3680 ( 
.A(n_3584),
.B(n_610),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3599),
.B(n_612),
.Y(n_3681)
);

NOR2xp33_ASAP7_75t_R g3682 ( 
.A(n_3587),
.B(n_291),
.Y(n_3682)
);

OR2x2_ASAP7_75t_L g3683 ( 
.A(n_3651),
.B(n_292),
.Y(n_3683)
);

INVx3_ASAP7_75t_L g3684 ( 
.A(n_3598),
.Y(n_3684)
);

HB1xp67_ASAP7_75t_L g3685 ( 
.A(n_3642),
.Y(n_3685)
);

INVx2_ASAP7_75t_L g3686 ( 
.A(n_3659),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3642),
.Y(n_3687)
);

INVxp67_ASAP7_75t_SL g3688 ( 
.A(n_3580),
.Y(n_3688)
);

BUFx3_ASAP7_75t_L g3689 ( 
.A(n_3630),
.Y(n_3689)
);

AND2x2_ASAP7_75t_L g3690 ( 
.A(n_3581),
.B(n_293),
.Y(n_3690)
);

BUFx12f_ASAP7_75t_L g3691 ( 
.A(n_3585),
.Y(n_3691)
);

AND2x2_ASAP7_75t_L g3692 ( 
.A(n_3657),
.B(n_296),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_SL g3693 ( 
.A(n_3605),
.B(n_613),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3595),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_SL g3695 ( 
.A(n_3604),
.B(n_614),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3616),
.Y(n_3696)
);

AND2x4_ASAP7_75t_SL g3697 ( 
.A(n_3585),
.B(n_615),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_SL g3698 ( 
.A(n_3652),
.B(n_3582),
.Y(n_3698)
);

NOR2xp33_ASAP7_75t_L g3699 ( 
.A(n_3629),
.B(n_615),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3597),
.B(n_616),
.Y(n_3700)
);

AND2x2_ASAP7_75t_L g3701 ( 
.A(n_3618),
.B(n_297),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3620),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3643),
.Y(n_3703)
);

AND2x2_ASAP7_75t_L g3704 ( 
.A(n_3646),
.B(n_298),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3603),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3638),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3606),
.Y(n_3707)
);

AOI22xp5_ASAP7_75t_L g3708 ( 
.A1(n_3592),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_3589),
.Y(n_3709)
);

NOR2xp33_ASAP7_75t_L g3710 ( 
.A(n_3610),
.B(n_1395),
.Y(n_3710)
);

INVx2_ASAP7_75t_L g3711 ( 
.A(n_3625),
.Y(n_3711)
);

AOI21xp5_ASAP7_75t_SL g3712 ( 
.A1(n_3586),
.A2(n_300),
.B(n_301),
.Y(n_3712)
);

BUFx2_ASAP7_75t_L g3713 ( 
.A(n_3611),
.Y(n_3713)
);

AND2x2_ASAP7_75t_L g3714 ( 
.A(n_3626),
.B(n_302),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3633),
.B(n_617),
.Y(n_3715)
);

AND2x2_ASAP7_75t_L g3716 ( 
.A(n_3648),
.B(n_303),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3628),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3632),
.B(n_618),
.Y(n_3718)
);

INVxp67_ASAP7_75t_SL g3719 ( 
.A(n_3649),
.Y(n_3719)
);

NOR2xp33_ASAP7_75t_L g3720 ( 
.A(n_3596),
.B(n_1399),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3601),
.B(n_619),
.Y(n_3721)
);

INVx2_ASAP7_75t_L g3722 ( 
.A(n_3641),
.Y(n_3722)
);

AND2x2_ASAP7_75t_L g3723 ( 
.A(n_3645),
.B(n_304),
.Y(n_3723)
);

AOI221xp5_ASAP7_75t_L g3724 ( 
.A1(n_3650),
.A2(n_307),
.B1(n_305),
.B2(n_306),
.C(n_308),
.Y(n_3724)
);

OR2x2_ASAP7_75t_L g3725 ( 
.A(n_3619),
.B(n_305),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3588),
.Y(n_3726)
);

INVx3_ASAP7_75t_L g3727 ( 
.A(n_3654),
.Y(n_3727)
);

AND2x4_ASAP7_75t_SL g3728 ( 
.A(n_3624),
.B(n_619),
.Y(n_3728)
);

AND2x6_ASAP7_75t_L g3729 ( 
.A(n_3608),
.B(n_306),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3602),
.B(n_620),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3612),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3639),
.B(n_306),
.Y(n_3732)
);

HB1xp67_ASAP7_75t_L g3733 ( 
.A(n_3623),
.Y(n_3733)
);

AND2x2_ASAP7_75t_L g3734 ( 
.A(n_3640),
.B(n_307),
.Y(n_3734)
);

HB1xp67_ASAP7_75t_L g3735 ( 
.A(n_3647),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3593),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3607),
.B(n_621),
.Y(n_3737)
);

NAND2x1p5_ASAP7_75t_SL g3738 ( 
.A(n_3591),
.B(n_310),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3658),
.Y(n_3739)
);

AND2x2_ASAP7_75t_L g3740 ( 
.A(n_3661),
.B(n_310),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3615),
.Y(n_3741)
);

BUFx3_ASAP7_75t_L g3742 ( 
.A(n_3660),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3600),
.B(n_622),
.Y(n_3743)
);

INVx2_ASAP7_75t_L g3744 ( 
.A(n_3644),
.Y(n_3744)
);

AND2x4_ASAP7_75t_L g3745 ( 
.A(n_3655),
.B(n_622),
.Y(n_3745)
);

AND2x2_ASAP7_75t_L g3746 ( 
.A(n_3655),
.B(n_311),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3615),
.Y(n_3747)
);

AND2x2_ASAP7_75t_L g3748 ( 
.A(n_3655),
.B(n_312),
.Y(n_3748)
);

OAI22xp5_ASAP7_75t_L g3749 ( 
.A1(n_3617),
.A2(n_314),
.B1(n_312),
.B2(n_313),
.Y(n_3749)
);

AND2x2_ASAP7_75t_L g3750 ( 
.A(n_3655),
.B(n_312),
.Y(n_3750)
);

HB1xp67_ASAP7_75t_L g3751 ( 
.A(n_3627),
.Y(n_3751)
);

INVx2_ASAP7_75t_L g3752 ( 
.A(n_3644),
.Y(n_3752)
);

BUFx2_ASAP7_75t_L g3753 ( 
.A(n_3655),
.Y(n_3753)
);

AND2x2_ASAP7_75t_L g3754 ( 
.A(n_3753),
.B(n_315),
.Y(n_3754)
);

NOR2x1p5_ASAP7_75t_L g3755 ( 
.A(n_3691),
.B(n_316),
.Y(n_3755)
);

INVxp67_ASAP7_75t_L g3756 ( 
.A(n_3694),
.Y(n_3756)
);

INVx2_ASAP7_75t_L g3757 ( 
.A(n_3677),
.Y(n_3757)
);

OA21x2_ASAP7_75t_L g3758 ( 
.A1(n_3687),
.A2(n_316),
.B(n_317),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_3705),
.B(n_623),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_3666),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3671),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3676),
.B(n_319),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_3706),
.B(n_624),
.Y(n_3763)
);

INVx2_ASAP7_75t_L g3764 ( 
.A(n_3673),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_3707),
.B(n_625),
.Y(n_3765)
);

NAND2x1_ASAP7_75t_L g3766 ( 
.A(n_3696),
.B(n_3664),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3711),
.B(n_626),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3741),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_3702),
.B(n_3701),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3747),
.Y(n_3770)
);

AND2x4_ASAP7_75t_L g3771 ( 
.A(n_3689),
.B(n_320),
.Y(n_3771)
);

AND2x4_ASAP7_75t_SL g3772 ( 
.A(n_3674),
.B(n_321),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3686),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3703),
.B(n_3719),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3668),
.Y(n_3775)
);

AND2x4_ASAP7_75t_SL g3776 ( 
.A(n_3745),
.B(n_321),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3667),
.B(n_628),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3751),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_3669),
.B(n_3709),
.Y(n_3779)
);

INVxp67_ASAP7_75t_SL g3780 ( 
.A(n_3685),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3665),
.Y(n_3781)
);

INVx1_ASAP7_75t_L g3782 ( 
.A(n_3672),
.Y(n_3782)
);

HB1xp67_ASAP7_75t_L g3783 ( 
.A(n_3744),
.Y(n_3783)
);

INVxp33_ASAP7_75t_L g3784 ( 
.A(n_3682),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3752),
.B(n_322),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3680),
.B(n_630),
.Y(n_3786)
);

AND2x2_ASAP7_75t_L g3787 ( 
.A(n_3670),
.B(n_323),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_3681),
.B(n_632),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3727),
.B(n_633),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3679),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3683),
.Y(n_3791)
);

HB1xp67_ASAP7_75t_L g3792 ( 
.A(n_3746),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3675),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3722),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_3663),
.B(n_633),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3748),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3743),
.B(n_634),
.Y(n_3797)
);

NAND3xp33_ASAP7_75t_L g3798 ( 
.A(n_3733),
.B(n_324),
.C(n_325),
.Y(n_3798)
);

CKINVDCx5p33_ASAP7_75t_R g3799 ( 
.A(n_3697),
.Y(n_3799)
);

HB1xp67_ASAP7_75t_L g3800 ( 
.A(n_3750),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3690),
.B(n_325),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_L g3802 ( 
.A(n_3735),
.B(n_637),
.Y(n_3802)
);

INVx3_ASAP7_75t_L g3803 ( 
.A(n_3692),
.Y(n_3803)
);

AND2x2_ASAP7_75t_L g3804 ( 
.A(n_3704),
.B(n_326),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3700),
.Y(n_3805)
);

OR2x2_ASAP7_75t_L g3806 ( 
.A(n_3739),
.B(n_327),
.Y(n_3806)
);

NAND2x1_ASAP7_75t_SL g3807 ( 
.A(n_3699),
.B(n_328),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3726),
.Y(n_3808)
);

AND2x2_ASAP7_75t_L g3809 ( 
.A(n_3698),
.B(n_329),
.Y(n_3809)
);

AND2x2_ASAP7_75t_L g3810 ( 
.A(n_3736),
.B(n_329),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3715),
.Y(n_3811)
);

OR2x6_ASAP7_75t_SL g3812 ( 
.A(n_3731),
.B(n_638),
.Y(n_3812)
);

OAI221xp5_ASAP7_75t_SL g3813 ( 
.A1(n_3708),
.A2(n_642),
.B1(n_640),
.B2(n_641),
.C(n_644),
.Y(n_3813)
);

AND2x2_ASAP7_75t_L g3814 ( 
.A(n_3716),
.B(n_3717),
.Y(n_3814)
);

HB1xp67_ASAP7_75t_L g3815 ( 
.A(n_3695),
.Y(n_3815)
);

INVx2_ASAP7_75t_L g3816 ( 
.A(n_3693),
.Y(n_3816)
);

INVx2_ASAP7_75t_L g3817 ( 
.A(n_3714),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_3710),
.B(n_644),
.Y(n_3818)
);

AND2x2_ASAP7_75t_L g3819 ( 
.A(n_3720),
.B(n_645),
.Y(n_3819)
);

AND2x2_ASAP7_75t_L g3820 ( 
.A(n_3732),
.B(n_645),
.Y(n_3820)
);

AND2x2_ASAP7_75t_L g3821 ( 
.A(n_3734),
.B(n_646),
.Y(n_3821)
);

OR2x2_ASAP7_75t_L g3822 ( 
.A(n_3718),
.B(n_648),
.Y(n_3822)
);

INVx2_ASAP7_75t_L g3823 ( 
.A(n_3725),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3729),
.B(n_649),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3723),
.Y(n_3825)
);

AND2x2_ASAP7_75t_L g3826 ( 
.A(n_3740),
.B(n_650),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_3721),
.B(n_651),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3730),
.Y(n_3828)
);

AND2x2_ASAP7_75t_L g3829 ( 
.A(n_3728),
.B(n_652),
.Y(n_3829)
);

AND2x2_ASAP7_75t_L g3830 ( 
.A(n_3737),
.B(n_655),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_SL g3831 ( 
.A(n_3678),
.B(n_656),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3724),
.B(n_656),
.Y(n_3832)
);

AND2x2_ASAP7_75t_L g3833 ( 
.A(n_3749),
.B(n_658),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_L g3834 ( 
.A(n_3738),
.B(n_658),
.Y(n_3834)
);

OR2x2_ASAP7_75t_L g3835 ( 
.A(n_3688),
.B(n_660),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3662),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3662),
.Y(n_3837)
);

AND2x2_ASAP7_75t_L g3838 ( 
.A(n_3753),
.B(n_661),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_SL g3839 ( 
.A(n_3684),
.B(n_663),
.Y(n_3839)
);

OR2x2_ASAP7_75t_L g3840 ( 
.A(n_3688),
.B(n_663),
.Y(n_3840)
);

AND2x2_ASAP7_75t_L g3841 ( 
.A(n_3753),
.B(n_664),
.Y(n_3841)
);

INVx3_ASAP7_75t_L g3842 ( 
.A(n_3674),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3662),
.Y(n_3843)
);

AND4x1_ASAP7_75t_L g3844 ( 
.A(n_3712),
.B(n_667),
.C(n_665),
.D(n_666),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3688),
.B(n_666),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3662),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3688),
.B(n_669),
.Y(n_3847)
);

INVxp67_ASAP7_75t_SL g3848 ( 
.A(n_3753),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_3688),
.B(n_670),
.Y(n_3849)
);

AND2x2_ASAP7_75t_L g3850 ( 
.A(n_3753),
.B(n_671),
.Y(n_3850)
);

INVx3_ASAP7_75t_L g3851 ( 
.A(n_3674),
.Y(n_3851)
);

OR2x2_ASAP7_75t_L g3852 ( 
.A(n_3688),
.B(n_671),
.Y(n_3852)
);

AND2x2_ASAP7_75t_L g3853 ( 
.A(n_3753),
.B(n_672),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_SL g3854 ( 
.A(n_3684),
.B(n_673),
.Y(n_3854)
);

AND2x2_ASAP7_75t_L g3855 ( 
.A(n_3753),
.B(n_673),
.Y(n_3855)
);

INVx2_ASAP7_75t_SL g3856 ( 
.A(n_3742),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3662),
.Y(n_3857)
);

AND2x2_ASAP7_75t_L g3858 ( 
.A(n_3753),
.B(n_675),
.Y(n_3858)
);

AND2x4_ASAP7_75t_L g3859 ( 
.A(n_3677),
.B(n_675),
.Y(n_3859)
);

OAI221xp5_ASAP7_75t_L g3860 ( 
.A1(n_3713),
.A2(n_679),
.B1(n_676),
.B2(n_678),
.C(n_680),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3753),
.B(n_681),
.Y(n_3861)
);

AND2x2_ASAP7_75t_L g3862 ( 
.A(n_3753),
.B(n_681),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3781),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3782),
.Y(n_3864)
);

INVx1_ASAP7_75t_SL g3865 ( 
.A(n_3807),
.Y(n_3865)
);

NAND3xp33_ASAP7_75t_L g3866 ( 
.A(n_3844),
.B(n_684),
.C(n_686),
.Y(n_3866)
);

AO21x2_ASAP7_75t_L g3867 ( 
.A1(n_3774),
.A2(n_686),
.B(n_687),
.Y(n_3867)
);

AOI22xp33_ASAP7_75t_L g3868 ( 
.A1(n_3816),
.A2(n_690),
.B1(n_688),
.B2(n_689),
.Y(n_3868)
);

AND2x4_ASAP7_75t_L g3869 ( 
.A(n_3842),
.B(n_691),
.Y(n_3869)
);

AND2x2_ASAP7_75t_L g3870 ( 
.A(n_3848),
.B(n_693),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_3851),
.Y(n_3871)
);

AOI22xp33_ASAP7_75t_SL g3872 ( 
.A1(n_3815),
.A2(n_696),
.B1(n_694),
.B2(n_695),
.Y(n_3872)
);

INVxp67_ASAP7_75t_SL g3873 ( 
.A(n_3792),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3768),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3770),
.Y(n_3875)
);

BUFx3_ASAP7_75t_L g3876 ( 
.A(n_3772),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3808),
.B(n_3794),
.Y(n_3877)
);

AND2x2_ASAP7_75t_L g3878 ( 
.A(n_3757),
.B(n_698),
.Y(n_3878)
);

OAI221xp5_ASAP7_75t_L g3879 ( 
.A1(n_3756),
.A2(n_702),
.B1(n_699),
.B2(n_701),
.C(n_703),
.Y(n_3879)
);

AND2x4_ASAP7_75t_L g3880 ( 
.A(n_3856),
.B(n_699),
.Y(n_3880)
);

NOR2x1_ASAP7_75t_L g3881 ( 
.A(n_3758),
.B(n_701),
.Y(n_3881)
);

NAND4xp25_ASAP7_75t_SL g3882 ( 
.A(n_3798),
.B(n_709),
.C(n_707),
.D(n_708),
.Y(n_3882)
);

AOI221xp5_ASAP7_75t_L g3883 ( 
.A1(n_3860),
.A2(n_710),
.B1(n_708),
.B2(n_709),
.C(n_711),
.Y(n_3883)
);

NAND4xp25_ASAP7_75t_L g3884 ( 
.A(n_3813),
.B(n_712),
.C(n_713),
.D(n_711),
.Y(n_3884)
);

OR2x2_ASAP7_75t_L g3885 ( 
.A(n_3769),
.B(n_710),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3775),
.Y(n_3886)
);

AOI31xp33_ASAP7_75t_L g3887 ( 
.A1(n_3784),
.A2(n_719),
.A3(n_717),
.B(n_718),
.Y(n_3887)
);

NAND2x1p5_ASAP7_75t_L g3888 ( 
.A(n_3766),
.B(n_722),
.Y(n_3888)
);

OR2x2_ASAP7_75t_SL g3889 ( 
.A(n_3800),
.B(n_723),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3836),
.Y(n_3890)
);

OAI22xp5_ASAP7_75t_L g3891 ( 
.A1(n_3812),
.A2(n_728),
.B1(n_725),
.B2(n_727),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3837),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_3843),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3846),
.Y(n_3894)
);

NOR3xp33_ASAP7_75t_L g3895 ( 
.A(n_3831),
.B(n_733),
.C(n_734),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3857),
.Y(n_3896)
);

NOR2x1_ASAP7_75t_R g3897 ( 
.A(n_3799),
.B(n_735),
.Y(n_3897)
);

OAI33xp33_ASAP7_75t_L g3898 ( 
.A1(n_3802),
.A2(n_739),
.A3(n_741),
.B1(n_737),
.B2(n_738),
.B3(n_740),
.Y(n_3898)
);

BUFx2_ASAP7_75t_L g3899 ( 
.A(n_3780),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3791),
.Y(n_3900)
);

BUFx2_ASAP7_75t_L g3901 ( 
.A(n_3803),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3773),
.Y(n_3902)
);

INVx4_ASAP7_75t_L g3903 ( 
.A(n_3771),
.Y(n_3903)
);

NAND3xp33_ASAP7_75t_SL g3904 ( 
.A(n_3834),
.B(n_745),
.C(n_746),
.Y(n_3904)
);

OAI21xp33_ASAP7_75t_L g3905 ( 
.A1(n_3832),
.A2(n_747),
.B(n_748),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3778),
.Y(n_3906)
);

NOR2xp33_ASAP7_75t_SL g3907 ( 
.A(n_3859),
.B(n_747),
.Y(n_3907)
);

INVx2_ASAP7_75t_L g3908 ( 
.A(n_3760),
.Y(n_3908)
);

A2O1A1Ixp33_ASAP7_75t_SL g3909 ( 
.A1(n_3759),
.A2(n_751),
.B(n_749),
.C(n_750),
.Y(n_3909)
);

NAND2xp5_ASAP7_75t_L g3910 ( 
.A(n_3811),
.B(n_3828),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3805),
.B(n_753),
.Y(n_3911)
);

AND2x4_ASAP7_75t_L g3912 ( 
.A(n_3790),
.B(n_755),
.Y(n_3912)
);

NOR3xp33_ASAP7_75t_L g3913 ( 
.A(n_3795),
.B(n_755),
.C(n_756),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3793),
.B(n_757),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3761),
.Y(n_3915)
);

AND2x4_ASAP7_75t_SL g3916 ( 
.A(n_3787),
.B(n_758),
.Y(n_3916)
);

HB1xp67_ASAP7_75t_L g3917 ( 
.A(n_3783),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3764),
.Y(n_3918)
);

AND2x4_ASAP7_75t_L g3919 ( 
.A(n_3796),
.B(n_759),
.Y(n_3919)
);

BUFx3_ASAP7_75t_L g3920 ( 
.A(n_3776),
.Y(n_3920)
);

OAI31xp33_ASAP7_75t_L g3921 ( 
.A1(n_3755),
.A2(n_3833),
.A3(n_3809),
.B(n_3824),
.Y(n_3921)
);

BUFx2_ASAP7_75t_SL g3922 ( 
.A(n_3754),
.Y(n_3922)
);

NAND3xp33_ASAP7_75t_L g3923 ( 
.A(n_3797),
.B(n_759),
.C(n_760),
.Y(n_3923)
);

NOR2x1_ASAP7_75t_L g3924 ( 
.A(n_3835),
.B(n_3840),
.Y(n_3924)
);

OR2x2_ASAP7_75t_L g3925 ( 
.A(n_3779),
.B(n_763),
.Y(n_3925)
);

AND2x2_ASAP7_75t_L g3926 ( 
.A(n_3823),
.B(n_3825),
.Y(n_3926)
);

INVxp67_ASAP7_75t_SL g3927 ( 
.A(n_3817),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3785),
.Y(n_3928)
);

INVxp67_ASAP7_75t_L g3929 ( 
.A(n_3814),
.Y(n_3929)
);

NOR2x1_ASAP7_75t_L g3930 ( 
.A(n_3852),
.B(n_764),
.Y(n_3930)
);

OAI22xp5_ASAP7_75t_SL g3931 ( 
.A1(n_3789),
.A2(n_767),
.B1(n_765),
.B2(n_766),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3838),
.B(n_768),
.Y(n_3932)
);

NOR2xp33_ASAP7_75t_L g3933 ( 
.A(n_3806),
.B(n_769),
.Y(n_3933)
);

OAI31xp33_ASAP7_75t_SL g3934 ( 
.A1(n_3839),
.A2(n_772),
.A3(n_773),
.B(n_771),
.Y(n_3934)
);

INVx2_ASAP7_75t_SL g3935 ( 
.A(n_3841),
.Y(n_3935)
);

AOI221x1_ASAP7_75t_L g3936 ( 
.A1(n_3767),
.A2(n_772),
.B1(n_770),
.B2(n_771),
.C(n_773),
.Y(n_3936)
);

OAI31xp33_ASAP7_75t_L g3937 ( 
.A1(n_3819),
.A2(n_776),
.A3(n_774),
.B(n_775),
.Y(n_3937)
);

NAND3xp33_ASAP7_75t_L g3938 ( 
.A(n_3763),
.B(n_777),
.C(n_778),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3873),
.Y(n_3939)
);

NAND3xp33_ASAP7_75t_L g3940 ( 
.A(n_3934),
.B(n_3765),
.C(n_3827),
.Y(n_3940)
);

OAI21xp33_ASAP7_75t_L g3941 ( 
.A1(n_3884),
.A2(n_3818),
.B(n_3822),
.Y(n_3941)
);

AND2x2_ASAP7_75t_L g3942 ( 
.A(n_3922),
.B(n_3762),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3899),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_L g3944 ( 
.A(n_3865),
.B(n_3935),
.Y(n_3944)
);

NOR2x1_ASAP7_75t_L g3945 ( 
.A(n_3867),
.B(n_3853),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3917),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_SL g3947 ( 
.A(n_3888),
.B(n_3845),
.Y(n_3947)
);

INVx4_ASAP7_75t_L g3948 ( 
.A(n_3869),
.Y(n_3948)
);

AND2x2_ASAP7_75t_L g3949 ( 
.A(n_3871),
.B(n_3850),
.Y(n_3949)
);

OR2x2_ASAP7_75t_L g3950 ( 
.A(n_3927),
.B(n_3847),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3926),
.Y(n_3951)
);

INVx1_ASAP7_75t_SL g3952 ( 
.A(n_3876),
.Y(n_3952)
);

AND2x2_ASAP7_75t_L g3953 ( 
.A(n_3901),
.B(n_3855),
.Y(n_3953)
);

AND2x2_ASAP7_75t_L g3954 ( 
.A(n_3903),
.B(n_3858),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3881),
.B(n_3810),
.Y(n_3955)
);

AND2x2_ASAP7_75t_L g3956 ( 
.A(n_3928),
.B(n_3861),
.Y(n_3956)
);

INVx4_ASAP7_75t_L g3957 ( 
.A(n_3880),
.Y(n_3957)
);

BUFx2_ASAP7_75t_L g3958 ( 
.A(n_3920),
.Y(n_3958)
);

INVx2_ASAP7_75t_L g3959 ( 
.A(n_3889),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_SL g3960 ( 
.A(n_3924),
.B(n_3849),
.Y(n_3960)
);

AND2x2_ASAP7_75t_L g3961 ( 
.A(n_3929),
.B(n_3862),
.Y(n_3961)
);

INVxp67_ASAP7_75t_L g3962 ( 
.A(n_3897),
.Y(n_3962)
);

INVxp33_ASAP7_75t_L g3963 ( 
.A(n_3921),
.Y(n_3963)
);

INVx2_ASAP7_75t_SL g3964 ( 
.A(n_3916),
.Y(n_3964)
);

OR2x6_ASAP7_75t_L g3965 ( 
.A(n_3930),
.B(n_3829),
.Y(n_3965)
);

BUFx2_ASAP7_75t_L g3966 ( 
.A(n_3870),
.Y(n_3966)
);

NOR2xp33_ASAP7_75t_L g3967 ( 
.A(n_3925),
.B(n_3786),
.Y(n_3967)
);

OR2x2_ASAP7_75t_L g3968 ( 
.A(n_3877),
.B(n_3788),
.Y(n_3968)
);

INVx1_ASAP7_75t_SL g3969 ( 
.A(n_3932),
.Y(n_3969)
);

OAI21xp5_ASAP7_75t_L g3970 ( 
.A1(n_3866),
.A2(n_3854),
.B(n_3830),
.Y(n_3970)
);

OR2x2_ASAP7_75t_L g3971 ( 
.A(n_3885),
.B(n_3777),
.Y(n_3971)
);

BUFx3_ASAP7_75t_L g3972 ( 
.A(n_3919),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3874),
.Y(n_3973)
);

NAND2x1p5_ASAP7_75t_L g3974 ( 
.A(n_3878),
.B(n_3801),
.Y(n_3974)
);

INVx2_ASAP7_75t_SL g3975 ( 
.A(n_3912),
.Y(n_3975)
);

INVx1_ASAP7_75t_L g3976 ( 
.A(n_3875),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3886),
.Y(n_3977)
);

AOI22xp5_ASAP7_75t_L g3978 ( 
.A1(n_3895),
.A2(n_3826),
.B1(n_3820),
.B2(n_3821),
.Y(n_3978)
);

HB1xp67_ASAP7_75t_L g3979 ( 
.A(n_3908),
.Y(n_3979)
);

AND2x2_ASAP7_75t_SL g3980 ( 
.A(n_3913),
.B(n_3804),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_3890),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3892),
.Y(n_3982)
);

OR2x2_ASAP7_75t_L g3983 ( 
.A(n_3910),
.B(n_1392),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_3933),
.B(n_779),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3893),
.Y(n_3985)
);

NAND3xp33_ASAP7_75t_L g3986 ( 
.A(n_3883),
.B(n_781),
.C(n_782),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3894),
.Y(n_3987)
);

AND2x4_ASAP7_75t_L g3988 ( 
.A(n_3863),
.B(n_1401),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3864),
.B(n_786),
.Y(n_3989)
);

INVxp67_ASAP7_75t_L g3990 ( 
.A(n_3907),
.Y(n_3990)
);

OR2x2_ASAP7_75t_L g3991 ( 
.A(n_3900),
.B(n_1389),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_L g3992 ( 
.A(n_3959),
.B(n_3891),
.Y(n_3992)
);

INVx2_ASAP7_75t_L g3993 ( 
.A(n_3958),
.Y(n_3993)
);

INVx2_ASAP7_75t_L g3994 ( 
.A(n_3964),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3942),
.B(n_3906),
.Y(n_3995)
);

HB1xp67_ASAP7_75t_L g3996 ( 
.A(n_3965),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_L g3997 ( 
.A(n_3966),
.B(n_3887),
.Y(n_3997)
);

INVx1_ASAP7_75t_SL g3998 ( 
.A(n_3952),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3939),
.Y(n_3999)
);

NOR2xp33_ASAP7_75t_L g4000 ( 
.A(n_3962),
.B(n_3911),
.Y(n_4000)
);

NOR2xp33_ASAP7_75t_SL g4001 ( 
.A(n_3948),
.B(n_3937),
.Y(n_4001)
);

AND2x2_ASAP7_75t_L g4002 ( 
.A(n_3954),
.B(n_3915),
.Y(n_4002)
);

AND2x2_ASAP7_75t_L g4003 ( 
.A(n_3953),
.B(n_3918),
.Y(n_4003)
);

NOR2xp33_ASAP7_75t_L g4004 ( 
.A(n_3957),
.B(n_3914),
.Y(n_4004)
);

HB1xp67_ASAP7_75t_L g4005 ( 
.A(n_3965),
.Y(n_4005)
);

INVx2_ASAP7_75t_SL g4006 ( 
.A(n_3972),
.Y(n_4006)
);

AND2x2_ASAP7_75t_L g4007 ( 
.A(n_3949),
.B(n_3902),
.Y(n_4007)
);

NAND2xp5_ASAP7_75t_L g4008 ( 
.A(n_3980),
.B(n_3905),
.Y(n_4008)
);

OR2x2_ASAP7_75t_L g4009 ( 
.A(n_3969),
.B(n_3904),
.Y(n_4009)
);

NAND2x1_ASAP7_75t_L g4010 ( 
.A(n_3945),
.B(n_3896),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_L g4011 ( 
.A(n_3990),
.B(n_3923),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_SL g4012 ( 
.A(n_3955),
.B(n_3872),
.Y(n_4012)
);

OR2x2_ASAP7_75t_L g4013 ( 
.A(n_3943),
.B(n_3938),
.Y(n_4013)
);

NOR2xp33_ASAP7_75t_L g4014 ( 
.A(n_3963),
.B(n_3931),
.Y(n_4014)
);

INVx2_ASAP7_75t_L g4015 ( 
.A(n_3974),
.Y(n_4015)
);

OR2x2_ASAP7_75t_L g4016 ( 
.A(n_3944),
.B(n_3882),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3946),
.Y(n_4017)
);

NOR2xp33_ASAP7_75t_L g4018 ( 
.A(n_3941),
.B(n_3898),
.Y(n_4018)
);

NOR2x1_ASAP7_75t_L g4019 ( 
.A(n_3986),
.B(n_3879),
.Y(n_4019)
);

BUFx2_ASAP7_75t_L g4020 ( 
.A(n_3975),
.Y(n_4020)
);

INVx2_ASAP7_75t_SL g4021 ( 
.A(n_3988),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3956),
.B(n_3936),
.Y(n_4022)
);

NAND2x1_ASAP7_75t_L g4023 ( 
.A(n_3961),
.B(n_3868),
.Y(n_4023)
);

OR2x2_ASAP7_75t_L g4024 ( 
.A(n_3950),
.B(n_3909),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3991),
.Y(n_4025)
);

OR2x2_ASAP7_75t_L g4026 ( 
.A(n_3951),
.B(n_3960),
.Y(n_4026)
);

NAND2x1p5_ASAP7_75t_L g4027 ( 
.A(n_3947),
.B(n_790),
.Y(n_4027)
);

BUFx2_ASAP7_75t_L g4028 ( 
.A(n_3979),
.Y(n_4028)
);

AND2x2_ASAP7_75t_L g4029 ( 
.A(n_3967),
.B(n_792),
.Y(n_4029)
);

AND2x2_ASAP7_75t_L g4030 ( 
.A(n_3971),
.B(n_792),
.Y(n_4030)
);

NOR2x1_ASAP7_75t_L g4031 ( 
.A(n_3983),
.B(n_793),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3973),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3976),
.Y(n_4033)
);

AND2x2_ASAP7_75t_L g4034 ( 
.A(n_3968),
.B(n_795),
.Y(n_4034)
);

INVxp67_ASAP7_75t_SL g4035 ( 
.A(n_3978),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_3977),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3981),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_SL g4038 ( 
.A(n_3940),
.B(n_3970),
.Y(n_4038)
);

OR2x2_ASAP7_75t_L g4039 ( 
.A(n_3989),
.B(n_799),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_3982),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_3985),
.B(n_800),
.Y(n_4041)
);

INVx2_ASAP7_75t_L g4042 ( 
.A(n_3987),
.Y(n_4042)
);

OR2x2_ASAP7_75t_L g4043 ( 
.A(n_3984),
.B(n_801),
.Y(n_4043)
);

INVxp67_ASAP7_75t_L g4044 ( 
.A(n_4001),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_4028),
.Y(n_4045)
);

NAND2xp33_ASAP7_75t_L g4046 ( 
.A(n_3998),
.B(n_802),
.Y(n_4046)
);

HB1xp67_ASAP7_75t_L g4047 ( 
.A(n_4010),
.Y(n_4047)
);

INVx2_ASAP7_75t_L g4048 ( 
.A(n_3993),
.Y(n_4048)
);

INVx2_ASAP7_75t_SL g4049 ( 
.A(n_4020),
.Y(n_4049)
);

OR2x6_ASAP7_75t_L g4050 ( 
.A(n_4006),
.B(n_803),
.Y(n_4050)
);

BUFx2_ASAP7_75t_SL g4051 ( 
.A(n_3994),
.Y(n_4051)
);

HB1xp67_ASAP7_75t_L g4052 ( 
.A(n_3996),
.Y(n_4052)
);

OAI211xp5_ASAP7_75t_L g4053 ( 
.A1(n_4038),
.A2(n_806),
.B(n_804),
.C(n_805),
.Y(n_4053)
);

NAND3xp33_ASAP7_75t_L g4054 ( 
.A(n_4014),
.B(n_804),
.C(n_805),
.Y(n_4054)
);

AOI22xp5_ASAP7_75t_L g4055 ( 
.A1(n_4019),
.A2(n_809),
.B1(n_807),
.B2(n_808),
.Y(n_4055)
);

OAI22xp5_ASAP7_75t_L g4056 ( 
.A1(n_4035),
.A2(n_812),
.B1(n_813),
.B2(n_811),
.Y(n_4056)
);

OAI21xp5_ASAP7_75t_L g4057 ( 
.A1(n_4018),
.A2(n_810),
.B(n_811),
.Y(n_4057)
);

AOI221xp5_ASAP7_75t_L g4058 ( 
.A1(n_4005),
.A2(n_813),
.B1(n_810),
.B2(n_812),
.C(n_814),
.Y(n_4058)
);

OAI22xp5_ASAP7_75t_L g4059 ( 
.A1(n_4008),
.A2(n_816),
.B1(n_817),
.B2(n_815),
.Y(n_4059)
);

AOI21xp33_ASAP7_75t_L g4060 ( 
.A1(n_4009),
.A2(n_816),
.B(n_818),
.Y(n_4060)
);

OR2x2_ASAP7_75t_L g4061 ( 
.A(n_3992),
.B(n_819),
.Y(n_4061)
);

AOI21xp5_ASAP7_75t_L g4062 ( 
.A1(n_4012),
.A2(n_819),
.B(n_820),
.Y(n_4062)
);

AOI22xp5_ASAP7_75t_SL g4063 ( 
.A1(n_4027),
.A2(n_824),
.B1(n_825),
.B2(n_823),
.Y(n_4063)
);

INVxp67_ASAP7_75t_SL g4064 ( 
.A(n_3997),
.Y(n_4064)
);

NOR2xp67_ASAP7_75t_L g4065 ( 
.A(n_4021),
.B(n_1390),
.Y(n_4065)
);

INVxp67_ASAP7_75t_L g4066 ( 
.A(n_4031),
.Y(n_4066)
);

NOR2xp33_ASAP7_75t_L g4067 ( 
.A(n_4016),
.B(n_1391),
.Y(n_4067)
);

AND2x4_ASAP7_75t_L g4068 ( 
.A(n_4015),
.B(n_825),
.Y(n_4068)
);

AOI21xp33_ASAP7_75t_L g4069 ( 
.A1(n_4024),
.A2(n_826),
.B(n_828),
.Y(n_4069)
);

INVxp67_ASAP7_75t_L g4070 ( 
.A(n_4000),
.Y(n_4070)
);

OR2x2_ASAP7_75t_L g4071 ( 
.A(n_4022),
.B(n_829),
.Y(n_4071)
);

OR2x2_ASAP7_75t_L g4072 ( 
.A(n_4026),
.B(n_829),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_4030),
.B(n_830),
.Y(n_4073)
);

BUFx2_ASAP7_75t_L g4074 ( 
.A(n_4003),
.Y(n_4074)
);

AND2x2_ASAP7_75t_L g4075 ( 
.A(n_4002),
.B(n_831),
.Y(n_4075)
);

OAI22xp33_ASAP7_75t_L g4076 ( 
.A1(n_4023),
.A2(n_836),
.B1(n_832),
.B2(n_835),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_L g4077 ( 
.A(n_4034),
.B(n_837),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_4025),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_3999),
.Y(n_4079)
);

OAI22xp33_ASAP7_75t_L g4080 ( 
.A1(n_4013),
.A2(n_841),
.B1(n_839),
.B2(n_840),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_3995),
.Y(n_4081)
);

INVxp67_ASAP7_75t_L g4082 ( 
.A(n_4004),
.Y(n_4082)
);

OAI22xp33_ASAP7_75t_L g4083 ( 
.A1(n_4011),
.A2(n_843),
.B1(n_841),
.B2(n_842),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_4017),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_4029),
.B(n_845),
.Y(n_4085)
);

AND2x2_ASAP7_75t_L g4086 ( 
.A(n_4007),
.B(n_1385),
.Y(n_4086)
);

INVxp67_ASAP7_75t_SL g4087 ( 
.A(n_4043),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_4039),
.Y(n_4088)
);

INVx2_ASAP7_75t_L g4089 ( 
.A(n_4042),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_4041),
.B(n_848),
.Y(n_4090)
);

AOI21xp5_ASAP7_75t_L g4091 ( 
.A1(n_4032),
.A2(n_851),
.B(n_852),
.Y(n_4091)
);

INVxp67_ASAP7_75t_L g4092 ( 
.A(n_4033),
.Y(n_4092)
);

INVxp33_ASAP7_75t_L g4093 ( 
.A(n_4036),
.Y(n_4093)
);

HB1xp67_ASAP7_75t_L g4094 ( 
.A(n_4037),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_4040),
.Y(n_4095)
);

INVx1_ASAP7_75t_SL g4096 ( 
.A(n_3998),
.Y(n_4096)
);

AOI21xp33_ASAP7_75t_SL g4097 ( 
.A1(n_4076),
.A2(n_853),
.B(n_854),
.Y(n_4097)
);

INVxp67_ASAP7_75t_L g4098 ( 
.A(n_4051),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_4052),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_4074),
.B(n_858),
.Y(n_4100)
);

AOI21xp33_ASAP7_75t_L g4101 ( 
.A1(n_4071),
.A2(n_1382),
.B(n_1381),
.Y(n_4101)
);

NOR3xp33_ASAP7_75t_L g4102 ( 
.A(n_4070),
.B(n_860),
.C(n_862),
.Y(n_4102)
);

AOI22xp5_ASAP7_75t_L g4103 ( 
.A1(n_4067),
.A2(n_864),
.B1(n_862),
.B2(n_863),
.Y(n_4103)
);

NAND2x1_ASAP7_75t_L g4104 ( 
.A(n_4050),
.B(n_1384),
.Y(n_4104)
);

OAI22xp5_ASAP7_75t_L g4105 ( 
.A1(n_4047),
.A2(n_4055),
.B1(n_4054),
.B2(n_4057),
.Y(n_4105)
);

INVx1_ASAP7_75t_L g4106 ( 
.A(n_4045),
.Y(n_4106)
);

OAI31xp33_ASAP7_75t_L g4107 ( 
.A1(n_4083),
.A2(n_871),
.A3(n_869),
.B(n_870),
.Y(n_4107)
);

INVx1_ASAP7_75t_SL g4108 ( 
.A(n_4063),
.Y(n_4108)
);

INVx1_ASAP7_75t_SL g4109 ( 
.A(n_4046),
.Y(n_4109)
);

OR2x2_ASAP7_75t_L g4110 ( 
.A(n_4061),
.B(n_871),
.Y(n_4110)
);

NOR3xp33_ASAP7_75t_L g4111 ( 
.A(n_4082),
.B(n_872),
.C(n_873),
.Y(n_4111)
);

AOI221x1_ASAP7_75t_L g4112 ( 
.A1(n_4060),
.A2(n_876),
.B1(n_874),
.B2(n_875),
.C(n_877),
.Y(n_4112)
);

O2A1O1Ixp33_ASAP7_75t_L g4113 ( 
.A1(n_4069),
.A2(n_1388),
.B(n_1391),
.C(n_1387),
.Y(n_4113)
);

AOI22xp5_ASAP7_75t_L g4114 ( 
.A1(n_4048),
.A2(n_880),
.B1(n_878),
.B2(n_879),
.Y(n_4114)
);

AOI221xp5_ASAP7_75t_L g4115 ( 
.A1(n_4093),
.A2(n_894),
.B1(n_898),
.B2(n_887),
.C(n_879),
.Y(n_4115)
);

O2A1O1Ixp33_ASAP7_75t_L g4116 ( 
.A1(n_4056),
.A2(n_1377),
.B(n_1378),
.C(n_1376),
.Y(n_4116)
);

OAI31xp33_ASAP7_75t_L g4117 ( 
.A1(n_4053),
.A2(n_883),
.A3(n_880),
.B(n_881),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_4068),
.B(n_4075),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_4086),
.Y(n_4119)
);

AOI22xp5_ASAP7_75t_SL g4120 ( 
.A1(n_4059),
.A2(n_886),
.B1(n_884),
.B2(n_885),
.Y(n_4120)
);

NOR2x1_ASAP7_75t_L g4121 ( 
.A(n_4072),
.B(n_4080),
.Y(n_4121)
);

AOI32xp33_ASAP7_75t_L g4122 ( 
.A1(n_4058),
.A2(n_891),
.A3(n_889),
.B1(n_890),
.B2(n_892),
.Y(n_4122)
);

A2O1A1Ixp33_ASAP7_75t_L g4123 ( 
.A1(n_4062),
.A2(n_895),
.B(n_892),
.C(n_894),
.Y(n_4123)
);

AOI21xp33_ASAP7_75t_L g4124 ( 
.A1(n_4087),
.A2(n_1380),
.B(n_1379),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_4094),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_4073),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_SL g4127 ( 
.A(n_4088),
.B(n_899),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_4077),
.Y(n_4128)
);

AOI22xp5_ASAP7_75t_L g4129 ( 
.A1(n_4081),
.A2(n_904),
.B1(n_902),
.B2(n_903),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_4085),
.Y(n_4130)
);

AOI21xp5_ASAP7_75t_L g4131 ( 
.A1(n_4091),
.A2(n_906),
.B(n_908),
.Y(n_4131)
);

AOI221xp5_ASAP7_75t_SL g4132 ( 
.A1(n_4092),
.A2(n_912),
.B1(n_910),
.B2(n_911),
.C(n_913),
.Y(n_4132)
);

INVx2_ASAP7_75t_SL g4133 ( 
.A(n_4089),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_4078),
.B(n_916),
.Y(n_4134)
);

INVx2_ASAP7_75t_L g4135 ( 
.A(n_4084),
.Y(n_4135)
);

INVx2_ASAP7_75t_L g4136 ( 
.A(n_4079),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_4090),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_4095),
.Y(n_4138)
);

AND2x4_ASAP7_75t_L g4139 ( 
.A(n_4049),
.B(n_918),
.Y(n_4139)
);

AOI21xp33_ASAP7_75t_L g4140 ( 
.A1(n_4066),
.A2(n_1381),
.B(n_1380),
.Y(n_4140)
);

OAI21xp33_ASAP7_75t_L g4141 ( 
.A1(n_4096),
.A2(n_919),
.B(n_920),
.Y(n_4141)
);

HB1xp67_ASAP7_75t_L g4142 ( 
.A(n_4065),
.Y(n_4142)
);

INVx2_ASAP7_75t_L g4143 ( 
.A(n_4049),
.Y(n_4143)
);

AOI321xp33_ASAP7_75t_L g4144 ( 
.A1(n_4064),
.A2(n_925),
.A3(n_927),
.B1(n_923),
.B2(n_924),
.C(n_926),
.Y(n_4144)
);

INVxp67_ASAP7_75t_L g4145 ( 
.A(n_4051),
.Y(n_4145)
);

INVxp67_ASAP7_75t_L g4146 ( 
.A(n_4051),
.Y(n_4146)
);

INVxp67_ASAP7_75t_L g4147 ( 
.A(n_4051),
.Y(n_4147)
);

OAI22xp33_ASAP7_75t_L g4148 ( 
.A1(n_4044),
.A2(n_931),
.B1(n_928),
.B2(n_929),
.Y(n_4148)
);

AOI222xp33_ASAP7_75t_L g4149 ( 
.A1(n_4066),
.A2(n_952),
.B1(n_936),
.B2(n_961),
.C1(n_942),
.C2(n_933),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_4052),
.Y(n_4150)
);

O2A1O1Ixp33_ASAP7_75t_L g4151 ( 
.A1(n_4047),
.A2(n_1374),
.B(n_1382),
.C(n_1373),
.Y(n_4151)
);

NOR2xp67_ASAP7_75t_SL g4152 ( 
.A(n_4051),
.B(n_934),
.Y(n_4152)
);

AOI22xp5_ASAP7_75t_L g4153 ( 
.A1(n_4044),
.A2(n_938),
.B1(n_935),
.B2(n_937),
.Y(n_4153)
);

AOI22xp5_ASAP7_75t_L g4154 ( 
.A1(n_4108),
.A2(n_1369),
.B1(n_1370),
.B2(n_1368),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_4142),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_4152),
.B(n_941),
.Y(n_4156)
);

AOI21xp5_ASAP7_75t_L g4157 ( 
.A1(n_4131),
.A2(n_944),
.B(n_945),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_4098),
.B(n_947),
.Y(n_4158)
);

NAND2x1p5_ASAP7_75t_L g4159 ( 
.A(n_4104),
.B(n_949),
.Y(n_4159)
);

INVx1_ASAP7_75t_SL g4160 ( 
.A(n_4109),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_4145),
.B(n_947),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_4146),
.B(n_949),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_4147),
.B(n_951),
.Y(n_4163)
);

AOI221x1_ASAP7_75t_L g4164 ( 
.A1(n_4099),
.A2(n_955),
.B1(n_953),
.B2(n_954),
.C(n_956),
.Y(n_4164)
);

AOI222xp33_ASAP7_75t_L g4165 ( 
.A1(n_4105),
.A2(n_960),
.B1(n_962),
.B2(n_957),
.C1(n_958),
.C2(n_961),
.Y(n_4165)
);

OAI21xp33_ASAP7_75t_L g4166 ( 
.A1(n_4143),
.A2(n_963),
.B(n_964),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_4139),
.Y(n_4167)
);

OAI21xp33_ASAP7_75t_L g4168 ( 
.A1(n_4121),
.A2(n_965),
.B(n_966),
.Y(n_4168)
);

OAI32xp33_ASAP7_75t_L g4169 ( 
.A1(n_4125),
.A2(n_976),
.A3(n_983),
.B1(n_969),
.B2(n_967),
.Y(n_4169)
);

OA21x2_ASAP7_75t_L g4170 ( 
.A1(n_4112),
.A2(n_4100),
.B(n_4134),
.Y(n_4170)
);

OAI221xp5_ASAP7_75t_SL g4171 ( 
.A1(n_4117),
.A2(n_973),
.B1(n_971),
.B2(n_972),
.C(n_975),
.Y(n_4171)
);

AOI322xp5_ASAP7_75t_L g4172 ( 
.A1(n_4132),
.A2(n_980),
.A3(n_979),
.B1(n_977),
.B2(n_971),
.C1(n_972),
.C2(n_978),
.Y(n_4172)
);

OAI21xp5_ASAP7_75t_SL g4173 ( 
.A1(n_4150),
.A2(n_981),
.B(n_982),
.Y(n_4173)
);

OAI21xp5_ASAP7_75t_SL g4174 ( 
.A1(n_4122),
.A2(n_986),
.B(n_988),
.Y(n_4174)
);

A2O1A1O1Ixp25_ASAP7_75t_L g4175 ( 
.A1(n_4144),
.A2(n_1002),
.B(n_1005),
.C(n_995),
.D(n_990),
.Y(n_4175)
);

OAI21xp33_ASAP7_75t_L g4176 ( 
.A1(n_4118),
.A2(n_990),
.B(n_991),
.Y(n_4176)
);

OAI21xp33_ASAP7_75t_L g4177 ( 
.A1(n_4119),
.A2(n_993),
.B(n_994),
.Y(n_4177)
);

AOI22xp5_ASAP7_75t_L g4178 ( 
.A1(n_4106),
.A2(n_1365),
.B1(n_1367),
.B2(n_1364),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_4097),
.B(n_996),
.Y(n_4179)
);

NOR2xp33_ASAP7_75t_L g4180 ( 
.A(n_4141),
.B(n_996),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_4110),
.Y(n_4181)
);

O2A1O1Ixp33_ASAP7_75t_L g4182 ( 
.A1(n_4151),
.A2(n_4123),
.B(n_4113),
.C(n_4140),
.Y(n_4182)
);

NAND2x1_ASAP7_75t_L g4183 ( 
.A(n_4133),
.B(n_1000),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_4149),
.B(n_4120),
.Y(n_4184)
);

NOR2xp33_ASAP7_75t_SL g4185 ( 
.A(n_4107),
.B(n_1007),
.Y(n_4185)
);

NOR2xp33_ASAP7_75t_SL g4186 ( 
.A(n_4101),
.B(n_1007),
.Y(n_4186)
);

AOI21xp5_ASAP7_75t_L g4187 ( 
.A1(n_4157),
.A2(n_4127),
.B(n_4124),
.Y(n_4187)
);

OAI21xp33_ASAP7_75t_L g4188 ( 
.A1(n_4184),
.A2(n_4130),
.B(n_4128),
.Y(n_4188)
);

OAI21xp5_ASAP7_75t_SL g4189 ( 
.A1(n_4174),
.A2(n_4126),
.B(n_4137),
.Y(n_4189)
);

O2A1O1Ixp33_ASAP7_75t_L g4190 ( 
.A1(n_4175),
.A2(n_4102),
.B(n_4116),
.C(n_4111),
.Y(n_4190)
);

OAI321xp33_ASAP7_75t_L g4191 ( 
.A1(n_4155),
.A2(n_4138),
.A3(n_4135),
.B1(n_4136),
.B2(n_4148),
.C(n_4115),
.Y(n_4191)
);

AOI221xp5_ASAP7_75t_L g4192 ( 
.A1(n_4182),
.A2(n_4153),
.B1(n_4114),
.B2(n_4129),
.C(n_4103),
.Y(n_4192)
);

OAI221xp5_ASAP7_75t_L g4193 ( 
.A1(n_4185),
.A2(n_1011),
.B1(n_1008),
.B2(n_1010),
.C(n_1012),
.Y(n_4193)
);

OAI22xp5_ASAP7_75t_L g4194 ( 
.A1(n_4154),
.A2(n_1015),
.B1(n_1013),
.B2(n_1014),
.Y(n_4194)
);

AOI22xp5_ASAP7_75t_L g4195 ( 
.A1(n_4186),
.A2(n_1018),
.B1(n_1016),
.B2(n_1017),
.Y(n_4195)
);

O2A1O1Ixp33_ASAP7_75t_L g4196 ( 
.A1(n_4171),
.A2(n_1022),
.B(n_1019),
.C(n_1020),
.Y(n_4196)
);

OAI211xp5_ASAP7_75t_L g4197 ( 
.A1(n_4172),
.A2(n_1025),
.B(n_1023),
.C(n_1024),
.Y(n_4197)
);

NOR2xp33_ASAP7_75t_L g4198 ( 
.A(n_4176),
.B(n_4177),
.Y(n_4198)
);

NAND2x1_ASAP7_75t_L g4199 ( 
.A(n_4181),
.B(n_1029),
.Y(n_4199)
);

INVx2_ASAP7_75t_SL g4200 ( 
.A(n_4183),
.Y(n_4200)
);

NAND3xp33_ASAP7_75t_SL g4201 ( 
.A(n_4165),
.B(n_1032),
.C(n_1031),
.Y(n_4201)
);

O2A1O1Ixp33_ASAP7_75t_L g4202 ( 
.A1(n_4169),
.A2(n_1035),
.B(n_1033),
.C(n_1034),
.Y(n_4202)
);

AOI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_4156),
.A2(n_1036),
.B(n_1037),
.Y(n_4203)
);

NOR2xp33_ASAP7_75t_L g4204 ( 
.A(n_4166),
.B(n_1037),
.Y(n_4204)
);

OAI221xp5_ASAP7_75t_L g4205 ( 
.A1(n_4173),
.A2(n_4158),
.B1(n_4163),
.B2(n_4162),
.C(n_4161),
.Y(n_4205)
);

AOI21xp5_ASAP7_75t_L g4206 ( 
.A1(n_4179),
.A2(n_1040),
.B(n_1041),
.Y(n_4206)
);

AOI21xp33_ASAP7_75t_SL g4207 ( 
.A1(n_4170),
.A2(n_1045),
.B(n_1044),
.Y(n_4207)
);

AOI22xp5_ASAP7_75t_L g4208 ( 
.A1(n_4180),
.A2(n_1051),
.B1(n_1049),
.B2(n_1050),
.Y(n_4208)
);

OAI21xp5_ASAP7_75t_L g4209 ( 
.A1(n_4170),
.A2(n_1056),
.B(n_1057),
.Y(n_4209)
);

AOI22xp5_ASAP7_75t_L g4210 ( 
.A1(n_4178),
.A2(n_1061),
.B1(n_1059),
.B2(n_1060),
.Y(n_4210)
);

NAND4xp25_ASAP7_75t_L g4211 ( 
.A(n_4160),
.B(n_1065),
.C(n_1063),
.D(n_1064),
.Y(n_4211)
);

AOI21xp5_ASAP7_75t_L g4212 ( 
.A1(n_4157),
.A2(n_1066),
.B(n_1067),
.Y(n_4212)
);

AOI221xp5_ASAP7_75t_L g4213 ( 
.A1(n_4168),
.A2(n_1075),
.B1(n_1072),
.B2(n_1073),
.C(n_1076),
.Y(n_4213)
);

AOI21xp5_ASAP7_75t_SL g4214 ( 
.A1(n_4164),
.A2(n_1078),
.B(n_1079),
.Y(n_4214)
);

OAI211xp5_ASAP7_75t_L g4215 ( 
.A1(n_4175),
.A2(n_1081),
.B(n_1079),
.C(n_1080),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_4167),
.Y(n_4216)
);

AOI221xp5_ASAP7_75t_L g4217 ( 
.A1(n_4168),
.A2(n_1083),
.B1(n_1080),
.B2(n_1082),
.C(n_1084),
.Y(n_4217)
);

NAND2xp5_ASAP7_75t_L g4218 ( 
.A(n_4167),
.B(n_1089),
.Y(n_4218)
);

INVx2_ASAP7_75t_L g4219 ( 
.A(n_4159),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4167),
.Y(n_4220)
);

OAI221xp5_ASAP7_75t_L g4221 ( 
.A1(n_4168),
.A2(n_1094),
.B1(n_1092),
.B2(n_1093),
.C(n_1095),
.Y(n_4221)
);

AOI221xp5_ASAP7_75t_L g4222 ( 
.A1(n_4168),
.A2(n_1098),
.B1(n_1096),
.B2(n_1097),
.C(n_1099),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_4167),
.B(n_1103),
.Y(n_4223)
);

AOI221x1_ASAP7_75t_L g4224 ( 
.A1(n_4168),
.A2(n_1107),
.B1(n_1104),
.B2(n_1106),
.C(n_1108),
.Y(n_4224)
);

OAI211xp5_ASAP7_75t_SL g4225 ( 
.A1(n_4160),
.A2(n_1110),
.B(n_1106),
.C(n_1108),
.Y(n_4225)
);

AOI21xp33_ASAP7_75t_L g4226 ( 
.A1(n_4200),
.A2(n_1114),
.B(n_1113),
.Y(n_4226)
);

OAI221xp5_ASAP7_75t_L g4227 ( 
.A1(n_4209),
.A2(n_1118),
.B1(n_1116),
.B2(n_1117),
.C(n_1119),
.Y(n_4227)
);

NOR4xp25_ASAP7_75t_L g4228 ( 
.A(n_4191),
.B(n_4188),
.C(n_4205),
.D(n_4189),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_4199),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_L g4230 ( 
.A(n_4207),
.B(n_1120),
.Y(n_4230)
);

AO22x1_ASAP7_75t_L g4231 ( 
.A1(n_4219),
.A2(n_1124),
.B1(n_1122),
.B2(n_1123),
.Y(n_4231)
);

AOI22xp5_ASAP7_75t_L g4232 ( 
.A1(n_4215),
.A2(n_1125),
.B1(n_1123),
.B2(n_1124),
.Y(n_4232)
);

A2O1A1Ixp33_ASAP7_75t_L g4233 ( 
.A1(n_4190),
.A2(n_4196),
.B(n_4202),
.C(n_4225),
.Y(n_4233)
);

OAI31xp33_ASAP7_75t_SL g4234 ( 
.A1(n_4201),
.A2(n_1130),
.A3(n_1127),
.B(n_1129),
.Y(n_4234)
);

AOI21xp33_ASAP7_75t_L g4235 ( 
.A1(n_4198),
.A2(n_1133),
.B(n_1132),
.Y(n_4235)
);

AOI21xp5_ASAP7_75t_L g4236 ( 
.A1(n_4214),
.A2(n_1134),
.B(n_1135),
.Y(n_4236)
);

OAI31xp33_ASAP7_75t_L g4237 ( 
.A1(n_4197),
.A2(n_1138),
.A3(n_1136),
.B(n_1137),
.Y(n_4237)
);

AOI21xp33_ASAP7_75t_L g4238 ( 
.A1(n_4216),
.A2(n_1141),
.B(n_1140),
.Y(n_4238)
);

AND2x2_ASAP7_75t_L g4239 ( 
.A(n_4220),
.B(n_1143),
.Y(n_4239)
);

AOI221xp5_ASAP7_75t_L g4240 ( 
.A1(n_4192),
.A2(n_1149),
.B1(n_1151),
.B2(n_1147),
.C(n_1150),
.Y(n_4240)
);

OAI22xp5_ASAP7_75t_L g4241 ( 
.A1(n_4193),
.A2(n_1155),
.B1(n_1153),
.B2(n_1154),
.Y(n_4241)
);

AOI221xp5_ASAP7_75t_L g4242 ( 
.A1(n_4187),
.A2(n_1158),
.B1(n_1160),
.B2(n_1157),
.C(n_1159),
.Y(n_4242)
);

OAI22xp5_ASAP7_75t_L g4243 ( 
.A1(n_4221),
.A2(n_4208),
.B1(n_4210),
.B2(n_4195),
.Y(n_4243)
);

OAI22xp33_ASAP7_75t_SL g4244 ( 
.A1(n_4218),
.A2(n_1172),
.B1(n_1170),
.B2(n_1171),
.Y(n_4244)
);

AOI21xp5_ASAP7_75t_L g4245 ( 
.A1(n_4212),
.A2(n_1170),
.B(n_1171),
.Y(n_4245)
);

AOI221xp5_ASAP7_75t_L g4246 ( 
.A1(n_4206),
.A2(n_1174),
.B1(n_1172),
.B2(n_1173),
.C(n_1175),
.Y(n_4246)
);

NOR2x1_ASAP7_75t_L g4247 ( 
.A(n_4211),
.B(n_1173),
.Y(n_4247)
);

AOI21xp5_ASAP7_75t_SL g4248 ( 
.A1(n_4224),
.A2(n_1174),
.B(n_1175),
.Y(n_4248)
);

AOI22xp5_ASAP7_75t_L g4249 ( 
.A1(n_4204),
.A2(n_1178),
.B1(n_1176),
.B2(n_1177),
.Y(n_4249)
);

AOI21xp5_ASAP7_75t_L g4250 ( 
.A1(n_4203),
.A2(n_1176),
.B(n_1177),
.Y(n_4250)
);

AOI221xp5_ASAP7_75t_L g4251 ( 
.A1(n_4194),
.A2(n_1363),
.B1(n_1181),
.B2(n_1179),
.C(n_1180),
.Y(n_4251)
);

NOR3xp33_ASAP7_75t_L g4252 ( 
.A(n_4223),
.B(n_1362),
.C(n_1182),
.Y(n_4252)
);

AND4x2_ASAP7_75t_L g4253 ( 
.A(n_4236),
.B(n_4217),
.C(n_4222),
.D(n_4213),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_4229),
.Y(n_4254)
);

OAI211xp5_ASAP7_75t_L g4255 ( 
.A1(n_4228),
.A2(n_4234),
.B(n_4248),
.C(n_4232),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4239),
.Y(n_4256)
);

OAI22xp5_ASAP7_75t_L g4257 ( 
.A1(n_4233),
.A2(n_1185),
.B1(n_1183),
.B2(n_1184),
.Y(n_4257)
);

AND2x2_ASAP7_75t_L g4258 ( 
.A(n_4247),
.B(n_1186),
.Y(n_4258)
);

OAI221xp5_ASAP7_75t_SL g4259 ( 
.A1(n_4237),
.A2(n_1189),
.B1(n_1187),
.B2(n_1188),
.C(n_1190),
.Y(n_4259)
);

XOR2xp5_ASAP7_75t_L g4260 ( 
.A(n_4243),
.B(n_1191),
.Y(n_4260)
);

NAND2xp5_ASAP7_75t_L g4261 ( 
.A(n_4231),
.B(n_1191),
.Y(n_4261)
);

OAI22xp5_ASAP7_75t_L g4262 ( 
.A1(n_4249),
.A2(n_1194),
.B1(n_1192),
.B2(n_1193),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4230),
.Y(n_4263)
);

AOI21xp5_ASAP7_75t_L g4264 ( 
.A1(n_4250),
.A2(n_1198),
.B(n_1199),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4244),
.Y(n_4265)
);

NOR2x1_ASAP7_75t_L g4266 ( 
.A(n_4227),
.B(n_1201),
.Y(n_4266)
);

OR2x2_ASAP7_75t_L g4267 ( 
.A(n_4241),
.B(n_1202),
.Y(n_4267)
);

O2A1O1Ixp33_ASAP7_75t_L g4268 ( 
.A1(n_4257),
.A2(n_4226),
.B(n_4238),
.C(n_4245),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_4261),
.Y(n_4269)
);

OAI211xp5_ASAP7_75t_L g4270 ( 
.A1(n_4255),
.A2(n_4240),
.B(n_4242),
.C(n_4246),
.Y(n_4270)
);

AOI211xp5_ASAP7_75t_L g4271 ( 
.A1(n_4259),
.A2(n_4235),
.B(n_4252),
.C(n_4251),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4260),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_L g4273 ( 
.A(n_4254),
.B(n_1204),
.Y(n_4273)
);

AOI22xp33_ASAP7_75t_L g4274 ( 
.A1(n_4265),
.A2(n_1207),
.B1(n_1205),
.B2(n_1206),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4258),
.Y(n_4275)
);

INVx2_ASAP7_75t_SL g4276 ( 
.A(n_4256),
.Y(n_4276)
);

INVx1_ASAP7_75t_SL g4277 ( 
.A(n_4267),
.Y(n_4277)
);

OAI222xp33_ASAP7_75t_L g4278 ( 
.A1(n_4266),
.A2(n_1215),
.B1(n_1217),
.B2(n_1213),
.C1(n_1214),
.C2(n_1216),
.Y(n_4278)
);

CKINVDCx5p33_ASAP7_75t_R g4279 ( 
.A(n_4277),
.Y(n_4279)
);

AO22x2_ASAP7_75t_L g4280 ( 
.A1(n_4276),
.A2(n_4263),
.B1(n_4264),
.B2(n_4262),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_4273),
.Y(n_4281)
);

NOR2xp33_ASAP7_75t_L g4282 ( 
.A(n_4278),
.B(n_4253),
.Y(n_4282)
);

AO22x2_ASAP7_75t_L g4283 ( 
.A1(n_4275),
.A2(n_1222),
.B1(n_1218),
.B2(n_1220),
.Y(n_4283)
);

AOI22xp5_ASAP7_75t_L g4284 ( 
.A1(n_4279),
.A2(n_4270),
.B1(n_4272),
.B2(n_4269),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4283),
.Y(n_4285)
);

AOI22xp5_ASAP7_75t_L g4286 ( 
.A1(n_4282),
.A2(n_4271),
.B1(n_4274),
.B2(n_4268),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_4280),
.Y(n_4287)
);

AOI221xp5_ASAP7_75t_L g4288 ( 
.A1(n_4287),
.A2(n_4281),
.B1(n_1225),
.B2(n_1223),
.C(n_1224),
.Y(n_4288)
);

NAND5xp2_ASAP7_75t_L g4289 ( 
.A(n_4284),
.B(n_1229),
.C(n_1226),
.D(n_1228),
.E(n_1230),
.Y(n_4289)
);

AOI222xp33_ASAP7_75t_L g4290 ( 
.A1(n_4285),
.A2(n_1233),
.B1(n_1235),
.B2(n_1231),
.C1(n_1232),
.C2(n_1234),
.Y(n_4290)
);

OAI221xp5_ASAP7_75t_L g4291 ( 
.A1(n_4286),
.A2(n_1237),
.B1(n_1235),
.B2(n_1236),
.C(n_1238),
.Y(n_4291)
);

AND3x4_ASAP7_75t_L g4292 ( 
.A(n_4289),
.B(n_1241),
.C(n_1242),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4292),
.Y(n_4293)
);

INVxp67_ASAP7_75t_SL g4294 ( 
.A(n_4293),
.Y(n_4294)
);

AOI31xp33_ASAP7_75t_SL g4295 ( 
.A1(n_4294),
.A2(n_4288),
.A3(n_4290),
.B(n_4291),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4295),
.Y(n_4296)
);

OAI21xp33_ASAP7_75t_L g4297 ( 
.A1(n_4296),
.A2(n_1243),
.B(n_1244),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_L g4298 ( 
.A(n_4297),
.B(n_1245),
.Y(n_4298)
);

AOI21xp33_ASAP7_75t_L g4299 ( 
.A1(n_4298),
.A2(n_1246),
.B(n_1247),
.Y(n_4299)
);

AOI22xp5_ASAP7_75t_L g4300 ( 
.A1(n_4299),
.A2(n_1250),
.B1(n_1247),
.B2(n_1249),
.Y(n_4300)
);

OR2x2_ASAP7_75t_L g4301 ( 
.A(n_4300),
.B(n_1251),
.Y(n_4301)
);

AOI21xp5_ASAP7_75t_L g4302 ( 
.A1(n_4301),
.A2(n_1252),
.B(n_1253),
.Y(n_4302)
);

AOI211xp5_ASAP7_75t_L g4303 ( 
.A1(n_4302),
.A2(n_1256),
.B(n_1254),
.C(n_1255),
.Y(n_4303)
);


endmodule