module fake_jpeg_30892_n_99 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_44),
.Y(n_60)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_48),
.Y(n_58)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_50),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_14),
.Y(n_50)
);

NOR2x1_ASAP7_75t_R g51 ( 
.A(n_50),
.B(n_40),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_1),
.B(n_2),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_39),
.B1(n_34),
.B2(n_37),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_54),
.B1(n_5),
.B2(n_6),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_42),
.B1(n_38),
.B2(n_35),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_37),
.B1(n_46),
.B2(n_42),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_40),
.B1(n_16),
.B2(n_17),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_46),
.B1(n_47),
.B2(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_1),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_65),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_70),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_12),
.B1(n_31),
.B2(n_29),
.Y(n_67)
);

FAx1_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_7),
.CI(n_8),
.CON(n_75),
.SN(n_75)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_58),
.B(n_3),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_73),
.B(n_7),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_5),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_6),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_9),
.B(n_10),
.Y(n_85)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_80),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_61),
.C(n_60),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_78),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_60),
.C(n_21),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_65),
.Y(n_89)
);

XNOR2x1_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_89),
.Y(n_92)
);

AO221x1_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_81),
.B1(n_76),
.B2(n_75),
.C(n_9),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_88),
.B(n_84),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_86),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_92),
.C(n_87),
.Y(n_95)
);

OAI31xp33_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_91),
.A3(n_79),
.B(n_82),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_79),
.B1(n_19),
.B2(n_20),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_11),
.C(n_22),
.Y(n_98)
);

OAI221xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.C(n_32),
.Y(n_99)
);


endmodule