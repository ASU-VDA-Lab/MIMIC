module fake_jpeg_25442_n_52 (n_3, n_2, n_1, n_0, n_4, n_5, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx11_ASAP7_75t_SL g7 ( 
.A(n_2),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx9p33_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_17),
.B(n_11),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_18),
.B(n_15),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_25),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_11),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_20),
.A2(n_12),
.B1(n_10),
.B2(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_15),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_20),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_35),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_6),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_35),
.Y(n_41)
);

OAI321xp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_43),
.A3(n_40),
.B1(n_12),
.B2(n_26),
.C(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_38),
.B1(n_10),
.B2(n_19),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_45),
.B(n_46),
.Y(n_47)
);

OAI21x1_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_3),
.B(n_5),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_1),
.C(n_21),
.Y(n_49)
);

BUFx24_ASAP7_75t_SL g51 ( 
.A(n_49),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_50),
.Y(n_52)
);


endmodule