module fake_jpeg_17022_n_285 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_285);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_34),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_41),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_29),
.A2(n_12),
.B1(n_16),
.B2(n_19),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_14),
.B1(n_21),
.B2(n_13),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_12),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_47),
.Y(n_56)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_29),
.B1(n_35),
.B2(n_30),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_37),
.B1(n_50),
.B2(n_38),
.Y(n_74)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_58),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_63),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_16),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_25),
.Y(n_62)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_21),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_38),
.B(n_15),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_68),
.A2(n_69),
.B1(n_49),
.B2(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_80),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_59),
.B1(n_42),
.B2(n_68),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_43),
.C(n_33),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_50),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_13),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_45),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_54),
.A2(n_43),
.B1(n_49),
.B2(n_37),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_82),
.A2(n_59),
.B1(n_66),
.B2(n_64),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_37),
.B(n_43),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_49),
.B1(n_28),
.B2(n_42),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_87),
.A2(n_66),
.B1(n_64),
.B2(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_61),
.B(n_14),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_62),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_101),
.B1(n_73),
.B2(n_86),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_93),
.Y(n_123)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_63),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_96),
.B1(n_76),
.B2(n_82),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_69),
.B1(n_58),
.B2(n_28),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_102),
.Y(n_128)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_78),
.B(n_26),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_71),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_103),
.B(n_109),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_43),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_105),
.A2(n_83),
.B(n_81),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_83),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_106),
.A2(n_104),
.B1(n_105),
.B2(n_95),
.Y(n_112)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_39),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_116),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_122),
.Y(n_135)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_99),
.Y(n_136)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

OAI221xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_72),
.B1(n_70),
.B2(n_75),
.C(n_80),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_75),
.A3(n_72),
.B1(n_74),
.B2(n_77),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_96),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_74),
.C(n_34),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_125),
.C(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

OAI21x1_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_43),
.B(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_73),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_34),
.C(n_43),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_105),
.B1(n_109),
.B2(n_94),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_46),
.C(n_39),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_129),
.A2(n_108),
.B1(n_86),
.B2(n_89),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_99),
.B(n_88),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_131),
.B(n_93),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_122),
.A2(n_106),
.B1(n_105),
.B2(n_96),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_132),
.A2(n_117),
.B1(n_111),
.B2(n_108),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_121),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_134),
.A2(n_110),
.B1(n_120),
.B2(n_128),
.Y(n_164)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_97),
.Y(n_137)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_153),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_92),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

NAND2x1_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_101),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_152),
.B1(n_126),
.B2(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_118),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_154),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_90),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_151),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_90),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_39),
.C(n_46),
.Y(n_153)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_108),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_127),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_150),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_128),
.C(n_116),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_160),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_162),
.B(n_22),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_164),
.A2(n_135),
.B1(n_148),
.B2(n_154),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_151),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_146),
.B(n_115),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_173),
.B(n_132),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_111),
.B1(n_24),
.B2(n_23),
.Y(n_174)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_138),
.B1(n_143),
.B2(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_68),
.B1(n_60),
.B2(n_2),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_177),
.A2(n_179),
.B1(n_169),
.B2(n_171),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_52),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_140),
.A2(n_60),
.B1(n_1),
.B2(n_2),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_153),
.C(n_135),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_156),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_187),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_150),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_161),
.C(n_165),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_189),
.A2(n_192),
.B1(n_200),
.B2(n_201),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_198),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_169),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_191),
.B(n_199),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_145),
.B1(n_155),
.B2(n_11),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_173),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_168),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_5),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_32),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_195),
.A2(n_157),
.B1(n_177),
.B2(n_166),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_203),
.B(n_207),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_166),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_205),
.A2(n_206),
.B1(n_212),
.B2(n_17),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_186),
.A2(n_161),
.B1(n_170),
.B2(n_181),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_193),
.A2(n_186),
.B1(n_199),
.B2(n_196),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_209),
.C(n_211),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_161),
.C(n_179),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_175),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_175),
.B1(n_1),
.B2(n_2),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_189),
.A2(n_8),
.B(n_11),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_213),
.A2(n_204),
.B(n_220),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_52),
.C(n_39),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_219),
.C(n_220),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_52),
.C(n_39),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_39),
.C(n_42),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_194),
.B1(n_185),
.B2(n_183),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_11),
.B1(n_9),
.B2(n_3),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_6),
.B(n_10),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_229),
.B(n_5),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_32),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_214),
.C(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_227),
.Y(n_240)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_209),
.A2(n_5),
.B(n_9),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_24),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_22),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_231),
.B(n_235),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_39),
.C(n_46),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_233),
.C(n_216),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_46),
.C(n_26),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_236),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_247),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_228),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_243),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_232),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_244),
.B(n_246),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_214),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_245),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_22),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_17),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_24),
.B(n_23),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_224),
.B(n_229),
.Y(n_251)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_252),
.A2(n_246),
.B1(n_248),
.B2(n_17),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_230),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_255),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_222),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_228),
.C(n_240),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_8),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_242),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_233),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_32),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_262),
.B(n_269),
.Y(n_273)
);

AOI322xp5_ASAP7_75t_L g272 ( 
.A1(n_263),
.A2(n_265),
.A3(n_268),
.B1(n_18),
.B2(n_46),
.C1(n_3),
.C2(n_4),
.Y(n_272)
);

AOI31xp67_ASAP7_75t_L g265 ( 
.A1(n_250),
.A2(n_245),
.A3(n_20),
.B(n_23),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_23),
.B(n_18),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_18),
.B(n_17),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_261),
.B(n_253),
.Y(n_271)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_271),
.Y(n_276)
);

NOR3xp33_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_274),
.C(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_264),
.B(n_253),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g275 ( 
.A1(n_261),
.A2(n_256),
.A3(n_18),
.B1(n_32),
.B2(n_20),
.C1(n_6),
.C2(n_9),
.Y(n_275)
);

A2O1A1O1Ixp25_ASAP7_75t_L g278 ( 
.A1(n_273),
.A2(n_256),
.B(n_20),
.C(n_4),
.D(n_5),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_278),
.B(n_6),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_276),
.A2(n_270),
.B(n_4),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_280),
.B(n_277),
.C(n_1),
.Y(n_281)
);

AOI322xp5_ASAP7_75t_L g282 ( 
.A1(n_281),
.A2(n_0),
.A3(n_1),
.B1(n_6),
.B2(n_9),
.C1(n_11),
.C2(n_243),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_282),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_283),
.B(n_0),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_0),
.C(n_273),
.Y(n_285)
);


endmodule