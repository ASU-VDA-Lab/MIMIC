module fake_jpeg_497_n_406 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_406);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_406;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_7),
.B(n_0),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_0),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_53),
.B(n_54),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_8),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_56),
.Y(n_161)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_57),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_8),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_58),
.B(n_60),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_59),
.B(n_64),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_8),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_61),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_62),
.Y(n_157)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_19),
.B(n_10),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_65),
.B(n_77),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_23),
.B(n_15),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_66),
.B(n_85),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_68),
.Y(n_172)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_69),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_22),
.A2(n_0),
.B(n_1),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_70),
.A2(n_1),
.B(n_2),
.Y(n_110)
);

CKINVDCx10_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_71),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_73),
.Y(n_173)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_74),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_40),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_17),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_21),
.B(n_12),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_86),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_45),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_88),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_52),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_90),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_21),
.B(n_31),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_93),
.Y(n_136)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_29),
.B(n_12),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_51),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_SL g165 ( 
.A(n_94),
.B(n_99),
.Y(n_165)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_100),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_104),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_31),
.B(n_12),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_103),
.Y(n_148)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_108),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_107),
.Y(n_123)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_41),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_27),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_49),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_110),
.B(n_114),
.Y(n_220)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_57),
.B(n_51),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_111),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_79),
.A2(n_46),
.B1(n_28),
.B2(n_27),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_112),
.A2(n_120),
.B1(n_128),
.B2(n_129),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_68),
.B(n_28),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_70),
.A2(n_34),
.B1(n_43),
.B2(n_50),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_71),
.A2(n_44),
.B(n_41),
.C(n_17),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_67),
.A2(n_24),
.B1(n_50),
.B2(n_33),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_67),
.A2(n_34),
.B1(n_43),
.B2(n_33),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_63),
.A2(n_32),
.B1(n_44),
.B2(n_49),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_131),
.A2(n_137),
.B1(n_145),
.B2(n_150),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_132),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_55),
.A2(n_25),
.B1(n_35),
.B2(n_32),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_133),
.A2(n_169),
.B1(n_129),
.B2(n_161),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_82),
.B(n_25),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_135),
.B(n_144),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_69),
.A2(n_35),
.B1(n_39),
.B2(n_2),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_13),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_139),
.B(n_156),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_109),
.B(n_13),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_61),
.A2(n_39),
.B1(n_3),
.B2(n_13),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_56),
.A2(n_3),
.B1(n_62),
.B2(n_72),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_80),
.B(n_86),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_164),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_84),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_90),
.B(n_106),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_160),
.B(n_121),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_97),
.B(n_104),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_92),
.A2(n_99),
.B1(n_98),
.B2(n_76),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_167),
.A2(n_177),
.B1(n_153),
.B2(n_125),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_73),
.A2(n_51),
.B1(n_58),
.B2(n_36),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_75),
.A2(n_56),
.B1(n_55),
.B2(n_72),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_170),
.A2(n_167),
.B1(n_162),
.B2(n_173),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_78),
.B(n_54),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_175),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_58),
.B(n_66),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_79),
.A2(n_67),
.B1(n_63),
.B2(n_22),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_181),
.A2(n_188),
.B1(n_193),
.B2(n_204),
.Y(n_256)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_186),
.B(n_210),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_132),
.A2(n_156),
.B1(n_123),
.B2(n_141),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_110),
.B(n_111),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_189),
.B(n_203),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_140),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_190),
.B(n_209),
.Y(n_239)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_191),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_123),
.A2(n_174),
.B1(n_158),
.B2(n_139),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_114),
.B(n_147),
.C(n_154),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_195),
.B(n_213),
.Y(n_261)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

INVx6_ASAP7_75t_SL g236 ( 
.A(n_196),
.Y(n_236)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_198),
.Y(n_268)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_199),
.Y(n_244)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_119),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_138),
.Y(n_201)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_202),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_172),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_158),
.A2(n_112),
.B1(n_115),
.B2(n_178),
.Y(n_204)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

INVx4_ASAP7_75t_SL g251 ( 
.A(n_206),
.Y(n_251)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_124),
.Y(n_207)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_207),
.Y(n_271)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_178),
.Y(n_208)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_208),
.Y(n_273)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_142),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_155),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_170),
.A2(n_150),
.B1(n_131),
.B2(n_128),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_211),
.A2(n_221),
.B1(n_126),
.B2(n_161),
.Y(n_241)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_152),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_212),
.B(n_214),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_149),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_134),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_215),
.B(n_216),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_117),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_113),
.B(n_148),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_218),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_136),
.B(n_118),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_219),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_127),
.B(n_133),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_228),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_155),
.B(n_176),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_225),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_143),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_224),
.Y(n_246)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_163),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_230),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_166),
.A2(n_137),
.B1(n_165),
.B2(n_117),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_229),
.B1(n_194),
.B2(n_179),
.Y(n_253)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_143),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_168),
.B(n_119),
.Y(n_230)
);

INVx13_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_232),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_157),
.B(n_162),
.Y(n_232)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_119),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_234),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_168),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_126),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_228),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_241),
.A2(n_258),
.B1(n_238),
.B2(n_240),
.Y(n_277)
);

AND2x6_ASAP7_75t_L g242 ( 
.A(n_185),
.B(n_157),
.Y(n_242)
);

A2O1A1O1Ixp25_ASAP7_75t_L g305 ( 
.A1(n_242),
.A2(n_243),
.B(n_274),
.C(n_247),
.D(n_266),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_189),
.A2(n_173),
.B(n_220),
.C(n_187),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_197),
.A2(n_179),
.B1(n_205),
.B2(n_211),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_245),
.B(n_253),
.Y(n_308)
);

A2O1A1Ixp33_ASAP7_75t_SL g247 ( 
.A1(n_219),
.A2(n_220),
.B(n_194),
.C(n_229),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_247),
.A2(n_259),
.B(n_198),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_220),
.B1(n_222),
.B2(n_216),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_258),
.A2(n_264),
.B1(n_259),
.B2(n_256),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_195),
.A2(n_183),
.B(n_187),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_191),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_203),
.A2(n_213),
.B1(n_182),
.B2(n_235),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_207),
.B(n_209),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_269),
.Y(n_288)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_199),
.B(n_212),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_190),
.B(n_214),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_272),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_215),
.B(n_180),
.Y(n_272)
);

AND2x6_ASAP7_75t_L g274 ( 
.A(n_206),
.B(n_196),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_269),
.Y(n_276)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_276),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_277),
.A2(n_286),
.B1(n_293),
.B2(n_303),
.Y(n_318)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_278),
.Y(n_315)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_279),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_236),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_280),
.B(n_283),
.Y(n_324)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_281),
.Y(n_317)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

NOR2x1_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_192),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_284),
.Y(n_313)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_285),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_241),
.A2(n_238),
.B1(n_243),
.B2(n_245),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_236),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_287),
.B(n_299),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_202),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_290),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_201),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_248),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_295),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_302),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_226),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_296),
.A2(n_298),
.B(n_304),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_249),
.A2(n_224),
.B(n_184),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_255),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_248),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_251),
.B(n_210),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_301),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_225),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_247),
.A2(n_208),
.B1(n_200),
.B2(n_233),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_240),
.A2(n_231),
.B1(n_260),
.B2(n_246),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_242),
.B(n_274),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_254),
.B(n_247),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_239),
.Y(n_312)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_257),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_307),
.A2(n_246),
.B1(n_291),
.B2(n_279),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_314),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_250),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_316),
.A2(n_319),
.B(n_283),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_306),
.A2(n_263),
.B(n_251),
.Y(n_319)
);

OA22x2_ASAP7_75t_L g323 ( 
.A1(n_286),
.A2(n_257),
.B1(n_273),
.B2(n_262),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_303),
.Y(n_343)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_328),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_293),
.A2(n_273),
.B1(n_268),
.B2(n_262),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_329),
.A2(n_331),
.B1(n_282),
.B2(n_285),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_276),
.A2(n_278),
.B1(n_308),
.B2(n_277),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_332),
.A2(n_349),
.B1(n_329),
.B2(n_326),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_333),
.B(n_346),
.Y(n_357)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_309),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_334),
.B(n_341),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_318),
.A2(n_308),
.B1(n_296),
.B2(n_288),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_336),
.A2(n_348),
.B1(n_315),
.B2(n_320),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_309),
.A2(n_305),
.B(n_308),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_337),
.Y(n_352)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_317),
.Y(n_338)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_338),
.Y(n_353)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_340),
.Y(n_356)
);

AO22x1_ASAP7_75t_L g341 ( 
.A1(n_324),
.A2(n_297),
.B1(n_292),
.B2(n_302),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_327),
.Y(n_342)
);

NAND3xp33_ASAP7_75t_L g360 ( 
.A(n_342),
.B(n_345),
.C(n_347),
.Y(n_360)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_343),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_311),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_344),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_310),
.B(n_290),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_319),
.A2(n_331),
.B(n_312),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_311),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_318),
.A2(n_288),
.B1(n_289),
.B2(n_295),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_316),
.A2(n_298),
.B(n_281),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_325),
.Y(n_350)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_350),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_358),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_339),
.B(n_314),
.C(n_320),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_354),
.B(n_355),
.C(n_358),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_330),
.C(n_322),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_346),
.B(n_330),
.C(n_322),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_362),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_359),
.A2(n_332),
.B1(n_336),
.B2(n_349),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_365),
.A2(n_368),
.B1(n_374),
.B2(n_362),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_360),
.B(n_341),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_367),
.B(n_369),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_352),
.A2(n_341),
.B1(n_337),
.B2(n_333),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_348),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_364),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_373),
.Y(n_379)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_363),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_372),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_SL g373 ( 
.A(n_357),
.B(n_340),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_364),
.B(n_350),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_375),
.Y(n_376)
);

XNOR2x1_ASAP7_75t_L g387 ( 
.A(n_377),
.B(n_381),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_371),
.A2(n_359),
.B1(n_351),
.B2(n_335),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_378),
.A2(n_382),
.B1(n_356),
.B2(n_353),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_368),
.A2(n_352),
.B(n_343),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_380),
.B(n_323),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_371),
.A2(n_357),
.B(n_335),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_365),
.A2(n_374),
.B1(n_361),
.B2(n_353),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_381),
.B(n_366),
.C(n_354),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_386),
.C(n_380),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_382),
.B(n_366),
.C(n_356),
.Y(n_386)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_383),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_388),
.B(n_390),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_389),
.B(n_391),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_384),
.B(n_313),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_386),
.B(n_379),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_392),
.B(n_394),
.Y(n_400)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_385),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_393),
.B(n_387),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_397),
.B(n_398),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_392),
.B(n_363),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_394),
.A2(n_376),
.B(n_387),
.Y(n_399)
);

AOI322xp5_ASAP7_75t_L g401 ( 
.A1(n_399),
.A2(n_396),
.A3(n_393),
.B1(n_395),
.B2(n_347),
.C1(n_344),
.C2(n_338),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_401),
.B(n_396),
.Y(n_403)
);

INVxp33_ASAP7_75t_L g404 ( 
.A(n_403),
.Y(n_404)
);

OAI221xp5_ASAP7_75t_L g405 ( 
.A1(n_404),
.A2(n_402),
.B1(n_400),
.B2(n_395),
.C(n_307),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_405),
.B(n_323),
.Y(n_406)
);


endmodule