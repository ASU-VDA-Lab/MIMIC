module real_aes_742_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_0), .B(n_139), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_1), .A2(n_121), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_2), .B(n_820), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_3), .A2(n_11), .B1(n_812), .B2(n_813), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_3), .Y(n_813) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_4), .B(n_129), .Y(n_185) );
INVx1_ASAP7_75t_L g126 ( .A(n_5), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_6), .B(n_129), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_7), .B(n_116), .Y(n_466) );
INVx1_ASAP7_75t_L g494 ( .A(n_8), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g820 ( .A(n_9), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_10), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_11), .Y(n_812) );
NAND2xp33_ASAP7_75t_L g166 ( .A(n_12), .B(n_133), .Y(n_166) );
INVx2_ASAP7_75t_L g118 ( .A(n_13), .Y(n_118) );
AOI221x1_ASAP7_75t_L g208 ( .A1(n_14), .A2(n_27), .B1(n_121), .B2(n_139), .C(n_209), .Y(n_208) );
CKINVDCx16_ASAP7_75t_R g429 ( .A(n_15), .Y(n_429) );
NOR3xp33_ASAP7_75t_L g818 ( .A(n_15), .B(n_819), .C(n_821), .Y(n_818) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_16), .B(n_139), .Y(n_162) );
AO21x2_ASAP7_75t_L g159 ( .A1(n_17), .A2(n_160), .B(n_161), .Y(n_159) );
INVx1_ASAP7_75t_L g475 ( .A(n_18), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_19), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_20), .B(n_152), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_21), .B(n_129), .Y(n_128) );
AO21x1_ASAP7_75t_L g180 ( .A1(n_22), .A2(n_139), .B(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g432 ( .A(n_23), .Y(n_432) );
INVx1_ASAP7_75t_L g473 ( .A(n_24), .Y(n_473) );
INVx1_ASAP7_75t_SL g459 ( .A(n_25), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_26), .B(n_140), .Y(n_553) );
NAND2x1_ASAP7_75t_L g194 ( .A(n_28), .B(n_129), .Y(n_194) );
AOI33xp33_ASAP7_75t_L g521 ( .A1(n_29), .A2(n_55), .A3(n_449), .B1(n_456), .B2(n_522), .B3(n_523), .Y(n_521) );
NAND2x1_ASAP7_75t_L g148 ( .A(n_30), .B(n_133), .Y(n_148) );
INVx1_ASAP7_75t_L g503 ( .A(n_31), .Y(n_503) );
OR2x2_ASAP7_75t_L g117 ( .A(n_32), .B(n_89), .Y(n_117) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_32), .A2(n_89), .B(n_118), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_33), .B(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_34), .B(n_133), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_35), .B(n_129), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_36), .B(n_133), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_37), .A2(n_121), .B(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g122 ( .A(n_38), .B(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g137 ( .A(n_38), .B(n_126), .Y(n_137) );
INVx1_ASAP7_75t_L g455 ( .A(n_38), .Y(n_455) );
OR2x6_ASAP7_75t_L g430 ( .A(n_39), .B(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g821 ( .A(n_39), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_40), .Y(n_505) );
XNOR2xp5_ASAP7_75t_L g775 ( .A(n_41), .B(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_42), .B(n_139), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_43), .B(n_447), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_44), .A2(n_116), .B1(n_156), .B2(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_45), .B(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_46), .A2(n_775), .B1(n_780), .B2(n_784), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_47), .B(n_140), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_48), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_49), .B(n_133), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_50), .B(n_160), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_51), .B(n_140), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_52), .A2(n_121), .B(n_147), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_53), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_54), .B(n_133), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_56), .B(n_140), .Y(n_533) );
INVx1_ASAP7_75t_L g125 ( .A(n_57), .Y(n_125) );
INVx1_ASAP7_75t_L g135 ( .A(n_57), .Y(n_135) );
AND2x2_ASAP7_75t_L g534 ( .A(n_58), .B(n_152), .Y(n_534) );
AOI221xp5_ASAP7_75t_L g492 ( .A1(n_59), .A2(n_77), .B1(n_447), .B2(n_453), .C(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_60), .B(n_447), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_61), .B(n_129), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_62), .B(n_156), .Y(n_511) );
AOI21xp5_ASAP7_75t_SL g483 ( .A1(n_63), .A2(n_453), .B(n_484), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_64), .A2(n_121), .B(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g469 ( .A(n_65), .Y(n_469) );
AO21x1_ASAP7_75t_L g182 ( .A1(n_66), .A2(n_121), .B(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_67), .B(n_139), .Y(n_170) );
INVx1_ASAP7_75t_L g532 ( .A(n_68), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_69), .B(n_139), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_70), .A2(n_453), .B(n_531), .Y(n_530) );
INVxp33_ASAP7_75t_L g824 ( .A(n_71), .Y(n_824) );
AND2x2_ASAP7_75t_L g231 ( .A(n_72), .B(n_153), .Y(n_231) );
INVx1_ASAP7_75t_L g123 ( .A(n_73), .Y(n_123) );
INVx1_ASAP7_75t_L g131 ( .A(n_73), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_74), .A2(n_99), .B1(n_777), .B2(n_778), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_74), .Y(n_777) );
AND2x2_ASAP7_75t_L g154 ( .A(n_75), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_76), .B(n_447), .Y(n_524) );
AND2x2_ASAP7_75t_L g462 ( .A(n_78), .B(n_155), .Y(n_462) );
INVx1_ASAP7_75t_L g470 ( .A(n_79), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_80), .A2(n_453), .B(n_458), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_81), .A2(n_453), .B(n_516), .C(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g433 ( .A(n_82), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_83), .B(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g168 ( .A(n_84), .B(n_155), .Y(n_168) );
AND2x2_ASAP7_75t_SL g481 ( .A(n_85), .B(n_155), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_86), .A2(n_453), .B1(n_519), .B2(n_520), .Y(n_518) );
OAI22xp5_ASAP7_75t_SL g808 ( .A1(n_87), .A2(n_809), .B1(n_810), .B2(n_811), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_87), .Y(n_809) );
AND2x2_ASAP7_75t_L g181 ( .A(n_88), .B(n_116), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_90), .B(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g198 ( .A(n_91), .B(n_155), .Y(n_198) );
INVx1_ASAP7_75t_L g485 ( .A(n_92), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_93), .B(n_129), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g120 ( .A1(n_94), .A2(n_121), .B(n_127), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_95), .B(n_133), .Y(n_210) );
AND2x2_ASAP7_75t_L g525 ( .A(n_96), .B(n_155), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_97), .B(n_129), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_98), .A2(n_501), .B(n_502), .C(n_504), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_99), .Y(n_778) );
BUFx2_ASAP7_75t_L g790 ( .A(n_100), .Y(n_790) );
BUFx2_ASAP7_75t_SL g801 ( .A(n_100), .Y(n_801) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_101), .A2(n_121), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_102), .B(n_140), .Y(n_486) );
AOI21xp33_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_814), .B(n_823), .Y(n_103) );
OA21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_787), .B(n_799), .Y(n_104) );
OAI21xp5_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_775), .B(n_779), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OAI22xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_425), .B1(n_434), .B2(n_438), .Y(n_107) );
INVx2_ASAP7_75t_L g781 ( .A(n_108), .Y(n_781) );
XNOR2x1_ASAP7_75t_L g807 ( .A(n_108), .B(n_808), .Y(n_807) );
OR2x6_ASAP7_75t_L g108 ( .A(n_109), .B(n_323), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_235), .C(n_290), .Y(n_109) );
AOI221xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_175), .B1(n_199), .B2(n_203), .C(n_213), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_158), .Y(n_111) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_112), .B(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g234 ( .A(n_112), .Y(n_234) );
AND2x2_ASAP7_75t_L g279 ( .A(n_112), .B(n_216), .Y(n_279) );
AND2x4_ASAP7_75t_L g112 ( .A(n_113), .B(n_143), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g267 ( .A(n_114), .Y(n_267) );
INVx1_ASAP7_75t_L g277 ( .A(n_114), .Y(n_277) );
AO21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_119), .B(n_141), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_115), .B(n_142), .Y(n_141) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_115), .A2(n_119), .B(n_141), .Y(n_241) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_116), .A2(n_162), .B(n_163), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_116), .B(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_116), .B(n_136), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_116), .A2(n_483), .B(n_487), .Y(n_482) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
AND2x2_ASAP7_75t_SL g153 ( .A(n_117), .B(n_118), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_138), .Y(n_119) );
AND2x6_ASAP7_75t_L g121 ( .A(n_122), .B(n_124), .Y(n_121) );
BUFx3_ASAP7_75t_L g451 ( .A(n_122), .Y(n_451) );
AND2x6_ASAP7_75t_L g133 ( .A(n_123), .B(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g457 ( .A(n_123), .Y(n_457) );
AND2x4_ASAP7_75t_L g453 ( .A(n_124), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
AND2x4_ASAP7_75t_L g129 ( .A(n_125), .B(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g449 ( .A(n_125), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_126), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_132), .B(n_136), .Y(n_127) );
INVxp67_ASAP7_75t_L g476 ( .A(n_129), .Y(n_476) );
AND2x4_ASAP7_75t_L g140 ( .A(n_130), .B(n_134), .Y(n_140) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVxp67_ASAP7_75t_L g474 ( .A(n_133), .Y(n_474) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_136), .A2(n_148), .B(n_149), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_136), .A2(n_165), .B(n_166), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_136), .A2(n_173), .B(n_174), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_136), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_136), .A2(n_194), .B(n_195), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_136), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_136), .A2(n_228), .B(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_SL g458 ( .A1(n_136), .A2(n_459), .B(n_460), .C(n_461), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_136), .A2(n_460), .B(n_485), .C(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_SL g493 ( .A1(n_136), .A2(n_460), .B(n_494), .C(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g519 ( .A(n_136), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_136), .A2(n_460), .B(n_532), .C(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_136), .A2(n_553), .B(n_554), .Y(n_552) );
INVx5_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g139 ( .A(n_137), .B(n_140), .Y(n_139) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_137), .Y(n_504) );
INVx1_ASAP7_75t_L g471 ( .A(n_140), .Y(n_471) );
OR2x2_ASAP7_75t_L g256 ( .A(n_143), .B(n_159), .Y(n_256) );
NAND2x1p5_ASAP7_75t_L g287 ( .A(n_143), .B(n_202), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_143), .B(n_167), .Y(n_300) );
INVx2_ASAP7_75t_L g309 ( .A(n_143), .Y(n_309) );
AND2x2_ASAP7_75t_L g330 ( .A(n_143), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g414 ( .A(n_143), .B(n_233), .Y(n_414) );
INVx4_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g242 ( .A(n_144), .B(n_167), .Y(n_242) );
AND2x2_ASAP7_75t_L g375 ( .A(n_144), .B(n_202), .Y(n_375) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_144), .Y(n_401) );
AO21x2_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_151), .B(n_154), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_151), .A2(n_445), .B(n_462), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_152), .A2(n_170), .B(n_171), .Y(n_169) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_152), .A2(n_208), .B(n_212), .Y(n_207) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_152), .A2(n_208), .B(n_212), .Y(n_219) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_155), .A2(n_197), .B1(n_500), .B2(n_505), .Y(n_499) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_156), .B(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx4f_ASAP7_75t_L g160 ( .A(n_157), .Y(n_160) );
AND2x4_ASAP7_75t_L g329 ( .A(n_158), .B(n_330), .Y(n_329) );
AOI321xp33_ASAP7_75t_L g343 ( .A1(n_158), .A2(n_272), .A3(n_273), .B1(n_305), .B2(n_344), .C(n_347), .Y(n_343) );
AND2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_167), .Y(n_158) );
BUFx3_ASAP7_75t_L g200 ( .A(n_159), .Y(n_200) );
INVx2_ASAP7_75t_L g233 ( .A(n_159), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_159), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g266 ( .A(n_159), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g299 ( .A(n_159), .Y(n_299) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_160), .A2(n_492), .B(n_496), .Y(n_491) );
INVx2_ASAP7_75t_SL g516 ( .A(n_160), .Y(n_516) );
INVx5_ASAP7_75t_L g202 ( .A(n_167), .Y(n_202) );
NOR2x1_ASAP7_75t_SL g251 ( .A(n_167), .B(n_241), .Y(n_251) );
BUFx2_ASAP7_75t_L g346 ( .A(n_167), .Y(n_346) );
OR2x6_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
INVxp67_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_188), .Y(n_176) );
NOR2xp33_ASAP7_75t_SL g244 ( .A(n_177), .B(n_245), .Y(n_244) );
NOR4xp25_ASAP7_75t_L g347 ( .A(n_177), .B(n_341), .C(n_345), .D(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g385 ( .A(n_177), .Y(n_385) );
AND2x2_ASAP7_75t_L g419 ( .A(n_177), .B(n_359), .Y(n_419) );
BUFx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g220 ( .A(n_178), .Y(n_220) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g274 ( .A(n_179), .Y(n_274) );
OAI21x1_ASAP7_75t_SL g179 ( .A1(n_180), .A2(n_182), .B(n_186), .Y(n_179) );
INVx1_ASAP7_75t_L g187 ( .A(n_181), .Y(n_187) );
AOI33xp33_ASAP7_75t_L g415 ( .A1(n_188), .A2(n_217), .A3(n_248), .B1(n_264), .B2(n_370), .B3(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g205 ( .A(n_189), .B(n_206), .Y(n_205) );
AND2x4_ASAP7_75t_L g215 ( .A(n_189), .B(n_216), .Y(n_215) );
BUFx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g222 ( .A(n_190), .Y(n_222) );
INVxp67_ASAP7_75t_L g303 ( .A(n_190), .Y(n_303) );
AND2x2_ASAP7_75t_L g359 ( .A(n_190), .B(n_224), .Y(n_359) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_197), .B(n_198), .Y(n_190) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_191), .A2(n_197), .B(n_198), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_192), .B(n_196), .Y(n_191) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_197), .A2(n_225), .B(n_231), .Y(n_224) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_197), .A2(n_225), .B(n_231), .Y(n_260) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_197), .A2(n_528), .B(n_534), .Y(n_527) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_197), .A2(n_528), .B(n_534), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_199), .A2(n_381), .B(n_382), .Y(n_380) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
AND2x2_ASAP7_75t_L g368 ( .A(n_200), .B(n_242), .Y(n_368) );
AND3x2_ASAP7_75t_L g370 ( .A(n_200), .B(n_254), .C(n_309), .Y(n_370) );
INVx3_ASAP7_75t_SL g322 ( .A(n_201), .Y(n_322) );
INVx4_ASAP7_75t_L g216 ( .A(n_202), .Y(n_216) );
AND2x2_ASAP7_75t_L g254 ( .A(n_202), .B(n_241), .Y(n_254) );
INVxp67_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
BUFx2_ASAP7_75t_L g248 ( .A(n_206), .Y(n_248) );
AND2x4_ASAP7_75t_L g273 ( .A(n_206), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g336 ( .A(n_206), .B(n_224), .Y(n_336) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g306 ( .A(n_207), .Y(n_306) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_207), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_R g213 ( .A1(n_214), .A2(n_217), .B(n_221), .C(n_232), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g265 ( .A(n_216), .B(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_216), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_216), .B(n_233), .Y(n_394) );
INVx1_ASAP7_75t_SL g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g376 ( .A(n_218), .B(n_366), .Y(n_376) );
AND2x2_ASAP7_75t_SL g218 ( .A(n_219), .B(n_220), .Y(n_218) );
AND2x2_ASAP7_75t_L g223 ( .A(n_219), .B(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g245 ( .A(n_219), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g261 ( .A(n_219), .B(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g294 ( .A(n_219), .B(n_274), .Y(n_294) );
AND2x4_ASAP7_75t_L g259 ( .A(n_220), .B(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g283 ( .A(n_220), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g321 ( .A(n_220), .B(n_246), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
AND2x2_ASAP7_75t_L g249 ( .A(n_222), .B(n_246), .Y(n_249) );
AND2x2_ASAP7_75t_L g264 ( .A(n_222), .B(n_224), .Y(n_264) );
BUFx2_ASAP7_75t_L g320 ( .A(n_222), .Y(n_320) );
AND2x2_ASAP7_75t_L g334 ( .A(n_222), .B(n_245), .Y(n_334) );
INVx2_ASAP7_75t_L g246 ( .A(n_224), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_226), .B(n_230), .Y(n_225) );
OAI22xp33_ASAP7_75t_L g282 ( .A1(n_232), .A2(n_283), .B1(n_285), .B2(n_289), .Y(n_282) );
INVx2_ASAP7_75t_SL g313 ( .A(n_232), .Y(n_313) );
OR2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
AND2x2_ASAP7_75t_L g288 ( .A(n_233), .B(n_241), .Y(n_288) );
INVx1_ASAP7_75t_L g395 ( .A(n_234), .Y(n_395) );
NOR3xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_268), .C(n_282), .Y(n_235) );
OAI221xp5_ASAP7_75t_SL g236 ( .A1(n_237), .A2(n_243), .B1(n_247), .B2(n_250), .C(n_252), .Y(n_236) );
INVx1_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_242), .Y(n_238) );
INVxp67_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g296 ( .A(n_240), .Y(n_296) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_240), .Y(n_424) );
INVx1_ASAP7_75t_L g387 ( .A(n_242), .Y(n_387) );
AND2x2_ASAP7_75t_SL g397 ( .A(n_242), .B(n_266), .Y(n_397) );
INVxp67_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_246), .B(n_274), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
OR2x2_ASAP7_75t_L g280 ( .A(n_248), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g358 ( .A(n_248), .Y(n_358) );
AND2x2_ASAP7_75t_L g293 ( .A(n_249), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g339 ( .A(n_251), .B(n_299), .Y(n_339) );
AND2x2_ASAP7_75t_L g416 ( .A(n_251), .B(n_414), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_257), .B1(n_264), .B2(n_265), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g275 ( .A(n_256), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_261), .Y(n_258) );
INVx2_ASAP7_75t_L g281 ( .A(n_259), .Y(n_281) );
AND2x4_ASAP7_75t_L g305 ( .A(n_259), .B(n_306), .Y(n_305) );
OAI21xp33_ASAP7_75t_SL g335 ( .A1(n_259), .A2(n_336), .B(n_337), .Y(n_335) );
AND2x2_ASAP7_75t_L g362 ( .A(n_259), .B(n_320), .Y(n_362) );
INVx2_ASAP7_75t_L g284 ( .A(n_260), .Y(n_284) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_260), .Y(n_317) );
INVx1_ASAP7_75t_SL g341 ( .A(n_261), .Y(n_341) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx2_ASAP7_75t_L g272 ( .A(n_263), .Y(n_272) );
AND2x4_ASAP7_75t_SL g366 ( .A(n_263), .B(n_284), .Y(n_366) );
AND2x2_ASAP7_75t_L g363 ( .A(n_266), .B(n_309), .Y(n_363) );
AND2x2_ASAP7_75t_L g389 ( .A(n_266), .B(n_375), .Y(n_389) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_267), .Y(n_311) );
INVx1_ASAP7_75t_L g331 ( .A(n_267), .Y(n_331) );
OAI22xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_275), .B1(n_278), .B2(n_280), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_273), .B(n_284), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_273), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g412 ( .A(n_273), .Y(n_412) );
INVx2_ASAP7_75t_SL g337 ( .A(n_275), .Y(n_337) );
AND2x2_ASAP7_75t_L g349 ( .A(n_277), .B(n_309), .Y(n_349) );
INVx2_ASAP7_75t_L g355 ( .A(n_277), .Y(n_355) );
INVxp33_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g314 ( .A(n_280), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_283), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g405 ( .A(n_283), .Y(n_405) );
INVx1_ASAP7_75t_L g333 ( .A(n_285), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_286), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g344 ( .A(n_288), .B(n_345), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_288), .A2(n_418), .B1(n_419), .B2(n_420), .Y(n_417) );
NOR3xp33_ASAP7_75t_L g290 ( .A(n_291), .B(n_312), .C(n_315), .Y(n_290) );
OAI221xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_295), .B1(n_297), .B2(n_301), .C(n_304), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_SL g410 ( .A(n_295), .Y(n_410) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g379 ( .A(n_296), .B(n_345), .Y(n_379) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g310 ( .A(n_299), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g381 ( .A(n_301), .Y(n_381) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g378 ( .A(n_302), .Y(n_378) );
INVx1_ASAP7_75t_L g384 ( .A(n_303), .Y(n_384) );
OR2x2_ASAP7_75t_L g407 ( .A(n_303), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
INVx1_ASAP7_75t_SL g316 ( .A(n_306), .Y(n_316) );
AND2x2_ASAP7_75t_L g386 ( .A(n_306), .B(n_366), .Y(n_386) );
AND2x2_ASAP7_75t_SL g418 ( .A(n_306), .B(n_319), .Y(n_418) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g423 ( .A(n_309), .Y(n_423) );
INVx1_ASAP7_75t_L g373 ( .A(n_311), .Y(n_373) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B(n_318), .C(n_322), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_316), .B(n_366), .Y(n_390) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_319), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x2_ASAP7_75t_L g327 ( .A(n_321), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g408 ( .A(n_321), .Y(n_408) );
NAND4xp75_ASAP7_75t_L g323 ( .A(n_324), .B(n_380), .C(n_396), .D(n_417), .Y(n_323) );
NOR3x1_ASAP7_75t_L g324 ( .A(n_325), .B(n_342), .C(n_364), .Y(n_324) );
NAND4xp75_ASAP7_75t_L g325 ( .A(n_326), .B(n_332), .C(n_335), .D(n_338), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_327), .B(n_329), .Y(n_326) );
AND2x2_ASAP7_75t_L g377 ( .A(n_328), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g402 ( .A(n_329), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_SL g391 ( .A(n_334), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_350), .Y(n_342) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_346), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_356), .B(n_360), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI322xp33_ASAP7_75t_L g382 ( .A1(n_354), .A2(n_383), .A3(n_387), .B1(n_388), .B2(n_390), .C1(n_391), .C2(n_392), .Y(n_382) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_355), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_358), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_359), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
OAI211xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_367), .B(n_369), .C(n_371), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_376), .B1(n_377), .B2(n_379), .Y(n_371) );
NOR2xp33_ASAP7_75t_SL g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx2_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B(n_386), .Y(n_383) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_389), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_393), .B(n_395), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g399 ( .A(n_394), .B(n_400), .Y(n_399) );
O2A1O1Ixp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B(n_403), .C(n_406), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_399), .B(n_402), .Y(n_398) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI221xp5_ASAP7_75t_SL g406 ( .A1(n_407), .A2(n_409), .B1(n_411), .B2(n_413), .C(n_415), .Y(n_406) );
INVxp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
CKINVDCx6p67_ASAP7_75t_R g425 ( .A(n_426), .Y(n_425) );
INVx4_ASAP7_75t_SL g782 ( .A(n_426), .Y(n_782) );
INVx3_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_428), .Y(n_427) );
AND2x6_ASAP7_75t_SL g428 ( .A(n_429), .B(n_430), .Y(n_428) );
OR2x6_ASAP7_75t_SL g436 ( .A(n_429), .B(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g786 ( .A(n_429), .B(n_430), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_429), .B(n_437), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_430), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_432), .B(n_433), .Y(n_822) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
CKINVDCx11_ASAP7_75t_R g435 ( .A(n_436), .Y(n_435) );
OAI22x1_ASAP7_75t_L g780 ( .A1(n_436), .A2(n_781), .B1(n_782), .B2(n_783), .Y(n_780) );
INVx1_ASAP7_75t_L g783 ( .A(n_438), .Y(n_783) );
OR3x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_640), .C(n_711), .Y(n_438) );
NAND3x1_ASAP7_75t_SL g439 ( .A(n_440), .B(n_567), .C(n_589), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_557), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_488), .B1(n_535), .B2(n_539), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_442), .A2(n_743), .B1(n_744), .B2(n_746), .Y(n_742) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_463), .Y(n_442) );
AND2x2_ASAP7_75t_L g558 ( .A(n_443), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_443), .B(n_605), .Y(n_624) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g542 ( .A(n_444), .Y(n_542) );
AND2x2_ASAP7_75t_L g592 ( .A(n_444), .B(n_465), .Y(n_592) );
INVx1_ASAP7_75t_L g631 ( .A(n_444), .Y(n_631) );
OR2x2_ASAP7_75t_L g668 ( .A(n_444), .B(n_480), .Y(n_668) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_444), .Y(n_680) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_444), .Y(n_704) );
AND2x2_ASAP7_75t_L g761 ( .A(n_444), .B(n_588), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_452), .Y(n_445) );
INVx1_ASAP7_75t_L g512 ( .A(n_447), .Y(n_512) );
AND2x4_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .Y(n_447) );
INVx1_ASAP7_75t_L g548 ( .A(n_448), .Y(n_548) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
OR2x6_ASAP7_75t_L g460 ( .A(n_449), .B(n_457), .Y(n_460) );
INVxp33_ASAP7_75t_L g522 ( .A(n_449), .Y(n_522) );
INVx1_ASAP7_75t_L g549 ( .A(n_451), .Y(n_549) );
INVxp67_ASAP7_75t_L g510 ( .A(n_453), .Y(n_510) );
NOR2x1p5_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g523 ( .A(n_456), .Y(n_523) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_460), .A2(n_469), .B1(n_470), .B2(n_471), .Y(n_468) );
INVxp67_ASAP7_75t_L g501 ( .A(n_460), .Y(n_501) );
INVx2_ASAP7_75t_L g555 ( .A(n_460), .Y(n_555) );
NOR2x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_478), .Y(n_463) );
INVx1_ASAP7_75t_L g636 ( .A(n_464), .Y(n_636) );
AND2x2_ASAP7_75t_L g662 ( .A(n_464), .B(n_480), .Y(n_662) );
NAND2x1_ASAP7_75t_L g678 ( .A(n_464), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g559 ( .A(n_465), .B(n_545), .Y(n_559) );
INVx3_ASAP7_75t_L g588 ( .A(n_465), .Y(n_588) );
NOR2x1_ASAP7_75t_SL g707 ( .A(n_465), .B(n_480), .Y(n_707) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_472), .B(n_477), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_471), .B(n_503), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B1(n_475), .B2(n_476), .Y(n_472) );
NOR2x1_ASAP7_75t_L g615 ( .A(n_478), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g586 ( .A(n_479), .B(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx4_ASAP7_75t_L g556 ( .A(n_480), .Y(n_556) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_480), .Y(n_601) );
AND2x2_ASAP7_75t_L g673 ( .A(n_480), .B(n_545), .Y(n_673) );
AND2x4_ASAP7_75t_L g690 ( .A(n_480), .B(n_634), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g737 ( .A(n_480), .B(n_632), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_480), .B(n_541), .Y(n_766) );
OR2x6_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_488), .A2(n_583), .B1(n_654), .B2(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_513), .Y(n_488) );
INVx2_ASAP7_75t_L g656 ( .A(n_489), .Y(n_656) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_497), .Y(n_489) );
BUFx3_ASAP7_75t_L g646 ( .A(n_490), .Y(n_646) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_491), .B(n_515), .Y(n_538) );
INVx2_ASAP7_75t_L g562 ( .A(n_491), .Y(n_562) );
INVx1_ASAP7_75t_L g574 ( .A(n_491), .Y(n_574) );
AND2x4_ASAP7_75t_L g581 ( .A(n_491), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g598 ( .A(n_491), .B(n_498), .Y(n_598) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_491), .Y(n_612) );
INVxp67_ASAP7_75t_L g620 ( .A(n_491), .Y(n_620) );
AND2x2_ASAP7_75t_L g649 ( .A(n_497), .B(n_565), .Y(n_649) );
AND2x2_ASAP7_75t_L g665 ( .A(n_497), .B(n_566), .Y(n_665) );
NOR2xp67_ASAP7_75t_L g752 ( .A(n_497), .B(n_565), .Y(n_752) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x4_ASAP7_75t_L g561 ( .A(n_498), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g572 ( .A(n_498), .Y(n_572) );
INVx1_ASAP7_75t_L g585 ( .A(n_498), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_498), .B(n_527), .Y(n_622) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_506), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_510), .B1(n_511), .B2(n_512), .Y(n_506) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g745 ( .A(n_513), .Y(n_745) );
AND2x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_526), .Y(n_513) );
AND2x2_ASAP7_75t_L g619 ( .A(n_514), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g648 ( .A(n_514), .Y(n_648) );
AND2x2_ASAP7_75t_L g750 ( .A(n_514), .B(n_565), .Y(n_750) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_515), .B(n_527), .Y(n_610) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B(n_525), .Y(n_515) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_516), .A2(n_517), .B(n_525), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_518), .B(n_524), .Y(n_517) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx3_ASAP7_75t_L g536 ( .A(n_526), .Y(n_536) );
NAND2x1p5_ASAP7_75t_L g725 ( .A(n_526), .B(n_646), .Y(n_725) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_527), .Y(n_639) );
AND2x2_ASAP7_75t_L g666 ( .A(n_527), .B(n_612), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
AND2x2_ASAP7_75t_L g580 ( .A(n_536), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g596 ( .A(n_536), .Y(n_596) );
AND2x2_ASAP7_75t_L g684 ( .A(n_536), .B(n_561), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_536), .B(n_704), .Y(n_709) );
AND2x2_ASAP7_75t_L g719 ( .A(n_536), .B(n_598), .Y(n_719) );
OR2x2_ASAP7_75t_L g756 ( .A(n_536), .B(n_656), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_537), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g716 ( .A(n_537), .B(n_572), .Y(n_716) );
AND2x2_ASAP7_75t_L g732 ( .A(n_537), .B(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g726 ( .A(n_538), .B(n_622), .Y(n_726) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_543), .Y(n_539) );
INVx1_ASAP7_75t_L g608 ( .A(n_540), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_540), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g706 ( .A(n_540), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_540), .B(n_587), .Y(n_731) );
INVx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_541), .Y(n_578) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_542), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_543), .A2(n_576), .B1(n_594), .B2(n_597), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_543), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_SL g710 ( .A(n_543), .Y(n_710) );
AND2x4_ASAP7_75t_SL g543 ( .A(n_544), .B(n_556), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x4_ASAP7_75t_L g587 ( .A(n_545), .B(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g607 ( .A(n_545), .Y(n_607) );
INVx1_ASAP7_75t_L g634 ( .A(n_545), .Y(n_634) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_551), .Y(n_545) );
NOR3xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .C(n_550), .Y(n_547) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_556), .Y(n_576) );
AND2x4_ASAP7_75t_L g633 ( .A(n_556), .B(n_634), .Y(n_633) );
NOR2x1_ASAP7_75t_L g694 ( .A(n_556), .B(n_663), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
AND2x2_ASAP7_75t_L g658 ( .A(n_558), .B(n_601), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g738 ( .A1(n_558), .A2(n_739), .B(n_740), .Y(n_738) );
INVx2_ASAP7_75t_L g616 ( .A(n_559), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_560), .A2(n_670), .B1(n_674), .B2(n_677), .Y(n_669) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_561), .Y(n_627) );
AND2x2_ASAP7_75t_L g637 ( .A(n_561), .B(n_638), .Y(n_637) );
INVx3_ASAP7_75t_L g676 ( .A(n_561), .Y(n_676) );
NAND2x1_ASAP7_75t_SL g701 ( .A(n_561), .B(n_570), .Y(n_701) );
AND2x2_ASAP7_75t_L g597 ( .A(n_563), .B(n_598), .Y(n_597) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NOR2x1_ASAP7_75t_L g573 ( .A(n_565), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g570 ( .A(n_566), .Y(n_570) );
INVx2_ASAP7_75t_L g582 ( .A(n_566), .Y(n_582) );
AOI21xp5_ASAP7_75t_SL g567 ( .A1(n_568), .A2(n_575), .B(n_579), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_570), .B(n_764), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_571), .A2(n_660), .B1(n_664), .B2(n_667), .Y(n_659) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
BUFx2_ASAP7_75t_L g764 ( .A(n_572), .Y(n_764) );
INVx1_ASAP7_75t_SL g771 ( .A(n_572), .Y(n_771) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_573), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OA21x2_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_583), .B(n_586), .Y(n_579) );
AND2x2_ASAP7_75t_L g583 ( .A(n_581), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g625 ( .A(n_581), .B(n_621), .Y(n_625) );
AND2x2_ASAP7_75t_L g740 ( .A(n_581), .B(n_638), .Y(n_740) );
AND2x2_ASAP7_75t_L g743 ( .A(n_581), .B(n_649), .Y(n_743) );
AND2x4_ASAP7_75t_L g751 ( .A(n_581), .B(n_752), .Y(n_751) );
OAI21xp33_ASAP7_75t_L g705 ( .A1(n_583), .A2(n_706), .B(n_708), .Y(n_705) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g733 ( .A(n_585), .Y(n_733) );
AND2x2_ASAP7_75t_L g749 ( .A(n_585), .B(n_750), .Y(n_749) );
INVx4_ASAP7_75t_L g663 ( .A(n_587), .Y(n_663) );
INVx1_ASAP7_75t_L g632 ( .A(n_588), .Y(n_632) );
AND2x2_ASAP7_75t_L g654 ( .A(n_588), .B(n_607), .Y(n_654) );
NOR2x1_ASAP7_75t_L g589 ( .A(n_590), .B(n_613), .Y(n_589) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_593), .B(n_599), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g600 ( .A(n_592), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_SL g753 ( .A(n_592), .B(n_605), .Y(n_753) );
AND2x2_ASAP7_75t_L g774 ( .A(n_592), .B(n_690), .Y(n_774) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g700 ( .A(n_597), .Y(n_700) );
OAI21xp5_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_602), .B(n_609), .Y(n_599) );
OR2x6_ASAP7_75t_L g652 ( .A(n_601), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_608), .Y(n_603) );
INVx2_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
OR2x2_ASAP7_75t_L g675 ( .A(n_610), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g772 ( .A(n_610), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_611), .B(n_745), .Y(n_744) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_626), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_617), .B1(n_623), .B2(n_625), .Y(n_614) );
OR2x2_ASAP7_75t_L g686 ( .A(n_616), .B(n_687), .Y(n_686) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_618), .Y(n_643) );
NAND2x1p5_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
INVx1_ASAP7_75t_L g692 ( .A(n_621), .Y(n_692) );
INVx2_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
INVxp67_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B1(n_635), .B2(n_637), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_633), .Y(n_629) );
AND2x4_ASAP7_75t_SL g630 ( .A(n_631), .B(n_632), .Y(n_630) );
AND2x2_ASAP7_75t_L g635 ( .A(n_633), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g696 ( .A(n_636), .B(n_690), .Y(n_696) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_641), .B(n_681), .Y(n_640) );
NOR2xp67_ASAP7_75t_L g641 ( .A(n_642), .B(n_655), .Y(n_641) );
AOI21xp33_ASAP7_75t_SL g642 ( .A1(n_643), .A2(n_644), .B(n_650), .Y(n_642) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx3_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2x1p5_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI22xp33_ASAP7_75t_SL g720 ( .A1(n_652), .A2(n_721), .B1(n_723), .B2(n_726), .Y(n_720) );
NOR2x1_ASAP7_75t_L g667 ( .A(n_653), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g703 ( .A(n_654), .B(n_704), .Y(n_703) );
OAI211xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B(n_659), .C(n_669), .Y(n_655) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp33_ASAP7_75t_SL g660 ( .A(n_661), .B(n_663), .Y(n_660) );
INVxp33_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g672 ( .A(n_663), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_664), .A2(n_684), .B1(n_685), .B2(n_688), .C(n_691), .Y(n_683) );
AND2x4_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx1_ASAP7_75t_L g724 ( .A(n_665), .Y(n_724) );
INVx2_ASAP7_75t_SL g722 ( .A(n_668), .Y(n_722) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
NAND2x1_ASAP7_75t_L g721 ( .A(n_672), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g718 ( .A(n_678), .Y(n_718) );
INVx1_ASAP7_75t_L g747 ( .A(n_679), .Y(n_747) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NOR2x1_ASAP7_75t_L g681 ( .A(n_682), .B(n_697), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_695), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g736 ( .A(n_687), .Y(n_736) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g757 ( .A(n_690), .B(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g762 ( .A(n_690), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVxp33_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
BUFx2_ASAP7_75t_L g715 ( .A(n_694), .Y(n_715) );
OAI21xp5_ASAP7_75t_SL g697 ( .A1(n_698), .A2(n_702), .B(n_705), .Y(n_697) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx2_ASAP7_75t_L g758 ( .A(n_704), .Y(n_758) );
AND2x2_ASAP7_75t_L g746 ( .A(n_707), .B(n_747), .Y(n_746) );
NOR2xp33_ASAP7_75t_R g708 ( .A(n_709), .B(n_710), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_727), .C(n_754), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_720), .Y(n_712) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_714), .B(n_717), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
OR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_728), .B(n_741), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g728 ( .A(n_729), .B(n_738), .Y(n_728) );
AOI22xp33_ASAP7_75t_SL g729 ( .A1(n_730), .A2(n_732), .B1(n_734), .B2(n_735), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NOR2x1_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVxp67_ASAP7_75t_SL g739 ( .A(n_737), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_742), .B(n_748), .Y(n_741) );
OAI21xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_751), .B(n_753), .Y(n_748) );
INVx1_ASAP7_75t_L g767 ( .A(n_751), .Y(n_767) );
AOI211xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_757), .B(n_759), .C(n_768), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_763), .B1(n_765), .B2(n_767), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_773), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
INVxp67_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
BUFx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_791), .Y(n_787) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVxp67_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g802 ( .A1(n_792), .A2(n_803), .B(n_806), .Y(n_802) );
NOR2xp33_ASAP7_75t_SL g792 ( .A(n_793), .B(n_798), .Y(n_792) );
INVx1_ASAP7_75t_SL g793 ( .A(n_794), .Y(n_793) );
BUFx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
BUFx3_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
BUFx2_ASAP7_75t_R g805 ( .A(n_797), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_802), .Y(n_799) );
INVx1_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_SL g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
INVx3_ASAP7_75t_SL g816 ( .A(n_817), .Y(n_816) );
CKINVDCx6p67_ASAP7_75t_R g827 ( .A(n_817), .Y(n_827) );
NAND2xp5_ASAP7_75t_SL g817 ( .A(n_818), .B(n_822), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
endmodule