module real_jpeg_1913_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_191;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_2),
.A2(n_82),
.B1(n_84),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_2),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_2),
.A2(n_67),
.B1(n_68),
.B2(n_110),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_110),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_110),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_4),
.B(n_84),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_4),
.B(n_111),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_4),
.A2(n_66),
.B(n_67),
.C(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_4),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_4),
.B(n_72),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_4),
.A2(n_67),
.B1(n_68),
.B2(n_160),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_4),
.B(n_31),
.C(n_34),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_160),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_4),
.B(n_45),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_4),
.B(n_60),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_5),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_5),
.A2(n_59),
.B1(n_67),
.B2(n_68),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_59),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_7),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_10),
.A2(n_81),
.B1(n_82),
.B2(n_84),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_10),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_10),
.A2(n_67),
.B1(n_68),
.B2(n_81),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_81),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_81),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_12),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_13),
.A2(n_82),
.B1(n_84),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_13),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_13),
.A2(n_67),
.B1(n_68),
.B2(n_95),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_95),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_95),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_14),
.A2(n_67),
.B1(n_68),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_14),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_75),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_75),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_15),
.A2(n_34),
.B1(n_35),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_137),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_136),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_112),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_21),
.B(n_112),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_97),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_41),
.B1(n_49),
.B2(n_50),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_33),
.B1(n_36),
.B2(n_39),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_25),
.A2(n_33),
.B1(n_153),
.B2(n_187),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_25),
.A2(n_155),
.B(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_26),
.A2(n_37),
.B1(n_58),
.B2(n_60),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_26),
.A2(n_58),
.B1(n_60),
.B2(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_26),
.A2(n_152),
.B(n_154),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_26),
.B(n_156),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

AO22x2_ASAP7_75t_L g72 ( 
.A1(n_28),
.A2(n_29),
.B1(n_66),
.B2(n_73),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_28),
.A2(n_73),
.B(n_160),
.Y(n_159)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_29),
.B(n_205),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_33),
.A2(n_175),
.B(n_176),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_33),
.A2(n_176),
.B(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_34),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_34),
.B(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_45),
.B(n_46),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_42),
.A2(n_45),
.B1(n_55),
.B2(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_42),
.A2(n_160),
.B(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_43),
.A2(n_44),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_43),
.A2(n_44),
.B1(n_134),
.B2(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_43),
.B(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_43),
.A2(n_191),
.B(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_43),
.A2(n_44),
.B1(n_191),
.B2(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_44),
.A2(n_150),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_44),
.B(n_164),
.Y(n_193)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_45),
.A2(n_163),
.B(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_61),
.B1(n_62),
.B2(n_96),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_52),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_53),
.A2(n_56),
.B1(n_57),
.B2(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_60),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_78),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_64),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_64),
.A2(n_127),
.B(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_65),
.A2(n_72),
.B1(n_126),
.B2(n_144),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B(n_71),
.C(n_72),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_67),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_68),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

AOI32xp33_ASAP7_75t_L g129 ( 
.A1(n_67),
.A2(n_82),
.A3(n_88),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_68),
.B(n_89),
.Y(n_131)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_72),
.B(n_107),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_76),
.B(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_76),
.A2(n_106),
.B(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_85),
.B(n_92),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_86),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_84),
.B1(n_88),
.B2(n_89),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_82),
.A2(n_85),
.B(n_160),
.C(n_169),
.Y(n_168)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_87),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_93),
.B(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_104),
.C(n_108),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_99),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_100),
.B(n_102),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_101),
.Y(n_175)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.C(n_119),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_113),
.B(n_117),
.Y(n_240)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_119),
.B(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_124),
.C(n_128),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_120),
.B(n_124),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_128),
.B(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_129),
.A2(n_132),
.B1(n_133),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI31xp33_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_237),
.A3(n_247),
.B(n_252),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_181),
.B(n_236),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_165),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_140),
.B(n_165),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_151),
.C(n_157),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_141),
.B(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_146),
.C(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_151),
.B(n_157),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_161),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_177),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_166),
.B(n_178),
.C(n_180),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_167),
.B(n_172),
.C(n_173),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_231),
.B(n_235),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_200),
.B(n_230),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_194),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_194),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.C(n_189),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_190),
.B1(n_209),
.B2(n_211),
.Y(n_208)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_198),
.C(n_199),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_212),
.B(n_229),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_208),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_208),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_223),
.B(n_228),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_218),
.B(n_222),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_221),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_220),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_226),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_234),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp33_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_241),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.C(n_245),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_251),
.Y(n_253)
);


endmodule