module fake_netlist_5_2141_n_70 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_70);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_70;

wire n_54;
wire n_29;
wire n_43;
wire n_47;
wire n_58;
wire n_67;
wire n_69;
wire n_36;
wire n_25;
wire n_53;
wire n_27;
wire n_42;
wire n_64;
wire n_22;
wire n_45;
wire n_24;
wire n_28;
wire n_46;
wire n_21;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_38;
wire n_61;
wire n_68;
wire n_32;
wire n_41;
wire n_35;
wire n_65;
wire n_56;
wire n_51;
wire n_63;
wire n_19;
wire n_57;
wire n_37;
wire n_59;
wire n_26;
wire n_30;
wire n_33;
wire n_55;
wire n_48;
wire n_31;
wire n_23;
wire n_50;
wire n_66;
wire n_52;
wire n_49;
wire n_60;
wire n_20;
wire n_39;

INVxp67_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NAND2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_30),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_32),
.B(n_28),
.Y(n_44)
);

OAI21x1_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_33),
.B(n_26),
.Y(n_45)
);

OAI21x1_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_33),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_43),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_43),
.B1(n_35),
.B2(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_42),
.Y(n_54)
);

AND2x4_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_39),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_33),
.B1(n_31),
.B2(n_22),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_40),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_36),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_2),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_55),
.B(n_59),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_60),
.B1(n_63),
.B2(n_62),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_60),
.B(n_56),
.Y(n_67)
);

AO21x1_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_20),
.B(n_31),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_68),
.Y(n_69)
);

NAND2x1p5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_6),
.Y(n_70)
);


endmodule