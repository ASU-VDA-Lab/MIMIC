module fake_jpeg_9138_n_209 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_209);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_33),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_19),
.B(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_14),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_47),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_21),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_29),
.B1(n_16),
.B2(n_22),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_29),
.B1(n_16),
.B2(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

OR2x2_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_31),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_56),
.Y(n_89)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_19),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_64),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_72),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_22),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_73),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_31),
.B(n_16),
.C(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_65),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_39),
.C(n_35),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_91),
.C(n_92),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_20),
.B(n_55),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_42),
.B1(n_41),
.B2(n_48),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_94),
.B1(n_20),
.B2(n_3),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_15),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_32),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_63),
.A2(n_41),
.B1(n_48),
.B2(n_26),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_62),
.A2(n_24),
.B1(n_23),
.B2(n_26),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_98),
.B1(n_66),
.B2(n_75),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_72),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_62),
.B(n_25),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_58),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_23),
.B1(n_14),
.B2(n_27),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_70),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_56),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_101),
.B(n_73),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_99),
.C(n_93),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_110),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_68),
.B1(n_52),
.B2(n_30),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_111),
.B1(n_117),
.B2(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_79),
.A2(n_57),
.B1(n_17),
.B2(n_50),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_0),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_114),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_25),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_121),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_1),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_2),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_88),
.B1(n_87),
.B2(n_113),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_125),
.C(n_135),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_78),
.C(n_84),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_139),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_130),
.B1(n_140),
.B2(n_86),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_78),
.C(n_88),
.Y(n_135)
);

OAI321xp33_ASAP7_75t_L g139 ( 
.A1(n_104),
.A2(n_82),
.A3(n_86),
.B1(n_80),
.B2(n_11),
.C(n_13),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_141),
.Y(n_150)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_111),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_87),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_151),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_146),
.A2(n_126),
.B1(n_143),
.B2(n_136),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_135),
.C(n_102),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_157),
.C(n_158),
.Y(n_162)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

XOR2x2_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_123),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_154),
.B1(n_3),
.B2(n_5),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_144),
.A2(n_112),
.B(n_118),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_134),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_137),
.A2(n_122),
.B1(n_120),
.B2(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_117),
.C(n_20),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_20),
.C(n_11),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_3),
.Y(n_161)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_167),
.C(n_173),
.Y(n_178)
);

BUFx12_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_165),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_154),
.B1(n_148),
.B2(n_150),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_127),
.C(n_126),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_127),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_174),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_129),
.C(n_10),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_158),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_162),
.C(n_167),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_150),
.B(n_160),
.Y(n_177)
);

AO21x1_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_165),
.B(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_161),
.Y(n_181)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_163),
.B(n_165),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_153),
.C(n_157),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_173),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_172),
.B(n_156),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_184),
.B(n_177),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_187),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_190),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_182),
.B(n_179),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_5),
.C(n_7),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_7),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_175),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_193),
.B(n_196),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_198),
.C(n_195),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_179),
.B1(n_8),
.B2(n_9),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_197),
.B(n_7),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_200),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_191),
.C(n_190),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_202),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_205),
.A2(n_8),
.B(n_203),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g206 ( 
.A1(n_204),
.A2(n_8),
.B(n_9),
.Y(n_206)
);

BUFx24_ASAP7_75t_SL g208 ( 
.A(n_206),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_207),
.Y(n_209)
);


endmodule