module fake_jpeg_29601_n_107 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_9),
.B(n_8),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_23),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_28),
.A2(n_34),
.B1(n_20),
.B2(n_25),
.Y(n_48)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_15),
.A2(n_22),
.B1(n_24),
.B2(n_18),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_21),
.B1(n_20),
.B2(n_25),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_3),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_36),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_12),
.A2(n_1),
.B1(n_2),
.B2(n_7),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_12),
.Y(n_35)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

AND2x6_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_35),
.B(n_31),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_17),
.B1(n_23),
.B2(n_19),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_16),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_17),
.B1(n_31),
.B2(n_7),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_16),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_4),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_63),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_59),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_31),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_64),
.C(n_65),
.Y(n_69)
);

NOR2x1_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_4),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_52),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_67),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_43),
.B(n_53),
.C(n_49),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_53),
.B(n_50),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_45),
.C(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_40),
.C(n_44),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_61),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_65),
.C(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

XNOR2x1_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_59),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_73),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_86),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_69),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_76),
.B(n_66),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_83),
.B(n_87),
.C(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_88),
.C(n_89),
.Y(n_96)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_98),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_90),
.A2(n_82),
.B(n_72),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_71),
.C(n_55),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_97),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_100),
.B(n_101),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_68),
.C(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_101),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_105),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_104),
.Y(n_107)
);


endmodule