module fake_jpeg_14023_n_432 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_432);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_432;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_48),
.Y(n_101)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_49),
.Y(n_121)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_28),
.B(n_1),
.C(n_2),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_54),
.B(n_57),
.Y(n_113)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_55),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_1),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_28),
.B(n_1),
.C(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_58),
.B(n_59),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_35),
.B(n_3),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_31),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_65),
.Y(n_112)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_16),
.B(n_3),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_67),
.B(n_75),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_70),
.Y(n_134)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_73),
.Y(n_135)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_16),
.B(n_14),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_4),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_78),
.B(n_79),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_33),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_24),
.B(n_14),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_85),
.Y(n_90)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_87),
.B1(n_21),
.B2(n_27),
.Y(n_94)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_43),
.Y(n_93)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_93),
.B(n_69),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_54),
.A2(n_41),
.B1(n_40),
.B2(n_38),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_100),
.A2(n_109),
.B1(n_119),
.B2(n_52),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_41),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_108),
.B(n_114),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_44),
.B1(n_27),
.B2(n_22),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_70),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_117),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_55),
.A2(n_18),
.B1(n_44),
.B2(n_21),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_120),
.B1(n_128),
.B2(n_138),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_36),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_51),
.B(n_36),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_81),
.A2(n_18),
.B1(n_44),
.B2(n_21),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_40),
.B1(n_38),
.B2(n_37),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_74),
.A2(n_18),
.B1(n_17),
.B2(n_22),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_48),
.B(n_37),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_4),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_52),
.B(n_32),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_115),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_77),
.A2(n_27),
.B1(n_22),
.B2(n_17),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_29),
.C(n_26),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_61),
.A2(n_17),
.B1(n_29),
.B2(n_26),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_143),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g215 ( 
.A1(n_144),
.A2(n_173),
.B1(n_180),
.B2(n_142),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_113),
.B(n_32),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_145),
.B(n_146),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_133),
.Y(n_146)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVxp67_ASAP7_75t_SL g226 ( 
.A(n_148),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_108),
.A2(n_46),
.B1(n_66),
.B2(n_72),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_149),
.A2(n_154),
.B1(n_170),
.B2(n_134),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_85),
.B1(n_88),
.B2(n_83),
.Y(n_150)
);

AO21x2_ASAP7_75t_L g233 ( 
.A1(n_150),
.A2(n_163),
.B(n_165),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_112),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_152),
.B(n_153),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_112),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_64),
.B1(n_45),
.B2(n_56),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_156),
.A2(n_170),
.B1(n_146),
.B2(n_145),
.Y(n_208)
);

AOI32xp33_ASAP7_75t_L g157 ( 
.A1(n_114),
.A2(n_85),
.A3(n_62),
.B1(n_73),
.B2(n_86),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_157),
.A2(n_161),
.B(n_156),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_102),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_158),
.B(n_159),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_123),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_160),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_174),
.Y(n_194)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

AO22x2_ASAP7_75t_L g163 ( 
.A1(n_109),
.A2(n_63),
.B1(n_60),
.B2(n_49),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_102),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_164),
.B(n_166),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_87),
.B1(n_82),
.B2(n_68),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_91),
.B(n_4),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

INVx13_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_169),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_90),
.A2(n_13),
.B1(n_6),
.B2(n_7),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

BUFx4f_ASAP7_75t_SL g203 ( 
.A(n_171),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_95),
.B1(n_97),
.B2(n_125),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_90),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_176),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_116),
.B(n_7),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_184),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_93),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_182),
.A2(n_124),
.B1(n_104),
.B2(n_142),
.Y(n_205)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_136),
.A2(n_9),
.B(n_11),
.C(n_12),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_92),
.B(n_9),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_135),
.C(n_121),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_92),
.B(n_11),
.Y(n_187)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_106),
.B(n_11),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_13),
.Y(n_213)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_127),
.B(n_12),
.Y(n_190)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_130),
.Y(n_192)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_192),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_134),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_193),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_200),
.B(n_215),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_171),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_209),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_205),
.B(n_213),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_144),
.A2(n_132),
.B1(n_126),
.B2(n_105),
.Y(n_207)
);

OA21x2_ASAP7_75t_L g266 ( 
.A1(n_207),
.A2(n_221),
.B(n_176),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_208),
.B(n_155),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_171),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_210),
.B(n_186),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g216 ( 
.A1(n_157),
.A2(n_131),
.B1(n_132),
.B2(n_105),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_219),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_149),
.A2(n_104),
.B1(n_124),
.B2(n_122),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_220),
.A2(n_229),
.B1(n_143),
.B2(n_172),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_151),
.A2(n_126),
.B1(n_122),
.B2(n_98),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_147),
.A2(n_96),
.B1(n_101),
.B2(n_121),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_121),
.C(n_135),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_181),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_178),
.B(n_103),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_188),
.Y(n_251)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_152),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_241),
.B(n_243),
.Y(n_295)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_242),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_153),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_217),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_268),
.Y(n_283)
);

OAI22x1_ASAP7_75t_SL g245 ( 
.A1(n_233),
.A2(n_151),
.B1(n_184),
.B2(n_163),
.Y(n_245)
);

A2O1A1Ixp33_ASAP7_75t_SL g292 ( 
.A1(n_245),
.A2(n_215),
.B(n_220),
.C(n_203),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_252),
.C(n_272),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_174),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_247),
.A2(n_257),
.B(n_258),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_233),
.A2(n_163),
.B1(n_159),
.B2(n_179),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_248),
.A2(n_204),
.B1(n_218),
.B2(n_236),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_250),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_256),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_SL g285 ( 
.A(n_253),
.B(n_234),
.C(n_215),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_211),
.A2(n_194),
.B(n_219),
.Y(n_254)
);

AO21x1_ASAP7_75t_L g290 ( 
.A1(n_254),
.A2(n_269),
.B(n_226),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_200),
.A2(n_233),
.B1(n_211),
.B2(n_237),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_273),
.B1(n_205),
.B2(n_233),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_161),
.Y(n_256)
);

A2O1A1O1Ixp25_ASAP7_75t_L g257 ( 
.A1(n_206),
.A2(n_166),
.B(n_185),
.C(n_186),
.D(n_163),
.Y(n_257)
);

A2O1A1O1Ixp25_ASAP7_75t_L g258 ( 
.A1(n_231),
.A2(n_163),
.B(n_182),
.C(n_148),
.D(n_115),
.Y(n_258)
);

OAI32xp33_ASAP7_75t_L g259 ( 
.A1(n_208),
.A2(n_162),
.A3(n_189),
.B1(n_168),
.B2(n_192),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_267),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_198),
.B(n_191),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_261),
.B(n_265),
.Y(n_288)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_196),
.Y(n_262)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

BUFx12_ASAP7_75t_L g263 ( 
.A(n_203),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_263),
.Y(n_286)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_197),
.Y(n_264)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_264),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_183),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_266),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_197),
.B(n_160),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_228),
.B(n_160),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_210),
.B(n_103),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_225),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_216),
.B(n_143),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_271),
.B(n_222),
.Y(n_305)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_171),
.C(n_98),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_195),
.Y(n_274)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_274),
.Y(n_306)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_236),
.Y(n_275)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_275),
.Y(n_307)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_195),
.Y(n_276)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_276),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_277),
.A2(n_279),
.B1(n_239),
.B2(n_255),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_249),
.A2(n_216),
.B1(n_215),
.B2(n_233),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_267),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_282),
.B(n_293),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_229),
.B(n_216),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_284),
.A2(n_290),
.B(n_249),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_285),
.B(n_260),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_238),
.B(n_199),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_291),
.B(n_250),
.Y(n_317)
);

AO22x1_ASAP7_75t_SL g314 ( 
.A1(n_292),
.A2(n_245),
.B1(n_249),
.B2(n_258),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_263),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_246),
.B(n_202),
.C(n_204),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_278),
.C(n_269),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_263),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_304),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_299),
.A2(n_302),
.B1(n_273),
.B2(n_242),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_271),
.A2(n_172),
.B1(n_218),
.B2(n_196),
.Y(n_302)
);

AND2x6_ASAP7_75t_L g304 ( 
.A(n_253),
.B(n_254),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_259),
.Y(n_323)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_264),
.Y(n_310)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_295),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_335),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_312),
.A2(n_327),
.B(n_300),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_283),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_313),
.B(n_321),
.Y(n_345)
);

OAI31xp33_ASAP7_75t_L g353 ( 
.A1(n_314),
.A2(n_285),
.A3(n_292),
.B(n_302),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_325),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_316),
.A2(n_329),
.B1(n_292),
.B2(n_287),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_317),
.B(n_288),
.Y(n_340)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_280),
.Y(n_320)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_320),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_278),
.B(n_252),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_322),
.B(n_326),
.C(n_328),
.Y(n_347)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_323),
.Y(n_352)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_324),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_281),
.B(n_251),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_296),
.A2(n_260),
.B(n_247),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_281),
.B(n_269),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_294),
.A2(n_266),
.B1(n_240),
.B2(n_257),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_256),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_332),
.C(n_333),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_272),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_290),
.B(n_275),
.C(n_276),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_277),
.A2(n_266),
.B1(n_262),
.B2(n_270),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_337),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_288),
.B(n_274),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_301),
.B(n_230),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_338),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_279),
.A2(n_225),
.B1(n_222),
.B2(n_224),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_290),
.B(n_223),
.Y(n_338)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_340),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_322),
.B(n_301),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_348),
.C(n_326),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_323),
.A2(n_294),
.B1(n_284),
.B2(n_305),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_342),
.A2(n_343),
.B1(n_334),
.B2(n_337),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_332),
.B(n_304),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_330),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_350),
.B(n_336),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_353),
.A2(n_361),
.B(n_312),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_286),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_354),
.B(n_357),
.Y(n_377)
);

OAI221xp5_ASAP7_75t_L g355 ( 
.A1(n_327),
.A2(n_310),
.B1(n_300),
.B2(n_287),
.C(n_292),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_355),
.A2(n_333),
.B1(n_338),
.B2(n_316),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_319),
.B(n_293),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_318),
.Y(n_358)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_358),
.Y(n_367)
);

INVx5_ASAP7_75t_L g360 ( 
.A(n_319),
.Y(n_360)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_360),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_375),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_363),
.A2(n_361),
.B(n_353),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_331),
.C(n_328),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_368),
.C(n_370),
.Y(n_384)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_365),
.Y(n_383)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_366),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_347),
.B(n_321),
.C(n_314),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_351),
.B(n_314),
.C(n_298),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_286),
.C(n_292),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_371),
.B(n_380),
.C(n_344),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_307),
.Y(n_372)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_372),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_373),
.A2(n_359),
.B1(n_352),
.B2(n_360),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_346),
.A2(n_307),
.B1(n_309),
.B2(n_306),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_374),
.A2(n_379),
.B1(n_358),
.B2(n_356),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_344),
.B(n_309),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_306),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_356),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_346),
.A2(n_289),
.B1(n_308),
.B2(n_303),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_341),
.B(n_303),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_385),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_377),
.B(n_340),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_386),
.B(n_395),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_364),
.B(n_345),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_396),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_388),
.A2(n_393),
.B(n_394),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_389),
.A2(n_390),
.B1(n_392),
.B2(n_378),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_378),
.A2(n_359),
.B1(n_379),
.B2(n_342),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_363),
.Y(n_393)
);

NOR2x1_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_348),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_374),
.B(n_349),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_384),
.B(n_370),
.C(n_371),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_401),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_387),
.B(n_369),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_384),
.B(n_362),
.C(n_368),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_402),
.B(n_404),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_403),
.A2(n_391),
.B1(n_392),
.B2(n_394),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_381),
.B(n_375),
.C(n_380),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_381),
.B(n_366),
.C(n_372),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_406),
.B(n_383),
.C(n_393),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_396),
.B(n_289),
.Y(n_407)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_407),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_L g408 ( 
.A(n_402),
.B(n_382),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_408),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_400),
.A2(n_383),
.B1(n_373),
.B2(n_388),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_413),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_399),
.A2(n_405),
.B(n_397),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_412),
.A2(n_415),
.B1(n_416),
.B2(n_367),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_398),
.A2(n_395),
.B(n_385),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_409),
.B(n_400),
.C(n_406),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_421),
.Y(n_423)
);

NOR2x1_ASAP7_75t_SL g425 ( 
.A(n_418),
.B(n_419),
.Y(n_425)
);

AOI221xp5_ASAP7_75t_L g419 ( 
.A1(n_414),
.A2(n_367),
.B1(n_355),
.B2(n_339),
.C(n_263),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_339),
.C(n_224),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_422),
.A2(n_415),
.B1(n_410),
.B2(n_411),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_424),
.B(n_203),
.C(n_223),
.Y(n_428)
);

NOR2x1_ASAP7_75t_L g426 ( 
.A(n_417),
.B(n_421),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_426),
.A2(n_420),
.B(n_308),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_427),
.B(n_428),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_429),
.B(n_426),
.Y(n_430)
);

AO21x1_ASAP7_75t_L g431 ( 
.A1(n_430),
.A2(n_423),
.B(n_425),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_431),
.B(n_230),
.Y(n_432)
);


endmodule