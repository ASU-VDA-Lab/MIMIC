module fake_jpeg_17323_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_30),
.Y(n_55)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_29),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_70),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_77),
.Y(n_84)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_31),
.B1(n_39),
.B2(n_38),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_64),
.B1(n_53),
.B2(n_33),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_31),
.B1(n_39),
.B2(n_38),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_26),
.B1(n_28),
.B2(n_24),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_73),
.B(n_81),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_0),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_44),
.B(n_33),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_23),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_17),
.B(n_15),
.C(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_24),
.Y(n_74)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_23),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_47),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_28),
.B1(n_15),
.B2(n_16),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_17),
.B1(n_27),
.B2(n_20),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_85),
.A2(n_110),
.B1(n_45),
.B2(n_34),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_52),
.C(n_47),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_52),
.C(n_47),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_62),
.B(n_58),
.CI(n_67),
.CON(n_90),
.SN(n_90)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_60),
.Y(n_113)
);

INVx5_ASAP7_75t_SL g96 ( 
.A(n_75),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_96),
.A2(n_99),
.B1(n_53),
.B2(n_56),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_64),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_61),
.A2(n_20),
.B1(n_19),
.B2(n_16),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_79),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_106),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_0),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_107),
.A2(n_108),
.B(n_97),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_0),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_69),
.A2(n_39),
.B1(n_33),
.B2(n_34),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g111 ( 
.A1(n_70),
.A2(n_19),
.B(n_18),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_73),
.C(n_29),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_112),
.B(n_123),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_132),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_137),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_69),
.Y(n_121)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_80),
.B1(n_68),
.B2(n_33),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_85),
.B1(n_96),
.B2(n_110),
.Y(n_142)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_126),
.A2(n_133),
.B1(n_93),
.B2(n_34),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_68),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_130),
.Y(n_144)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_45),
.Y(n_130)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_131),
.A2(n_115),
.B1(n_129),
.B2(n_128),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_94),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_59),
.Y(n_135)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_76),
.C(n_40),
.Y(n_168)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_53),
.B(n_23),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_93),
.B1(n_108),
.B2(n_98),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_140),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_142),
.A2(n_146),
.B1(n_149),
.B2(n_34),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_112),
.A2(n_95),
.B1(n_92),
.B2(n_86),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_104),
.B(n_108),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_147),
.A2(n_25),
.B1(n_29),
.B2(n_35),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_137),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_160),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_97),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_117),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_123),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_168),
.C(n_32),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_125),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_114),
.B(n_107),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_23),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_164),
.A2(n_131),
.B1(n_139),
.B2(n_115),
.Y(n_174)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_116),
.A2(n_107),
.B1(n_98),
.B2(n_34),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_138),
.B(n_119),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_122),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_76),
.Y(n_169)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_132),
.B(n_29),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_170),
.B(n_18),
.Y(n_198)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_172),
.A2(n_176),
.B(n_188),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_149),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_195),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_168),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_18),
.Y(n_180)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_163),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_182),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_163),
.Y(n_182)
);

AO21x2_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_82),
.B(n_43),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_183),
.A2(n_153),
.B1(n_156),
.B2(n_157),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_189),
.C(n_148),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_23),
.Y(n_185)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_29),
.Y(n_187)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_38),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_18),
.Y(n_191)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_144),
.A2(n_38),
.B(n_25),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_193),
.A2(n_194),
.B(n_197),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_151),
.A2(n_35),
.B1(n_43),
.B2(n_42),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_150),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_200),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_167),
.A2(n_40),
.B(n_32),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_198),
.B(n_141),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g200 ( 
.A1(n_154),
.A2(n_40),
.A3(n_32),
.B1(n_3),
.B2(n_4),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_155),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_203),
.A2(n_159),
.B(n_161),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_204),
.A2(n_213),
.B1(n_183),
.B2(n_200),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_184),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_216),
.C(n_223),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_175),
.Y(n_206)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_183),
.B1(n_190),
.B2(n_174),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_210),
.B(n_222),
.Y(n_248)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_173),
.Y(n_212)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_166),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_148),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_2),
.C(n_5),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_162),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_195),
.C(n_203),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_226),
.B(n_208),
.Y(n_249)
);

MAJx2_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_147),
.C(n_177),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_239),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_172),
.B(n_193),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_233),
.A2(n_226),
.B(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_211),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_217),
.Y(n_252)
);

XOR2x2_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_147),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_243),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_187),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_240),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_195),
.B1(n_197),
.B2(n_194),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_241),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_195),
.C(n_40),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_247),
.C(n_204),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_216),
.B(n_1),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_225),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_249),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_253),
.Y(n_269)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_230),
.Y(n_254)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_256),
.B(n_258),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_248),
.B(n_209),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_232),
.B(n_224),
.Y(n_260)
);

NOR2xp67_ASAP7_75t_R g274 ( 
.A(n_260),
.B(n_245),
.Y(n_274)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_246),
.B(n_6),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_235),
.A2(n_218),
.B1(n_221),
.B2(n_219),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_265),
.C(n_247),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_235),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_264),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_212),
.C(n_6),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_253),
.B(n_257),
.Y(n_281)
);

XNOR2x1_ASAP7_75t_SL g268 ( 
.A(n_251),
.B(n_238),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_268),
.B(n_249),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_237),
.C(n_255),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_273),
.C(n_9),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_275),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_237),
.C(n_244),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_250),
.B1(n_263),
.B2(n_262),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_243),
.C(n_231),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_5),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_256),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_286),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_283),
.B(n_288),
.Y(n_296)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_264),
.B(n_7),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_287),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_5),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_14),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_7),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_8),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_290),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_8),
.B(n_9),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_266),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_295),
.B(n_298),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_270),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_279),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_9),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_286),
.B(n_276),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_10),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_291),
.B(n_273),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_301),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_303),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_10),
.Y(n_303)
);

MAJx2_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_306),
.C(n_307),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_13),
.Y(n_307)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_308),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_311),
.A2(n_302),
.B(n_304),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_310),
.C(n_297),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_293),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_314),
.B(n_309),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_294),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_14),
.Y(n_317)
);


endmodule