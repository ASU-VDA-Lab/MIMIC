module fake_netlist_1_7060_n_23 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_23);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_23;
wire n_20;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
wire n_21;
CKINVDCx20_ASAP7_75t_R g11 ( .A(n_4), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_0), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_0), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_6), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_12), .Y(n_15) );
A2O1A1Ixp33_ASAP7_75t_L g16 ( .A1(n_13), .A2(n_1), .B(n_2), .C(n_3), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_15), .B(n_14), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_17), .B(n_11), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
AOI221xp5_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_16), .B1(n_11), .B2(n_3), .C(n_1), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
OAI22xp5_ASAP7_75t_SL g22 ( .A1(n_21), .A2(n_2), .B1(n_5), .B2(n_7), .Y(n_22) );
AOI22xp33_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_23) );
endmodule