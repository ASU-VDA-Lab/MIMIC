module fake_jpeg_3363_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_59),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_58),
.Y(n_60)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_48),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_65),
.B(n_50),
.C(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_47),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_42),
.B1(n_41),
.B2(n_43),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_68),
.A2(n_42),
.B1(n_47),
.B2(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

AO22x1_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_57),
.B1(n_40),
.B2(n_49),
.Y(n_73)
);

NOR2x1_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_64),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_80),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_79),
.Y(n_91)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_46),
.Y(n_79)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_83),
.Y(n_89)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp67_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_98),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_50),
.B(n_4),
.Y(n_100)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_17),
.Y(n_93)
);

A2O1A1O1Ixp25_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_20),
.B(n_33),
.C(n_31),
.D(n_29),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_97),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_1),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_2),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_102),
.Y(n_123)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_18),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_3),
.B(n_4),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_114),
.B(n_10),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_3),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_110),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_93),
.B1(n_90),
.B2(n_9),
.Y(n_116)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_5),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_113),
.A2(n_25),
.B1(n_27),
.B2(n_16),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_111),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_24),
.B(n_28),
.C(n_12),
.D(n_15),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_125),
.B1(n_107),
.B2(n_23),
.Y(n_132)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_128),
.Y(n_133)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_130),
.B1(n_132),
.B2(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_99),
.C(n_100),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_126),
.C(n_120),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_134),
.A2(n_120),
.B(n_118),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_131),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_137),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_135),
.B1(n_133),
.B2(n_106),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_122),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_26),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_36),
.B(n_10),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);


endmodule