module fake_jpeg_1812_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_28),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_45),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_49),
.B(n_55),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_53),
.B(n_35),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_41),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_48),
.B(n_46),
.C(n_40),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_49),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_46),
.B1(n_44),
.B2(n_37),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_64),
.B1(n_1),
.B2(n_2),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_55),
.A2(n_43),
.B1(n_37),
.B2(n_39),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_54),
.B1(n_52),
.B2(n_3),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_43),
.B1(n_39),
.B2(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_50),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_5),
.B(n_6),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_17),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_71),
.Y(n_82)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_54),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_78),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_4),
.Y(n_80)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_75),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_80),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_89),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_90),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_57),
.B(n_8),
.Y(n_85)
);

OA21x2_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_9),
.B(n_10),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_70),
.A2(n_20),
.B1(n_33),
.B2(n_31),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_22),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_7),
.B(n_8),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_7),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_73),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_9),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_107),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_21),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_99),
.C(n_13),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_104),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_87),
.C(n_85),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_103),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_12),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_12),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_114),
.C(n_117),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_16),
.C(n_19),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_23),
.B(n_25),
.Y(n_115)
);

NAND2xp33_ASAP7_75t_SL g120 ( 
.A(n_115),
.B(n_101),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_30),
.Y(n_117)
);

XOR2x2_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_34),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_98),
.C(n_103),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_109),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_121)
);

AO21x1_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_109),
.B(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_123),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_118),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_119),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_124),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_126),
.Y(n_131)
);


endmodule