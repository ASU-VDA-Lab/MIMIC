module fake_jpeg_14255_n_93 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_93);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_93;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_0),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_1),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_33),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_13),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_24),
.A2(n_29),
.B1(n_13),
.B2(n_19),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_16),
.B(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_30),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_19),
.A2(n_2),
.B1(n_3),
.B2(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_18),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_21),
.B1(n_31),
.B2(n_10),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_21),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_10),
.Y(n_61)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_23),
.B(n_24),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_34),
.B(n_41),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_54),
.B1(n_48),
.B2(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_37),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_10),
.B1(n_18),
.B2(n_26),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_59),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g57 ( 
.A(n_45),
.B(n_30),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_37),
.C(n_47),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_38),
.B(n_36),
.Y(n_60)
);

A2O1A1O1Ixp25_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_52),
.B(n_49),
.C(n_53),
.D(n_61),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_41),
.B(n_42),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_63),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_69),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_65),
.B(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_58),
.C(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_42),
.Y(n_69)
);

AOI22x1_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_48),
.B1(n_58),
.B2(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_73),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_61),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_78),
.B1(n_68),
.B2(n_69),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_82),
.B(n_74),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_62),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_83),
.A2(n_77),
.B1(n_81),
.B2(n_78),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_83),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_75),
.B1(n_71),
.B2(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_67),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_82),
.C(n_80),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_79),
.C(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_89),
.B(n_90),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_91),
.Y(n_92)
);

AOI221xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_88),
.B1(n_79),
.B2(n_8),
.C(n_51),
.Y(n_93)
);


endmodule