module fake_jpeg_28229_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_38),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_16),
.Y(n_53)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_44),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_0),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_30),
.Y(n_60)
);

CKINVDCx9p33_ASAP7_75t_R g46 ( 
.A(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_48),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_49),
.B(n_50),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_62),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_64),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NAND2x1_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_17),
.Y(n_61)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_46),
.Y(n_85)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_26),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_41),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_21),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_17),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_81),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_85),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_45),
.B1(n_26),
.B2(n_22),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_71),
.A2(n_78),
.B1(n_83),
.B2(n_94),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_26),
.B1(n_25),
.B2(n_32),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_25),
.B1(n_32),
.B2(n_18),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_76),
.A2(n_86),
.B1(n_47),
.B2(n_58),
.Y(n_123)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_25),
.B1(n_32),
.B2(n_35),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_79),
.B(n_80),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_65),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_35),
.B1(n_23),
.B2(n_19),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_23),
.B1(n_19),
.B2(n_29),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_90),
.B1(n_93),
.B2(n_98),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_18),
.B1(n_23),
.B2(n_27),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_87),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_38),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_23),
.B1(n_19),
.B2(n_29),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_42),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_47),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_29),
.B1(n_39),
.B2(n_33),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_27),
.B1(n_30),
.B2(n_39),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_52),
.A2(n_39),
.B1(n_30),
.B2(n_41),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_62),
.B1(n_47),
.B2(n_28),
.Y(n_130)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_42),
.C(n_61),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_58),
.C(n_52),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_61),
.A2(n_42),
.B(n_38),
.C(n_17),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_20),
.B(n_28),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_17),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_113),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_58),
.B1(n_52),
.B2(n_62),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_130),
.B1(n_95),
.B2(n_75),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_68),
.B(n_39),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_109),
.B(n_129),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_79),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_69),
.B(n_56),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_71),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_122),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_99),
.B(n_20),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_128),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_85),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_24),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_69),
.B(n_28),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_112),
.B(n_106),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_133),
.A2(n_137),
.B(n_138),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_121),
.A2(n_97),
.B1(n_85),
.B2(n_74),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_136),
.B(n_48),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_100),
.B(n_98),
.C(n_74),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_68),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_139),
.B(n_159),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_87),
.B(n_98),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_146),
.B(n_149),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_73),
.B(n_87),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_70),
.B1(n_87),
.B2(n_93),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_73),
.B1(n_90),
.B2(n_84),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_83),
.B(n_88),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_160),
.Y(n_182)
);

OR2x4_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_101),
.Y(n_148)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_109),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_88),
.B(n_101),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_88),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_48),
.B(n_17),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_116),
.A2(n_92),
.B1(n_77),
.B2(n_89),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_152),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_107),
.A2(n_92),
.B1(n_75),
.B2(n_33),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_154),
.B1(n_104),
.B2(n_108),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_102),
.A2(n_118),
.B1(n_125),
.B2(n_114),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_48),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_102),
.A2(n_34),
.B(n_33),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_0),
.Y(n_192)
);

XOR2x1_ASAP7_75t_SL g206 ( 
.A(n_165),
.B(n_149),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_138),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_167),
.B(n_168),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_108),
.Y(n_168)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_170),
.Y(n_216)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_172),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_157),
.B(n_129),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_178),
.B1(n_180),
.B2(n_145),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_111),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_175),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_111),
.C(n_117),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_186),
.C(n_191),
.Y(n_208)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_183),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_159),
.A2(n_117),
.B1(n_75),
.B2(n_34),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_147),
.A2(n_34),
.B1(n_20),
.B2(n_48),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_181),
.A2(n_140),
.B(n_142),
.Y(n_223)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_193),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_187),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_48),
.C(n_17),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_24),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_139),
.B(n_24),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_189),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_17),
.C(n_16),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_194),
.Y(n_200)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_131),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_132),
.B(n_0),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_135),
.B(n_16),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_176),
.C(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_198),
.B(n_201),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_164),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_182),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_150),
.B1(n_144),
.B2(n_153),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_202),
.A2(n_204),
.B1(n_225),
.B2(n_188),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_150),
.B1(n_138),
.B2(n_143),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_182),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_205),
.B(n_211),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_162),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_173),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_137),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_215),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_187),
.C(n_166),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_191),
.C(n_186),
.Y(n_226)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_217),
.B(n_219),
.Y(n_230)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_158),
.Y(n_221)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_223),
.A2(n_173),
.B(n_188),
.Y(n_229)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_224),
.B(n_198),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_166),
.A2(n_134),
.B1(n_133),
.B2(n_146),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_226),
.B(n_228),
.Y(n_263)
);

AO22x1_ASAP7_75t_L g227 ( 
.A1(n_212),
.A2(n_165),
.B1(n_179),
.B2(n_167),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_233),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_229),
.A2(n_240),
.B(n_200),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_236),
.B1(n_217),
.B2(n_225),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_232),
.A2(n_210),
.B1(n_207),
.B2(n_200),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_170),
.C(n_163),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_194),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_235),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_204),
.A2(n_134),
.B1(n_193),
.B2(n_3),
.Y(n_236)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_8),
.C(n_13),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_241),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_197),
.A2(n_1),
.B(n_2),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_218),
.B(n_14),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_14),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_245),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_213),
.C(n_206),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_248),
.A2(n_202),
.B1(n_197),
.B2(n_201),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_250),
.A2(n_251),
.B1(n_258),
.B2(n_269),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_248),
.A2(n_205),
.B1(n_199),
.B2(n_215),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_253),
.A2(n_261),
.B(n_227),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_255),
.A2(n_266),
.B1(n_230),
.B2(n_239),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_243),
.A2(n_223),
.B1(n_211),
.B2(n_214),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_221),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_268),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_242),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_12),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_231),
.A2(n_224),
.B1(n_219),
.B2(n_3),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_12),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_243),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_229),
.B(n_240),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_272),
.Y(n_298)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_236),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_273),
.A2(n_280),
.B(n_269),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_245),
.C(n_228),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_260),
.C(n_257),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_234),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_285),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_238),
.Y(n_277)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_277),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_255),
.A2(n_235),
.B1(n_244),
.B2(n_9),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_279),
.A2(n_10),
.B1(n_11),
.B2(n_6),
.Y(n_293)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_281),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_267),
.B(n_12),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_284),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_266),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_283),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_297)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_8),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_256),
.B1(n_259),
.B2(n_252),
.Y(n_286)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_286),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_273),
.C(n_278),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_257),
.C(n_268),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_275),
.C(n_285),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_264),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_292),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_291),
.A2(n_296),
.B1(n_270),
.B2(n_278),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_258),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_293),
.A2(n_297),
.B1(n_283),
.B2(n_271),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_303),
.C(n_304),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_305),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_281),
.C(n_10),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_298),
.A2(n_10),
.B(n_11),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_308),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_299),
.Y(n_307)
);

NOR2x1_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_301),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_295),
.C(n_292),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_287),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_297),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_315),
.Y(n_321)
);

AO21x2_ASAP7_75t_SL g316 ( 
.A1(n_309),
.A2(n_295),
.B(n_290),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_316),
.A2(n_7),
.B1(n_308),
.B2(n_311),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_7),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_318),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_7),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_322),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_318),
.Y(n_320)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_314),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_316),
.C(n_319),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_324),
.B(n_325),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_321),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_326),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_325),
.Y(n_330)
);


endmodule