module fake_jpeg_26539_n_31 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_31);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_31;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_29;
wire n_15;

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_3),
.A2(n_9),
.B1(n_4),
.B2(n_0),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_SL g18 ( 
.A(n_14),
.B(n_1),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_16),
.C(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_1),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_8),
.B1(n_11),
.B2(n_5),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_22),
.B1(n_15),
.B2(n_16),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_17),
.B(n_2),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_15),
.A2(n_6),
.B1(n_10),
.B2(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_18),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_24),
.B(n_26),
.Y(n_29)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_25),
.B(n_27),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_21),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_23),
.B1(n_16),
.B2(n_26),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_29),
.Y(n_31)
);


endmodule