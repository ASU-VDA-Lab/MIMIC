module fake_netlist_1_6154_n_47 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_47);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_47;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_46;
wire n_30;
wire n_16;
wire n_26;
wire n_33;
wire n_25;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
INVx2_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_7), .Y(n_17) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_7), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_2), .Y(n_19) );
OAI22xp5_ASAP7_75t_SL g20 ( .A1(n_14), .A2(n_10), .B1(n_5), .B2(n_9), .Y(n_20) );
OA21x2_ASAP7_75t_L g21 ( .A1(n_3), .A2(n_13), .B(n_5), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_4), .B(n_9), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_2), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_18), .B(n_0), .Y(n_24) );
OAI22xp5_ASAP7_75t_L g25 ( .A1(n_20), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_25) );
AND2x4_ASAP7_75t_L g26 ( .A(n_16), .B(n_1), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_16), .Y(n_27) );
OAI21x1_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_16), .B(n_21), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_26), .B(n_23), .Y(n_29) );
A2O1A1Ixp33_ASAP7_75t_L g30 ( .A1(n_26), .A2(n_19), .B(n_17), .C(n_23), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_29), .B(n_24), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_28), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_31), .B(n_29), .Y(n_33) );
NAND2xp33_ASAP7_75t_SL g34 ( .A(n_32), .B(n_20), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
A2O1A1Ixp33_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_30), .B(n_28), .C(n_32), .Y(n_36) );
NAND2xp33_ASAP7_75t_R g37 ( .A(n_33), .B(n_21), .Y(n_37) );
AOI322xp5_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_19), .A3(n_17), .B1(n_25), .B2(n_22), .C1(n_8), .C2(n_10), .Y(n_38) );
A2O1A1Ixp33_ASAP7_75t_L g39 ( .A1(n_36), .A2(n_28), .B(n_25), .C(n_21), .Y(n_39) );
A2O1A1Ixp33_ASAP7_75t_L g40 ( .A1(n_35), .A2(n_21), .B(n_6), .C(n_4), .Y(n_40) );
OAI221xp5_ASAP7_75t_L g41 ( .A1(n_38), .A2(n_37), .B1(n_6), .B2(n_12), .C(n_15), .Y(n_41) );
NAND2x1p5_ASAP7_75t_L g42 ( .A(n_40), .B(n_11), .Y(n_42) );
INVx1_ASAP7_75t_L g43 ( .A(n_39), .Y(n_43) );
INVx1_ASAP7_75t_L g44 ( .A(n_43), .Y(n_44) );
INVx1_ASAP7_75t_L g45 ( .A(n_42), .Y(n_45) );
INVx1_ASAP7_75t_L g46 ( .A(n_44), .Y(n_46) );
AO221x1_ASAP7_75t_L g47 ( .A1(n_46), .A2(n_45), .B1(n_44), .B2(n_42), .C(n_41), .Y(n_47) );
endmodule