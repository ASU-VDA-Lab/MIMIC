module fake_jpeg_6738_n_191 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_191);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_9),
.B(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_36),
.Y(n_60)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_38),
.Y(n_71)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_2),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_3),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_4),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_28),
.Y(n_57)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_31),
.B1(n_29),
.B2(n_28),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_51),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_33),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_30),
.C(n_22),
.Y(n_93)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_29),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_23),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_74),
.B(n_80),
.C(n_22),
.Y(n_95)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_67),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_14),
.B1(n_26),
.B2(n_24),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_61),
.A2(n_75),
.B1(n_77),
.B2(n_36),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_31),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_23),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_50),
.B1(n_39),
.B2(n_24),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_79),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_70),
.B(n_78),
.Y(n_86)
);

AO22x1_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_15),
.B1(n_19),
.B2(n_26),
.Y(n_74)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_23),
.B1(n_18),
.B2(n_22),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_15),
.B1(n_14),
.B2(n_19),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_33),
.B(n_30),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_101),
.Y(n_107)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_16),
.Y(n_88)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_97),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_80),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_22),
.Y(n_94)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_104),
.B(n_78),
.C(n_64),
.Y(n_125)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_70),
.Y(n_123)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_18),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_100),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_18),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_4),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_103),
.B(n_105),
.Y(n_115)
);

BUFx24_ASAP7_75t_SL g105 ( 
.A(n_65),
.Y(n_105)
);

OA21x2_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_75),
.B(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_119),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_75),
.B1(n_58),
.B2(n_74),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_118),
.B1(n_126),
.B2(n_102),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_116),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_60),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_81),
.C(n_69),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_90),
.C(n_102),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_53),
.B1(n_61),
.B2(n_68),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_88),
.B(n_64),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_123),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_23),
.Y(n_124)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_124),
.B(n_103),
.CI(n_86),
.CON(n_137),
.SN(n_137)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_127),
.B1(n_92),
.B2(n_84),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_100),
.B1(n_94),
.B2(n_97),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_85),
.A2(n_53),
.B1(n_79),
.B2(n_47),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_130),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_106),
.B(n_92),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_139),
.B(n_121),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_114),
.B(n_82),
.Y(n_130)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_89),
.B1(n_84),
.B2(n_86),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_135),
.A2(n_136),
.B1(n_5),
.B2(n_6),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_140),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_72),
.C(n_6),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_114),
.A2(n_90),
.B(n_47),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_99),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_142),
.Y(n_146)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

AO221x1_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_120),
.B1(n_126),
.B2(n_107),
.C(n_125),
.Y(n_150)
);

XOR2x2_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_116),
.Y(n_144)
);

A2O1A1O1Ixp25_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_110),
.B(n_118),
.C(n_120),
.D(n_115),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_91),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_145),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_149),
.B1(n_133),
.B2(n_128),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_121),
.B(n_109),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_157),
.Y(n_163)
);

A2O1A1O1Ixp25_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_144),
.B(n_137),
.C(n_132),
.D(n_135),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_138),
.C(n_141),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_156),
.B(n_137),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_130),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_136),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_158),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_161),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_143),
.C(n_132),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_165),
.C(n_167),
.Y(n_175)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_140),
.C(n_129),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_168),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_153),
.C(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_134),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_157),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_173),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_153),
.B(n_149),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_179),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_146),
.C(n_154),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_173),
.C(n_172),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_168),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_169),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_155),
.C(n_11),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_5),
.B(n_6),
.Y(n_181)
);

AOI21x1_ASAP7_75t_L g184 ( 
.A1(n_181),
.A2(n_8),
.B(n_9),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_182),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_SL g188 ( 
.A1(n_183),
.A2(n_184),
.B(n_180),
.C(n_12),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_SL g187 ( 
.A(n_185),
.B(n_179),
.C(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_188),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_12),
.C(n_13),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_190),
.Y(n_191)
);


endmodule