module fake_jpeg_11564_n_202 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_202);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_42),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_25),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_9),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_5),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_78),
.B(n_0),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_31),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_1),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_54),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_1),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_77),
.B1(n_61),
.B2(n_79),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_104),
.B1(n_71),
.B2(n_68),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_61),
.B1(n_72),
.B2(n_67),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_59),
.B1(n_66),
.B2(n_57),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_105),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_64),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_79),
.B1(n_67),
.B2(n_72),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

BUFx16f_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_104),
.A2(n_73),
.B1(n_58),
.B2(n_87),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_5),
.C(n_7),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_113),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_58),
.B1(n_76),
.B2(n_84),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_111),
.B1(n_120),
.B2(n_123),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_76),
.B1(n_59),
.B2(n_63),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_111),
.B1(n_107),
.B2(n_116),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_87),
.B1(n_66),
.B2(n_74),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_126),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_62),
.B1(n_56),
.B2(n_60),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_124),
.A2(n_125),
.B1(n_2),
.B2(n_3),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_56),
.B1(n_3),
.B2(n_4),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_91),
.B(n_2),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_106),
.B1(n_60),
.B2(n_4),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_141),
.B1(n_36),
.B2(n_39),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_133),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_121),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_121),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_136),
.Y(n_157)
);

HAxp5_ASAP7_75t_SL g135 ( 
.A(n_124),
.B(n_106),
.CON(n_135),
.SN(n_135)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_144),
.B(n_14),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_142),
.A2(n_12),
.B(n_13),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_115),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_10),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_145),
.B(n_146),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_11),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_12),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_148),
.B(n_149),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_37),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_156),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_38),
.B1(n_17),
.B2(n_20),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_151),
.A2(n_154),
.B(n_155),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_141),
.A2(n_23),
.B1(n_28),
.B2(n_30),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_159),
.Y(n_180)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_32),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_142),
.C(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_33),
.B(n_34),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_144),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_35),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_166),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_167),
.A2(n_137),
.B1(n_44),
.B2(n_46),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_170),
.B(n_178),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_173),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_135),
.C(n_138),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_41),
.C(n_47),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_177),
.A2(n_151),
.B1(n_155),
.B2(n_165),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_157),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_168),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_181),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_160),
.B(n_154),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_186),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_189),
.B1(n_169),
.B2(n_179),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_163),
.B(n_153),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_187),
.B(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_172),
.B1(n_180),
.B2(n_174),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_192),
.C(n_193),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_187),
.C(n_190),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g197 ( 
.A(n_196),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_183),
.B(n_188),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_186),
.B1(n_193),
.B2(n_170),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_199),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_177),
.B(n_50),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_49),
.Y(n_202)
);


endmodule