module fake_ibex_839_n_1325 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_247, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_267, n_268, n_8, n_118, n_224, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_264, n_124, n_37, n_256, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_263, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_262, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_14, n_0, n_239, n_94, n_134, n_12, n_266, n_42, n_77, n_112, n_257, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_258, n_80, n_172, n_215, n_250, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_261, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_260, n_99, n_269, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_270, n_230, n_96, n_185, n_271, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_265, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_259, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1325);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_247;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_267;
input n_268;
input n_8;
input n_118;
input n_224;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_264;
input n_124;
input n_37;
input n_256;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_263;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_262;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_266;
input n_42;
input n_77;
input n_112;
input n_257;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_258;
input n_80;
input n_172;
input n_215;
input n_250;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_261;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_260;
input n_99;
input n_269;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_270;
input n_230;
input n_96;
input n_185;
input n_271;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_265;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_259;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1325;

wire n_1084;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_280;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_875;
wire n_1307;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1133;
wire n_904;
wire n_355;
wire n_646;
wire n_448;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_573;
wire n_359;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_397;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_451;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1108;
wire n_382;
wire n_1239;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_1281;
wire n_695;
wire n_639;
wire n_482;
wire n_282;
wire n_870;
wire n_1298;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_657;
wire n_1156;
wire n_1293;
wire n_749;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1015;
wire n_663;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_840;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_483;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_413;
wire n_1069;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_998;
wire n_1115;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_291;
wire n_318;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_997;
wire n_891;
wire n_303;
wire n_717;
wire n_668;
wire n_871;
wire n_485;
wire n_1315;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1265;
wire n_1048;
wire n_774;
wire n_588;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_423;
wire n_357;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_377;
wire n_647;
wire n_1291;
wire n_317;
wire n_326;
wire n_276;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_1112;
wire n_1267;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1021;
wire n_746;
wire n_1188;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_804;
wire n_484;
wire n_480;
wire n_1057;
wire n_354;
wire n_516;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_277;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1139;
wire n_858;
wire n_1018;
wire n_385;
wire n_1324;
wire n_782;
wire n_616;
wire n_833;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1221;
wire n_284;
wire n_1047;
wire n_792;
wire n_1314;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_478;
wire n_336;
wire n_861;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1098;
wire n_584;
wire n_1187;
wire n_698;
wire n_1061;
wire n_682;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1023;
wire n_568;
wire n_813;
wire n_1211;
wire n_1284;
wire n_1116;
wire n_791;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1074;
wire n_759;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_735;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1033;
wire n_627;
wire n_990;
wire n_322;
wire n_888;
wire n_582;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1002;
wire n_1111;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1145;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1277;
wire n_1016;
wire n_680;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_908;
wire n_565;
wire n_1123;
wire n_1272;
wire n_984;
wire n_394;
wire n_364;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g272 ( 
.A(n_111),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_147),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_104),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_35),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_260),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_26),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_112),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_234),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_139),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_74),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_165),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_34),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_70),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_144),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_156),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_58),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_235),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_149),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_146),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_127),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_123),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_194),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_126),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_261),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_6),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_253),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_63),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_201),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_266),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_202),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_182),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_47),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_229),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_189),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_6),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_263),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_270),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_238),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_122),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_58),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_248),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_239),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_129),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_161),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_153),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_19),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_173),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_50),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_219),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_255),
.Y(n_323)
);

BUFx5_ASAP7_75t_L g324 ( 
.A(n_116),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_157),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_226),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_181),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_128),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_190),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_9),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_177),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_140),
.Y(n_332)
);

BUFx2_ASAP7_75t_SL g333 ( 
.A(n_163),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_64),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_45),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_204),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_180),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_99),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_271),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_251),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_228),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_246),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_167),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_155),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_78),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_64),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_48),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_88),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_240),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_215),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_231),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_178),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_162),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_109),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_233),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_32),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_230),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_227),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_203),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_158),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_259),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_174),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_262),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_1),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_138),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_101),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_225),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_197),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_159),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_218),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_172),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_142),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_74),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_120),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_252),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_232),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_199),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_223),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_151),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_207),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_49),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_96),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_98),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_130),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_88),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_195),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_224),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_60),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_209),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_51),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_84),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_171),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_170),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_62),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_264),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_210),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_212),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_241),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_43),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_66),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_52),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_17),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_244),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_243),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_257),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_61),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_83),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_57),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_216),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_131),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_198),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_206),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_93),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_184),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_60),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_89),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_50),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_245),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_72),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_117),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_249),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_179),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_136),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_92),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_73),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_12),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_51),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_39),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_34),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_46),
.Y(n_430)
);

BUFx10_ASAP7_75t_L g431 ( 
.A(n_72),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_9),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_102),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_62),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_28),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_135),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_269),
.Y(n_437)
);

BUFx10_ASAP7_75t_L g438 ( 
.A(n_237),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_164),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_247),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_84),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_250),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_141),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_103),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_97),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_20),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_30),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_236),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_56),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_196),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_258),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_191),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_33),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_40),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_211),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_267),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_55),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_242),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_14),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_213),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_12),
.Y(n_461)
);

INVx4_ASAP7_75t_R g462 ( 
.A(n_18),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_424),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_335),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_335),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_454),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_454),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_324),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_276),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_407),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_L g471 ( 
.A(n_356),
.B(n_0),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_315),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_461),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_277),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_284),
.B(n_0),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_419),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_308),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_349),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_354),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_427),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_440),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_324),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_345),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_324),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_431),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_282),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_331),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_L g488 ( 
.A(n_373),
.B(n_1),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_381),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_282),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_L g491 ( 
.A(n_385),
.B(n_2),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_394),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_279),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_332),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_283),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_431),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_285),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_431),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_286),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_400),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_402),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_406),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_417),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_289),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_298),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_300),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_324),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_313),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_319),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_311),
.B(n_2),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_425),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_321),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_426),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_R g514 ( 
.A(n_273),
.B(n_90),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_434),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_330),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_334),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_346),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_347),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_348),
.Y(n_520)
);

CKINVDCx14_ASAP7_75t_R g521 ( 
.A(n_297),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_446),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_453),
.B(n_459),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_364),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_390),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_297),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_297),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_438),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_391),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_272),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_509),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_468),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_476),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_530),
.B(n_287),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_526),
.B(n_388),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_465),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_474),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_477),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_483),
.B(n_489),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_482),
.B(n_287),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_492),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_482),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_484),
.B(n_507),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_480),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_500),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_484),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_507),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_521),
.B(n_399),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_521),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_501),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_502),
.B(n_290),
.Y(n_551)
);

AND2x6_ASAP7_75t_L g552 ( 
.A(n_527),
.B(n_326),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_466),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_503),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_475),
.B(n_290),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_511),
.B(n_293),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_528),
.B(n_293),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_493),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_513),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_467),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_504),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_522),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_473),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_512),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_463),
.B(n_294),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_518),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_523),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_471),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_488),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_491),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_518),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_495),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_510),
.B(n_296),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_470),
.B(n_388),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_515),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_485),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_514),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_497),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_505),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_SL g580 ( 
.A(n_496),
.B(n_401),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_472),
.B(n_326),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_506),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_516),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_519),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_525),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_529),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_487),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_472),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_496),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_490),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_498),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_498),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_499),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_499),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_508),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_508),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_517),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_517),
.Y(n_598)
);

NAND2xp33_ASAP7_75t_SL g599 ( 
.A(n_520),
.B(n_408),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_520),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_524),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_469),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_524),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_478),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_479),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_481),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_486),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_486),
.B(n_415),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_494),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_464),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_464),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_R g612 ( 
.A(n_472),
.B(n_416),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_464),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_468),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_464),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_464),
.Y(n_616)
);

OA21x2_ASAP7_75t_L g617 ( 
.A1(n_468),
.A2(n_339),
.B(n_299),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_464),
.Y(n_618)
);

NAND2xp33_ASAP7_75t_SL g619 ( 
.A(n_496),
.B(n_388),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_476),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_464),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_464),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_464),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_468),
.B(n_299),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_464),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_521),
.B(n_428),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_526),
.B(n_327),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_526),
.B(n_327),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_468),
.Y(n_629)
);

AND2x6_ASAP7_75t_L g630 ( 
.A(n_526),
.B(n_338),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_468),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_464),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_464),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_509),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_476),
.Y(n_635)
);

OA21x2_ASAP7_75t_L g636 ( 
.A1(n_468),
.A2(n_344),
.B(n_339),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_464),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_509),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_468),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_464),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_468),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_468),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_530),
.B(n_344),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_476),
.Y(n_644)
);

NAND2x1_ASAP7_75t_L g645 ( 
.A(n_526),
.B(n_462),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_468),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_470),
.A2(n_430),
.B1(n_432),
.B2(n_429),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_464),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_464),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_526),
.B(n_338),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_634),
.B(n_564),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_SL g652 ( 
.A(n_549),
.B(n_435),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_567),
.B(n_305),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_553),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_553),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_553),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_567),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_L g658 ( 
.A(n_552),
.B(n_324),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_576),
.B(n_396),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_634),
.B(n_441),
.Y(n_660)
);

AND2x6_ASAP7_75t_L g661 ( 
.A(n_572),
.B(n_362),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_564),
.B(n_447),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_612),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_575),
.B(n_537),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_578),
.B(n_449),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_535),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_574),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_549),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_638),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_635),
.B(n_457),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_577),
.B(n_274),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_572),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_561),
.A2(n_288),
.B1(n_291),
.B2(n_275),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_R g674 ( 
.A(n_580),
.B(n_278),
.Y(n_674)
);

INVx6_ASAP7_75t_L g675 ( 
.A(n_587),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_533),
.B(n_544),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_583),
.B(n_362),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_584),
.B(n_375),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_536),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_610),
.Y(n_680)
);

INVx4_ASAP7_75t_SL g681 ( 
.A(n_581),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_548),
.B(n_280),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_626),
.B(n_281),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_611),
.Y(n_684)
);

XOR2x2_ASAP7_75t_L g685 ( 
.A(n_593),
.B(n_596),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_560),
.Y(n_686)
);

INVxp33_ASAP7_75t_L g687 ( 
.A(n_544),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_617),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_538),
.A2(n_333),
.B1(n_306),
.B2(n_307),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_620),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_620),
.Y(n_691)
);

INVx6_ASAP7_75t_L g692 ( 
.A(n_587),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_563),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_582),
.B(n_375),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_613),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_563),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_644),
.B(n_3),
.Y(n_697)
);

AND2x6_ASAP7_75t_L g698 ( 
.A(n_582),
.B(n_420),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_579),
.B(n_420),
.Y(n_699)
);

AND2x2_ASAP7_75t_SL g700 ( 
.A(n_566),
.B(n_303),
.Y(n_700)
);

BUFx10_ASAP7_75t_L g701 ( 
.A(n_587),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_615),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_588),
.B(n_292),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_644),
.Y(n_704)
);

AND2x6_ASAP7_75t_L g705 ( 
.A(n_585),
.B(n_312),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_568),
.B(n_295),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_616),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_627),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_628),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_618),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_546),
.Y(n_711)
);

INVx5_ASAP7_75t_L g712 ( 
.A(n_546),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_621),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_645),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_622),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_586),
.B(n_316),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_558),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_541),
.A2(n_545),
.B1(n_554),
.B2(n_550),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_623),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_650),
.B(n_558),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_631),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_559),
.B(n_302),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_625),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_617),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_636),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_589),
.B(n_3),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_581),
.Y(n_727)
);

OR2x6_ASAP7_75t_L g728 ( 
.A(n_590),
.B(n_317),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_562),
.B(n_304),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_636),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_649),
.Y(n_731)
);

CKINVDCx11_ASAP7_75t_R g732 ( 
.A(n_594),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_566),
.B(n_309),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_631),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_586),
.B(n_310),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_632),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_573),
.B(n_314),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_633),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_591),
.B(n_4),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_552),
.A2(n_322),
.B1(n_328),
.B2(n_318),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_639),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_573),
.B(n_565),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_593),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_639),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_637),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_646),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_552),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_640),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_539),
.B(n_320),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_648),
.Y(n_750)
);

NOR3xp33_ASAP7_75t_SL g751 ( 
.A(n_599),
.B(n_325),
.C(n_323),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_571),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_539),
.Y(n_753)
);

NOR2x1p5_ASAP7_75t_L g754 ( 
.A(n_602),
.B(n_337),
.Y(n_754)
);

OR2x6_ASAP7_75t_L g755 ( 
.A(n_590),
.B(n_329),
.Y(n_755)
);

AND2x6_ASAP7_75t_L g756 ( 
.A(n_606),
.B(n_336),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_630),
.Y(n_757)
);

OAI22x1_ASAP7_75t_L g758 ( 
.A1(n_595),
.A2(n_597),
.B1(n_601),
.B2(n_600),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_532),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_555),
.B(n_557),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_581),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_569),
.B(n_341),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_647),
.B(n_340),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_581),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_608),
.B(n_4),
.Y(n_765)
);

INVxp67_ASAP7_75t_SL g766 ( 
.A(n_534),
.Y(n_766)
);

NAND3xp33_ASAP7_75t_L g767 ( 
.A(n_619),
.B(n_351),
.C(n_350),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_630),
.A2(n_359),
.B1(n_365),
.B2(n_355),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_551),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_556),
.Y(n_770)
);

XNOR2xp5_ASAP7_75t_L g771 ( 
.A(n_607),
.B(n_5),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_602),
.Y(n_772)
);

BUFx10_ASAP7_75t_L g773 ( 
.A(n_604),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_555),
.B(n_342),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_643),
.Y(n_775)
);

AND2x6_ASAP7_75t_L g776 ( 
.A(n_605),
.B(n_370),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_592),
.B(n_5),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_570),
.B(n_374),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_630),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_598),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_630),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_557),
.B(n_343),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_603),
.B(n_352),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_609),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_630),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_542),
.A2(n_376),
.B1(n_387),
.B2(n_379),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_619),
.A2(n_393),
.B1(n_410),
.B2(n_392),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_547),
.B(n_353),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_540),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_614),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_629),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_624),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_624),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_641),
.B(n_358),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_642),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_543),
.B(n_360),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_553),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_567),
.B(n_414),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_575),
.B(n_361),
.Y(n_799)
);

INVx4_ASAP7_75t_SL g800 ( 
.A(n_581),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_553),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_553),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_553),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_553),
.Y(n_804)
);

BUFx10_ASAP7_75t_L g805 ( 
.A(n_549),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_553),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_567),
.B(n_363),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_634),
.B(n_7),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_567),
.B(n_422),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_531),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_567),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_553),
.Y(n_812)
);

INVx4_ASAP7_75t_L g813 ( 
.A(n_567),
.Y(n_813)
);

OAI221xp5_ASAP7_75t_L g814 ( 
.A1(n_717),
.A2(n_690),
.B1(n_720),
.B2(n_753),
.C(n_752),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_766),
.Y(n_815)
);

NAND2x1p5_ASAP7_75t_L g816 ( 
.A(n_651),
.B(n_423),
.Y(n_816)
);

AO22x2_ASAP7_75t_L g817 ( 
.A1(n_697),
.A2(n_436),
.B1(n_437),
.B2(n_433),
.Y(n_817)
);

AO22x2_ASAP7_75t_L g818 ( 
.A1(n_808),
.A2(n_456),
.B1(n_439),
.B2(n_384),
.Y(n_818)
);

AO22x2_ASAP7_75t_L g819 ( 
.A1(n_765),
.A2(n_384),
.B1(n_418),
.B2(n_357),
.Y(n_819)
);

XNOR2xp5_ASAP7_75t_L g820 ( 
.A(n_685),
.B(n_8),
.Y(n_820)
);

AO22x2_ASAP7_75t_L g821 ( 
.A1(n_662),
.A2(n_676),
.B1(n_813),
.B2(n_716),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_SL g822 ( 
.A1(n_691),
.A2(n_367),
.B1(n_368),
.B2(n_366),
.Y(n_822)
);

AO22x2_ASAP7_75t_L g823 ( 
.A1(n_716),
.A2(n_418),
.B1(n_455),
.B2(n_357),
.Y(n_823)
);

NOR2x1p5_ASAP7_75t_L g824 ( 
.A(n_704),
.B(n_369),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_769),
.Y(n_825)
);

OAI221xp5_ASAP7_75t_L g826 ( 
.A1(n_670),
.A2(n_460),
.B1(n_455),
.B2(n_371),
.C(n_372),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_770),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_669),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_805),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_700),
.A2(n_378),
.B1(n_380),
.B2(n_377),
.Y(n_830)
);

INVx1_ASAP7_75t_SL g831 ( 
.A(n_810),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_775),
.Y(n_832)
);

XNOR2xp5_ASAP7_75t_L g833 ( 
.A(n_663),
.B(n_8),
.Y(n_833)
);

AO22x2_ASAP7_75t_L g834 ( 
.A1(n_726),
.A2(n_460),
.B1(n_13),
.B2(n_10),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_668),
.B(n_11),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_687),
.B(n_382),
.Y(n_836)
);

AO22x2_ASAP7_75t_L g837 ( 
.A1(n_739),
.A2(n_15),
.B1(n_11),
.B2(n_13),
.Y(n_837)
);

AO22x2_ASAP7_75t_L g838 ( 
.A1(n_653),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_660),
.A2(n_386),
.B1(n_389),
.B2(n_383),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_743),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_653),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_657),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_811),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_805),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_798),
.B(n_395),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_667),
.Y(n_846)
);

OAI221xp5_ASAP7_75t_L g847 ( 
.A1(n_664),
.A2(n_397),
.B1(n_404),
.B2(n_403),
.C(n_398),
.Y(n_847)
);

AO22x2_ASAP7_75t_L g848 ( 
.A1(n_777),
.A2(n_19),
.B1(n_16),
.B2(n_18),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_668),
.B(n_20),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_679),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_733),
.B(n_21),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_680),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_665),
.B(n_405),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_672),
.B(n_728),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_684),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_672),
.B(n_21),
.Y(n_856)
);

AO22x2_ASAP7_75t_L g857 ( 
.A1(n_809),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_701),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_755),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_695),
.Y(n_860)
);

AO22x2_ASAP7_75t_L g861 ( 
.A1(n_809),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_702),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_707),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_718),
.A2(n_458),
.B1(n_411),
.B2(n_412),
.Y(n_864)
);

AO22x2_ASAP7_75t_L g865 ( 
.A1(n_665),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_742),
.B(n_409),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_754),
.B(n_27),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_710),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_713),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_715),
.Y(n_870)
);

AO22x2_ASAP7_75t_L g871 ( 
.A1(n_694),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_871)
);

AO22x2_ASAP7_75t_L g872 ( 
.A1(n_694),
.A2(n_33),
.B1(n_29),
.B2(n_31),
.Y(n_872)
);

OR2x2_ASAP7_75t_SL g873 ( 
.A(n_771),
.B(n_301),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_719),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_723),
.Y(n_875)
);

NAND2x1p5_ASAP7_75t_L g876 ( 
.A(n_708),
.B(n_709),
.Y(n_876)
);

AO22x2_ASAP7_75t_L g877 ( 
.A1(n_673),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_877)
);

AO22x2_ASAP7_75t_L g878 ( 
.A1(n_762),
.A2(n_41),
.B1(n_36),
.B2(n_38),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_701),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_795),
.Y(n_880)
);

AO22x2_ASAP7_75t_L g881 ( 
.A1(n_762),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_755),
.B(n_42),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_736),
.Y(n_883)
);

OAI221xp5_ASAP7_75t_L g884 ( 
.A1(n_689),
.A2(n_452),
.B1(n_413),
.B2(n_450),
.C(n_448),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_763),
.B(n_421),
.Y(n_885)
);

INVxp67_ASAP7_75t_L g886 ( 
.A(n_807),
.Y(n_886)
);

AO22x2_ASAP7_75t_L g887 ( 
.A1(n_778),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_887)
);

OAI221xp5_ASAP7_75t_L g888 ( 
.A1(n_786),
.A2(n_442),
.B1(n_445),
.B2(n_444),
.C(n_443),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_772),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_745),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_783),
.B(n_47),
.Y(n_891)
);

AO22x2_ASAP7_75t_L g892 ( 
.A1(n_778),
.A2(n_53),
.B1(n_49),
.B2(n_52),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_791),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_748),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_791),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_674),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_731),
.B(n_738),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_780),
.B(n_54),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_732),
.Y(n_899)
);

AO22x2_ASAP7_75t_L g900 ( 
.A1(n_677),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_750),
.Y(n_901)
);

AO22x2_ASAP7_75t_L g902 ( 
.A1(n_677),
.A2(n_63),
.B1(n_59),
.B2(n_61),
.Y(n_902)
);

AO22x2_ASAP7_75t_L g903 ( 
.A1(n_678),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_659),
.B(n_65),
.Y(n_904)
);

NAND3xp33_ASAP7_75t_L g905 ( 
.A(n_784),
.B(n_451),
.C(n_67),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_666),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_705),
.B(n_68),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_760),
.Y(n_908)
);

OR2x6_ASAP7_75t_L g909 ( 
.A(n_675),
.B(n_451),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_678),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_699),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_699),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_771),
.B(n_68),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_789),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_792),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_793),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_773),
.B(n_69),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_693),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_759),
.Y(n_919)
);

OAI221xp5_ASAP7_75t_L g920 ( 
.A1(n_652),
.A2(n_71),
.B1(n_73),
.B2(n_75),
.C(n_76),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_758),
.B(n_76),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_776),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_756),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_714),
.B(n_77),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_790),
.Y(n_925)
);

AO22x2_ASAP7_75t_L g926 ( 
.A1(n_767),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_926)
);

OAI221xp5_ASAP7_75t_L g927 ( 
.A1(n_751),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.C(n_83),
.Y(n_927)
);

AO22x2_ASAP7_75t_L g928 ( 
.A1(n_681),
.A2(n_82),
.B1(n_85),
.B2(n_86),
.Y(n_928)
);

BUFx8_ASAP7_75t_L g929 ( 
.A(n_661),
.Y(n_929)
);

NAND2x1p5_ASAP7_75t_L g930 ( 
.A(n_747),
.B(n_85),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_692),
.Y(n_931)
);

BUFx6f_ASAP7_75t_SL g932 ( 
.A(n_773),
.Y(n_932)
);

CKINVDCx16_ASAP7_75t_R g933 ( 
.A(n_661),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_692),
.Y(n_934)
);

NOR2xp67_ASAP7_75t_L g935 ( 
.A(n_787),
.B(n_86),
.Y(n_935)
);

AO22x2_ASAP7_75t_L g936 ( 
.A1(n_681),
.A2(n_800),
.B1(n_757),
.B2(n_776),
.Y(n_936)
);

AO22x2_ASAP7_75t_L g937 ( 
.A1(n_800),
.A2(n_757),
.B1(n_776),
.B2(n_698),
.Y(n_937)
);

NOR2xp67_ASAP7_75t_L g938 ( 
.A(n_735),
.B(n_706),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_844),
.B(n_829),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_844),
.B(n_779),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_879),
.B(n_779),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_859),
.B(n_785),
.Y(n_942)
);

NAND2xp33_ASAP7_75t_SL g943 ( 
.A(n_932),
.B(n_785),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_825),
.B(n_827),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_815),
.B(n_727),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_840),
.B(n_933),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_835),
.B(n_761),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_832),
.B(n_737),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_849),
.B(n_764),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_822),
.B(n_781),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_816),
.B(n_740),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_886),
.B(n_768),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_831),
.B(n_712),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_897),
.B(n_712),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_856),
.B(n_712),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_841),
.B(n_703),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_839),
.B(n_836),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_917),
.B(n_794),
.Y(n_958)
);

NAND2xp33_ASAP7_75t_SL g959 ( 
.A(n_896),
.B(n_688),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_898),
.B(n_796),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_858),
.B(n_688),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_830),
.B(n_682),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_929),
.B(n_683),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_864),
.B(n_853),
.Y(n_964)
);

NAND2xp33_ASAP7_75t_SL g965 ( 
.A(n_889),
.B(n_724),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_850),
.B(n_698),
.Y(n_966)
);

NAND2xp33_ASAP7_75t_SL g967 ( 
.A(n_824),
.B(n_725),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_828),
.B(n_845),
.Y(n_968)
);

NAND2xp33_ASAP7_75t_SL g969 ( 
.A(n_937),
.B(n_730),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_852),
.B(n_749),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_821),
.B(n_799),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_855),
.B(n_774),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_860),
.B(n_782),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_867),
.B(n_801),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_851),
.B(n_801),
.Y(n_975)
);

NAND2xp33_ASAP7_75t_SL g976 ( 
.A(n_937),
.B(n_722),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_923),
.B(n_804),
.Y(n_977)
);

NAND2xp33_ASAP7_75t_SL g978 ( 
.A(n_934),
.B(n_729),
.Y(n_978)
);

NAND2xp33_ASAP7_75t_SL g979 ( 
.A(n_936),
.B(n_812),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_821),
.B(n_671),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_882),
.B(n_788),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_930),
.B(n_806),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_891),
.B(n_812),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_862),
.B(n_658),
.Y(n_984)
);

NAND2xp33_ASAP7_75t_SL g985 ( 
.A(n_936),
.B(n_734),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_854),
.B(n_817),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_938),
.B(n_734),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_863),
.B(n_654),
.Y(n_988)
);

NAND2xp33_ASAP7_75t_SL g989 ( 
.A(n_907),
.B(n_744),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_868),
.B(n_869),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_935),
.B(n_744),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_870),
.B(n_655),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_924),
.B(n_744),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_904),
.B(n_746),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_874),
.B(n_746),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_875),
.B(n_656),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_883),
.B(n_686),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_890),
.B(n_696),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_894),
.B(n_797),
.Y(n_999)
);

NAND2xp33_ASAP7_75t_SL g1000 ( 
.A(n_901),
.B(n_921),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_911),
.B(n_802),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_912),
.B(n_803),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_893),
.B(n_711),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_823),
.B(n_721),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_895),
.B(n_741),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_823),
.B(n_87),
.Y(n_1006)
);

NAND2xp33_ASAP7_75t_SL g1007 ( 
.A(n_913),
.B(n_89),
.Y(n_1007)
);

NAND2xp33_ASAP7_75t_SL g1008 ( 
.A(n_919),
.B(n_91),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_854),
.B(n_94),
.Y(n_1009)
);

NAND2xp33_ASAP7_75t_SL g1010 ( 
.A(n_925),
.B(n_95),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_876),
.B(n_100),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_906),
.B(n_105),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_931),
.B(n_106),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_910),
.B(n_107),
.Y(n_1014)
);

NAND2xp33_ASAP7_75t_SL g1015 ( 
.A(n_866),
.B(n_108),
.Y(n_1015)
);

NAND2xp33_ASAP7_75t_SL g1016 ( 
.A(n_899),
.B(n_110),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_818),
.B(n_113),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_908),
.B(n_114),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_905),
.B(n_115),
.Y(n_1019)
);

NAND2xp33_ASAP7_75t_SL g1020 ( 
.A(n_820),
.B(n_118),
.Y(n_1020)
);

NAND2xp33_ASAP7_75t_SL g1021 ( 
.A(n_842),
.B(n_119),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_885),
.B(n_121),
.Y(n_1022)
);

NAND2xp33_ASAP7_75t_SL g1023 ( 
.A(n_843),
.B(n_124),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_922),
.B(n_125),
.Y(n_1024)
);

NAND2xp33_ASAP7_75t_SL g1025 ( 
.A(n_833),
.B(n_132),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_880),
.B(n_133),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_819),
.B(n_134),
.Y(n_1027)
);

NAND2xp33_ASAP7_75t_SL g1028 ( 
.A(n_846),
.B(n_137),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_819),
.B(n_143),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_818),
.B(n_145),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_990),
.Y(n_1031)
);

AO31x2_ASAP7_75t_L g1032 ( 
.A1(n_1027),
.A2(n_916),
.A3(n_914),
.B(n_915),
.Y(n_1032)
);

CKINVDCx6p67_ASAP7_75t_R g1033 ( 
.A(n_1009),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_944),
.Y(n_1034)
);

OAI22x1_ASAP7_75t_L g1035 ( 
.A1(n_986),
.A2(n_865),
.B1(n_838),
.B2(n_861),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_1009),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_944),
.Y(n_1037)
);

AO22x2_ASAP7_75t_L g1038 ( 
.A1(n_1017),
.A2(n_865),
.B1(n_903),
.B2(n_900),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_1009),
.B(n_918),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_965),
.Y(n_1040)
);

NAND2xp33_ASAP7_75t_L g1041 ( 
.A(n_985),
.B(n_928),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_944),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_948),
.A2(n_814),
.B(n_826),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_1018),
.A2(n_909),
.B(n_927),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_960),
.B(n_873),
.Y(n_1045)
);

NOR2xp67_ASAP7_75t_L g1046 ( 
.A(n_963),
.B(n_920),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_1026),
.A2(n_926),
.B(n_834),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1007),
.A2(n_834),
.B1(n_837),
.B2(n_848),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_972),
.B(n_848),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_964),
.A2(n_847),
.B(n_888),
.C(n_884),
.Y(n_1050)
);

OAI22x1_ASAP7_75t_L g1051 ( 
.A1(n_1030),
.A2(n_838),
.B1(n_861),
.B2(n_857),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_956),
.B(n_837),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_979),
.Y(n_1053)
);

BUFx12f_ASAP7_75t_L g1054 ( 
.A(n_981),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_R g1055 ( 
.A(n_943),
.B(n_900),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_939),
.B(n_148),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_946),
.Y(n_1057)
);

BUFx24_ASAP7_75t_L g1058 ( 
.A(n_969),
.Y(n_1058)
);

NAND3xp33_ASAP7_75t_L g1059 ( 
.A(n_1000),
.B(n_903),
.C(n_902),
.Y(n_1059)
);

AO21x2_ASAP7_75t_L g1060 ( 
.A1(n_1004),
.A2(n_902),
.B(n_872),
.Y(n_1060)
);

AND2x6_ASAP7_75t_SL g1061 ( 
.A(n_1006),
.B(n_878),
.Y(n_1061)
);

CKINVDCx16_ASAP7_75t_R g1062 ( 
.A(n_1016),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_961),
.A2(n_872),
.B(n_871),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_995),
.A2(n_871),
.B(n_857),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_994),
.A2(n_881),
.B(n_878),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_970),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_988),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_973),
.A2(n_892),
.B(n_887),
.C(n_881),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_957),
.B(n_887),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_952),
.B(n_892),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_974),
.B(n_877),
.Y(n_1071)
);

INVx5_ASAP7_75t_L g1072 ( 
.A(n_971),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_962),
.B(n_980),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_951),
.B(n_877),
.Y(n_1074)
);

AO31x2_ASAP7_75t_L g1075 ( 
.A1(n_1029),
.A2(n_150),
.A3(n_152),
.B(n_154),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_958),
.B(n_160),
.Y(n_1076)
);

CKINVDCx11_ASAP7_75t_R g1077 ( 
.A(n_978),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_992),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_967),
.B(n_959),
.Y(n_1079)
);

AO31x2_ASAP7_75t_L g1080 ( 
.A1(n_984),
.A2(n_166),
.A3(n_168),
.B(n_169),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_941),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_947),
.B(n_949),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_968),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_993),
.Y(n_1084)
);

OA21x2_ASAP7_75t_L g1085 ( 
.A1(n_1019),
.A2(n_175),
.B(n_176),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_991),
.B(n_268),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_955),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_R g1088 ( 
.A(n_1025),
.B(n_1020),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_996),
.Y(n_1089)
);

NOR2xp67_ASAP7_75t_L g1090 ( 
.A(n_953),
.B(n_183),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_976),
.B(n_185),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_966),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_950),
.B(n_186),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_SL g1094 ( 
.A1(n_982),
.A2(n_187),
.B(n_188),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_1042),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1031),
.B(n_942),
.Y(n_1096)
);

CKINVDCx20_ASAP7_75t_R g1097 ( 
.A(n_1033),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_1052),
.B(n_954),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1071),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1068),
.B(n_1001),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1066),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_1055),
.B(n_1021),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1043),
.A2(n_1024),
.B(n_975),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1038),
.B(n_1035),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1078),
.Y(n_1105)
);

OAI21xp33_ASAP7_75t_SL g1106 ( 
.A1(n_1039),
.A2(n_983),
.B(n_1013),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_1042),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1038),
.Y(n_1108)
);

NAND3xp33_ASAP7_75t_L g1109 ( 
.A(n_1059),
.B(n_987),
.C(n_1022),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1067),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1036),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_1042),
.Y(n_1112)
);

NOR2x1_ASAP7_75t_SL g1113 ( 
.A(n_1058),
.B(n_1079),
.Y(n_1113)
);

AO21x2_ASAP7_75t_L g1114 ( 
.A1(n_1047),
.A2(n_1014),
.B(n_1012),
.Y(n_1114)
);

NOR2xp67_ASAP7_75t_L g1115 ( 
.A(n_1051),
.B(n_940),
.Y(n_1115)
);

AOI221xp5_ASAP7_75t_L g1116 ( 
.A1(n_1069),
.A2(n_1015),
.B1(n_1028),
.B2(n_1023),
.C(n_1002),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1067),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_1053),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1040),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1048),
.A2(n_1011),
.B1(n_945),
.B2(n_977),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_1077),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1044),
.A2(n_1008),
.B(n_1010),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_1062),
.B(n_989),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_1034),
.Y(n_1124)
);

OAI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_1049),
.A2(n_999),
.B1(n_998),
.B2(n_997),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_1054),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_1088),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_1070),
.B(n_1003),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1081),
.Y(n_1129)
);

OR2x2_ASAP7_75t_L g1130 ( 
.A(n_1074),
.B(n_1005),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1063),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1045),
.B(n_265),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1037),
.B(n_1072),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1110),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1131),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1110),
.Y(n_1136)
);

AOI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1102),
.A2(n_1091),
.B(n_1065),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_1108),
.B(n_1072),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1117),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1103),
.A2(n_1046),
.B(n_1064),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_1095),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1099),
.B(n_1060),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_1118),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1117),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_1133),
.B(n_1072),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1101),
.Y(n_1146)
);

AOI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1102),
.A2(n_1122),
.B(n_1115),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_1105),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1129),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1104),
.B(n_1061),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_1126),
.Y(n_1151)
);

INVxp67_ASAP7_75t_SL g1152 ( 
.A(n_1119),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_1129),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1129),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1129),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1119),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1130),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1128),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_1111),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_1133),
.Y(n_1160)
);

OR2x6_ASAP7_75t_L g1161 ( 
.A(n_1123),
.B(n_1041),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1124),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_1121),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1133),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1096),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1148),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_1143),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1138),
.B(n_1113),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1146),
.Y(n_1169)
);

BUFx24_ASAP7_75t_SL g1170 ( 
.A(n_1163),
.Y(n_1170)
);

BUFx24_ASAP7_75t_SL g1171 ( 
.A(n_1150),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1157),
.B(n_1098),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_1143),
.Y(n_1173)
);

INVx8_ASAP7_75t_L g1174 ( 
.A(n_1145),
.Y(n_1174)
);

INVxp67_ASAP7_75t_L g1175 ( 
.A(n_1159),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_1159),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1138),
.B(n_1095),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1157),
.B(n_1073),
.Y(n_1178)
);

XNOR2xp5_ASAP7_75t_L g1179 ( 
.A(n_1151),
.B(n_1121),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1158),
.B(n_1100),
.Y(n_1180)
);

INVxp67_ASAP7_75t_L g1181 ( 
.A(n_1152),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1146),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_R g1183 ( 
.A(n_1147),
.B(n_1097),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_R g1184 ( 
.A(n_1147),
.B(n_1097),
.Y(n_1184)
);

INVxp67_ASAP7_75t_L g1185 ( 
.A(n_1141),
.Y(n_1185)
);

CKINVDCx12_ASAP7_75t_R g1186 ( 
.A(n_1161),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1138),
.B(n_1112),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1158),
.B(n_1126),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1138),
.B(n_1112),
.Y(n_1189)
);

BUFx8_ASAP7_75t_SL g1190 ( 
.A(n_1161),
.Y(n_1190)
);

BUFx10_ASAP7_75t_L g1191 ( 
.A(n_1145),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1165),
.B(n_1125),
.Y(n_1192)
);

BUFx8_ASAP7_75t_SL g1193 ( 
.A(n_1161),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1161),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_1176),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1182),
.B(n_1169),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_1183),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1180),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1166),
.B(n_1142),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1173),
.B(n_1142),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1175),
.B(n_1156),
.Y(n_1201)
);

OR2x2_ASAP7_75t_L g1202 ( 
.A(n_1167),
.B(n_1172),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1181),
.B(n_1156),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1192),
.B(n_1135),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1185),
.Y(n_1205)
);

INVxp67_ASAP7_75t_SL g1206 ( 
.A(n_1190),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1184),
.B(n_1127),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1193),
.A2(n_1161),
.B1(n_1140),
.B2(n_1164),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_1191),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1178),
.Y(n_1210)
);

BUFx2_ASAP7_75t_SL g1211 ( 
.A(n_1191),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1177),
.B(n_1135),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_1188),
.B(n_1134),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1186),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1174),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1171),
.A2(n_1164),
.B1(n_1109),
.B2(n_1120),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1194),
.A2(n_1174),
.B1(n_1168),
.B2(n_1160),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1203),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1206),
.Y(n_1219)
);

NAND3xp33_ASAP7_75t_L g1220 ( 
.A(n_1205),
.B(n_1165),
.C(n_1179),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1203),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1196),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1215),
.A2(n_1168),
.B1(n_1174),
.B2(n_1127),
.Y(n_1223)
);

AOI222xp33_ASAP7_75t_L g1224 ( 
.A1(n_1206),
.A2(n_1083),
.B1(n_1170),
.B2(n_1087),
.C1(n_1057),
.C2(n_1125),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1210),
.B(n_1198),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1195),
.B(n_1177),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1196),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1201),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1201),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1204),
.B(n_1187),
.Y(n_1230)
);

OA332x1_ASAP7_75t_L g1231 ( 
.A1(n_1202),
.A2(n_1137),
.A3(n_1189),
.B1(n_1187),
.B2(n_1160),
.B3(n_1123),
.C1(n_1162),
.C2(n_1141),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1218),
.B(n_1197),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1221),
.B(n_1198),
.Y(n_1233)
);

OR2x6_ASAP7_75t_SL g1234 ( 
.A(n_1220),
.B(n_1202),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1222),
.B(n_1200),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1228),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1229),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1225),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_1222),
.B(n_1199),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1227),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1219),
.B(n_1197),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1230),
.B(n_1212),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1226),
.B(n_1230),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1227),
.B(n_1195),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1224),
.B(n_1200),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1223),
.B(n_1199),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1234),
.A2(n_1215),
.B1(n_1209),
.B2(n_1214),
.Y(n_1247)
);

NOR2x1_ASAP7_75t_L g1248 ( 
.A(n_1241),
.B(n_1215),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1234),
.Y(n_1249)
);

INVx2_ASAP7_75t_SL g1250 ( 
.A(n_1241),
.Y(n_1250)
);

AO221x2_ASAP7_75t_L g1251 ( 
.A1(n_1245),
.A2(n_1214),
.B1(n_1231),
.B2(n_1211),
.C(n_1210),
.Y(n_1251)
);

NAND2xp33_ASAP7_75t_SL g1252 ( 
.A(n_1246),
.B(n_1209),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1248),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_1252),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1250),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1249),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1255),
.B(n_1251),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1254),
.A2(n_1247),
.B1(n_1232),
.B2(n_1242),
.Y(n_1258)
);

CKINVDCx16_ASAP7_75t_R g1259 ( 
.A(n_1257),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1258),
.B(n_1256),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1257),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1257),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1262),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1261),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1260),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1259),
.B(n_1253),
.Y(n_1266)
);

INVxp67_ASAP7_75t_L g1267 ( 
.A(n_1260),
.Y(n_1267)
);

INVxp67_ASAP7_75t_L g1268 ( 
.A(n_1260),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1262),
.Y(n_1269)
);

AOI211x1_ASAP7_75t_L g1270 ( 
.A1(n_1266),
.A2(n_1238),
.B(n_1207),
.C(n_1246),
.Y(n_1270)
);

O2A1O1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1268),
.A2(n_1232),
.B(n_1082),
.C(n_1132),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1263),
.B(n_1243),
.Y(n_1272)
);

NOR2xp67_ASAP7_75t_L g1273 ( 
.A(n_1269),
.B(n_1232),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1267),
.A2(n_1244),
.B1(n_1236),
.B2(n_1237),
.Y(n_1274)
);

AOI211xp5_ASAP7_75t_L g1275 ( 
.A1(n_1265),
.A2(n_1050),
.B(n_1106),
.C(n_1233),
.Y(n_1275)
);

AO21x1_ASAP7_75t_L g1276 ( 
.A1(n_1266),
.A2(n_1056),
.B(n_1242),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1264),
.Y(n_1277)
);

AOI221xp5_ASAP7_75t_L g1278 ( 
.A1(n_1277),
.A2(n_1216),
.B1(n_1240),
.B2(n_1242),
.C(n_1208),
.Y(n_1278)
);

OAI211xp5_ASAP7_75t_L g1279 ( 
.A1(n_1270),
.A2(n_1217),
.B(n_1094),
.C(n_1084),
.Y(n_1279)
);

NOR3xp33_ASAP7_75t_L g1280 ( 
.A(n_1271),
.B(n_1076),
.C(n_1090),
.Y(n_1280)
);

OAI311xp33_ASAP7_75t_L g1281 ( 
.A1(n_1274),
.A2(n_1239),
.A3(n_1116),
.B1(n_1213),
.C1(n_1235),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1272),
.Y(n_1282)
);

AOI221xp5_ASAP7_75t_L g1283 ( 
.A1(n_1276),
.A2(n_1093),
.B1(n_1107),
.B2(n_1162),
.C(n_1092),
.Y(n_1283)
);

OAI221xp5_ASAP7_75t_L g1284 ( 
.A1(n_1273),
.A2(n_1137),
.B1(n_1231),
.B2(n_1213),
.C(n_1160),
.Y(n_1284)
);

NOR2x1_ASAP7_75t_L g1285 ( 
.A(n_1275),
.B(n_1086),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1282),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1285),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1278),
.B(n_1189),
.Y(n_1288)
);

XOR2x1_ASAP7_75t_L g1289 ( 
.A(n_1281),
.B(n_1145),
.Y(n_1289)
);

NOR2x1_ASAP7_75t_L g1290 ( 
.A(n_1279),
.B(n_1085),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1283),
.B(n_1160),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1280),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1284),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1282),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_R g1295 ( 
.A(n_1294),
.B(n_192),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1293),
.B(n_1081),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_R g1297 ( 
.A(n_1292),
.B(n_193),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1289),
.B(n_1145),
.Y(n_1298)
);

NAND3xp33_ASAP7_75t_L g1299 ( 
.A(n_1287),
.B(n_1288),
.C(n_1290),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_R g1300 ( 
.A(n_1291),
.B(n_200),
.Y(n_1300)
);

NOR3xp33_ASAP7_75t_SL g1301 ( 
.A(n_1286),
.B(n_205),
.C(n_208),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1295),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1299),
.A2(n_1153),
.B1(n_1154),
.B2(n_1155),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1298),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1301),
.B(n_1032),
.Y(n_1305)
);

O2A1O1Ixp33_ASAP7_75t_SL g1306 ( 
.A1(n_1296),
.A2(n_1089),
.B(n_1154),
.C(n_1149),
.Y(n_1306)
);

BUFx10_ASAP7_75t_L g1307 ( 
.A(n_1297),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1300),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1304),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1308),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1302),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1303),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_1307),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1310),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1311),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1313),
.A2(n_1305),
.B1(n_1306),
.B2(n_1144),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1309),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1312),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1314),
.A2(n_1144),
.B1(n_1139),
.B2(n_1136),
.Y(n_1319)
);

AOI31xp33_ASAP7_75t_L g1320 ( 
.A1(n_1318),
.A2(n_1315),
.A3(n_1317),
.B(n_1316),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1320),
.B(n_214),
.Y(n_1321)
);

AOI222xp33_ASAP7_75t_SL g1322 ( 
.A1(n_1321),
.A2(n_1319),
.B1(n_1080),
.B2(n_1075),
.C1(n_1139),
.C2(n_1136),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1322),
.Y(n_1323)
);

AOI221xp5_ASAP7_75t_L g1324 ( 
.A1(n_1323),
.A2(n_1134),
.B1(n_1114),
.B2(n_1075),
.C(n_222),
.Y(n_1324)
);

AOI211xp5_ASAP7_75t_L g1325 ( 
.A1(n_1324),
.A2(n_217),
.B(n_220),
.C(n_221),
.Y(n_1325)
);


endmodule