module fake_aes_4670_n_788 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_96, n_39, n_788);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_96;
input n_39;
output n_788;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_57), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_39), .Y(n_99) );
INVx1_ASAP7_75t_SL g100 ( .A(n_28), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_46), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_65), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_7), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_43), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_31), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_35), .Y(n_106) );
BUFx2_ASAP7_75t_L g107 ( .A(n_48), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_76), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_50), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_15), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_5), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_38), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_13), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_62), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_32), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_86), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_7), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_8), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_89), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_12), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_13), .Y(n_121) );
CKINVDCx14_ASAP7_75t_R g122 ( .A(n_67), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_85), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_94), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_96), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_92), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_95), .Y(n_127) );
INVxp33_ASAP7_75t_L g128 ( .A(n_88), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_17), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_66), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_2), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_54), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_68), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_81), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_99), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_99), .Y(n_136) );
AOI22xp5_ASAP7_75t_L g137 ( .A1(n_101), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_118), .Y(n_138) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_101), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_106), .Y(n_140) );
BUFx2_ASAP7_75t_L g141 ( .A(n_107), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_107), .B(n_3), .Y(n_142) );
INVx4_ASAP7_75t_L g143 ( .A(n_98), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_110), .B(n_4), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_104), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_106), .Y(n_146) );
OAI22x1_ASAP7_75t_R g147 ( .A1(n_103), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_102), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_102), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_115), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_124), .B(n_6), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_118), .Y(n_153) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_116), .A2(n_49), .B(n_93), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_116), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_120), .Y(n_156) );
OAI21xp33_ASAP7_75t_SL g157 ( .A1(n_145), .A2(n_110), .B(n_129), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_144), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_138), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
OR2x6_ASAP7_75t_L g161 ( .A(n_142), .B(n_129), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_143), .B(n_114), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_141), .B(n_114), .Y(n_163) );
INVx2_ASAP7_75t_SL g164 ( .A(n_141), .Y(n_164) );
INVx1_ASAP7_75t_SL g165 ( .A(n_142), .Y(n_165) );
INVx2_ASAP7_75t_SL g166 ( .A(n_142), .Y(n_166) );
NAND3xp33_ASAP7_75t_L g167 ( .A(n_152), .B(n_117), .C(n_111), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_143), .B(n_128), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_144), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_138), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_138), .Y(n_173) );
AO22x2_ASAP7_75t_L g174 ( .A1(n_148), .A2(n_155), .B1(n_149), .B2(n_151), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_148), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_135), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_143), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_156), .B(n_125), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_137), .A2(n_113), .B1(n_131), .B2(n_121), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_149), .B(n_122), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_138), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
NAND2xp33_ASAP7_75t_L g183 ( .A(n_150), .B(n_108), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_136), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_153), .Y(n_186) );
INVxp67_ASAP7_75t_L g187 ( .A(n_150), .Y(n_187) );
INVxp67_ASAP7_75t_SL g188 ( .A(n_151), .Y(n_188) );
AOI22xp33_ASAP7_75t_SL g189 ( .A1(n_147), .A2(n_121), .B1(n_120), .B2(n_118), .Y(n_189) );
OR2x6_ASAP7_75t_L g190 ( .A(n_154), .B(n_118), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_155), .B(n_118), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_139), .A2(n_134), .B1(n_133), .B2(n_125), .Y(n_192) );
BUFx10_ASAP7_75t_L g193 ( .A(n_153), .Y(n_193) );
NAND3xp33_ASAP7_75t_L g194 ( .A(n_136), .B(n_134), .C(n_133), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_174), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_174), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_170), .B(n_156), .Y(n_197) );
INVx4_ASAP7_75t_L g198 ( .A(n_174), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_174), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_163), .B(n_156), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_157), .A2(n_146), .B(n_140), .C(n_126), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_177), .B(n_109), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_187), .B(n_112), .Y(n_203) );
OAI22xp5_ASAP7_75t_SL g204 ( .A1(n_189), .A2(n_126), .B1(n_146), .B2(n_140), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_161), .A2(n_100), .B1(n_105), .B2(n_132), .Y(n_205) );
NOR2x1p5_ASAP7_75t_L g206 ( .A(n_163), .B(n_119), .Y(n_206) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_164), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_177), .B(n_123), .Y(n_208) );
INVx1_ASAP7_75t_SL g209 ( .A(n_165), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_166), .B(n_127), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_166), .B(n_130), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_180), .B(n_154), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_160), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_162), .B(n_47), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_188), .Y(n_215) );
INVxp67_ASAP7_75t_SL g216 ( .A(n_164), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_167), .B(n_51), .Y(n_217) );
AND2x2_ASAP7_75t_SL g218 ( .A(n_158), .B(n_153), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_161), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_190), .A2(n_97), .B(n_45), .Y(n_220) );
INVxp67_ASAP7_75t_SL g221 ( .A(n_168), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_161), .B(n_9), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_161), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_171), .B(n_11), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_175), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_190), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_160), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_176), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_183), .B(n_14), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_183), .B(n_14), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_192), .B(n_55), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_178), .B(n_15), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_191), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_176), .Y(n_234) );
OR2x2_ASAP7_75t_L g235 ( .A(n_179), .B(n_16), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_185), .Y(n_236) );
INVxp67_ASAP7_75t_L g237 ( .A(n_185), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_191), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_212), .A2(n_190), .B(n_194), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_199), .A2(n_190), .B1(n_159), .B2(n_181), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_213), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_221), .A2(n_181), .B(n_186), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_200), .B(n_16), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_228), .A2(n_173), .B(n_186), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_228), .A2(n_184), .B(n_182), .Y(n_245) );
NAND2x1p5_ASAP7_75t_L g246 ( .A(n_222), .B(n_17), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_215), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_213), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_234), .A2(n_184), .B(n_182), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_199), .A2(n_173), .B1(n_172), .B2(n_169), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_215), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_216), .B(n_18), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_200), .B(n_18), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_234), .A2(n_172), .B(n_169), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_226), .B(n_193), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_222), .A2(n_193), .B1(n_159), .B2(n_21), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_209), .B(n_193), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_207), .B(n_19), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_209), .B(n_237), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_238), .Y(n_260) );
AOI33xp33_ASAP7_75t_L g261 ( .A1(n_201), .A2(n_20), .A3(n_22), .B1(n_23), .B2(n_24), .B3(n_25), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_197), .A2(n_225), .B(n_211), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_238), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_225), .A2(n_26), .B(n_27), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_233), .B(n_29), .Y(n_265) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_199), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_233), .B(n_91), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_210), .A2(n_30), .B(n_33), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_227), .A2(n_34), .B(n_36), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_206), .B(n_37), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_233), .B(n_90), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_227), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_SL g273 ( .A1(n_220), .A2(n_40), .B(n_41), .C(n_42), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_247), .B(n_222), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_259), .B(n_206), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_266), .Y(n_276) );
AOI31xp67_ASAP7_75t_L g277 ( .A1(n_256), .A2(n_232), .A3(n_236), .B(n_229), .Y(n_277) );
OAI21xp5_ASAP7_75t_L g278 ( .A1(n_239), .A2(n_195), .B(n_196), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_241), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_248), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_240), .A2(n_226), .B(n_220), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_246), .A2(n_222), .B1(n_198), .B2(n_196), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_272), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_251), .B(n_235), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_262), .A2(n_226), .B(n_218), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_260), .B(n_235), .Y(n_286) );
OAI21xp5_ASAP7_75t_L g287 ( .A1(n_242), .A2(n_224), .B(n_218), .Y(n_287) );
OA21x2_ASAP7_75t_L g288 ( .A1(n_264), .A2(n_195), .B(n_230), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_266), .Y(n_289) );
BUFx10_ASAP7_75t_L g290 ( .A(n_266), .Y(n_290) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_269), .A2(n_236), .B(n_214), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_266), .B(n_198), .Y(n_292) );
AND3x1_ASAP7_75t_L g293 ( .A(n_270), .B(n_223), .C(n_231), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_L g294 ( .A1(n_252), .A2(n_217), .B(n_223), .C(n_219), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_263), .B(n_204), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_252), .B(n_204), .Y(n_296) );
AO32x2_ASAP7_75t_L g297 ( .A1(n_250), .A2(n_198), .A3(n_218), .B1(n_226), .B2(n_205), .Y(n_297) );
OA21x2_ASAP7_75t_L g298 ( .A1(n_291), .A2(n_265), .B(n_271), .Y(n_298) );
OAI21x1_ASAP7_75t_L g299 ( .A1(n_291), .A2(n_268), .B(n_267), .Y(n_299) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_281), .A2(n_246), .B(n_249), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_292), .B(n_198), .Y(n_301) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_278), .A2(n_294), .B(n_285), .Y(n_302) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_278), .A2(n_245), .B(n_244), .Y(n_303) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_287), .A2(n_273), .B(n_253), .Y(n_304) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_288), .A2(n_254), .B(n_243), .Y(n_305) );
AO31x2_ASAP7_75t_L g306 ( .A1(n_282), .A2(n_258), .A3(n_261), .B(n_273), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_283), .B(n_226), .Y(n_307) );
OAI21x1_ASAP7_75t_SL g308 ( .A1(n_283), .A2(n_257), .B(n_261), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_290), .Y(n_309) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_292), .B(n_276), .Y(n_310) );
OA21x2_ASAP7_75t_L g311 ( .A1(n_277), .A2(n_255), .B(n_258), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_283), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_279), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_279), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_296), .B(n_255), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_295), .B(n_203), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_279), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_292), .Y(n_318) );
OAI21x1_ASAP7_75t_SL g319 ( .A1(n_280), .A2(n_44), .B(n_52), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_274), .B(n_208), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_280), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_288), .A2(n_280), .B(n_274), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_312), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_312), .B(n_293), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_314), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_309), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_314), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_313), .B(n_286), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_314), .Y(n_329) );
AND2x4_ASAP7_75t_L g330 ( .A(n_301), .B(n_292), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_309), .Y(n_331) );
OAI21x1_ASAP7_75t_L g332 ( .A1(n_299), .A2(n_288), .B(n_277), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_313), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_317), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_317), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_321), .B(n_302), .Y(n_336) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_309), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_321), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_310), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_315), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_315), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_307), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_302), .B(n_293), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_316), .B(n_284), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_307), .Y(n_345) );
CKINVDCx8_ASAP7_75t_R g346 ( .A(n_301), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_307), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_322), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_316), .B(n_288), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_318), .B(n_289), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_305), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_318), .B(n_289), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_322), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_300), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_305), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_310), .Y(n_356) );
OAI21x1_ASAP7_75t_L g357 ( .A1(n_299), .A2(n_275), .B(n_276), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_320), .A2(n_276), .B1(n_290), .B2(n_202), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_320), .B(n_297), .Y(n_359) );
AO21x2_ASAP7_75t_L g360 ( .A1(n_308), .A2(n_297), .B(n_276), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_310), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_320), .B(n_297), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_325), .Y(n_363) );
NOR2x1_ASAP7_75t_SL g364 ( .A(n_356), .B(n_276), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_340), .B(n_316), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_359), .B(n_310), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_359), .B(n_301), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_351), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_334), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_334), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_337), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_326), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_335), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_362), .B(n_301), .Y(n_374) );
BUFx3_ASAP7_75t_L g375 ( .A(n_331), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_325), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_331), .Y(n_377) );
NOR2x1_ASAP7_75t_L g378 ( .A(n_331), .B(n_311), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_335), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_351), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_351), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_362), .B(n_301), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_355), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_333), .B(n_311), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_336), .B(n_300), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_323), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_333), .B(n_311), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_346), .A2(n_311), .B1(n_308), .B2(n_297), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_333), .B(n_311), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_355), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_324), .B(n_304), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_355), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_325), .Y(n_393) );
INVx3_ASAP7_75t_L g394 ( .A(n_354), .Y(n_394) );
NOR2x1p5_ASAP7_75t_L g395 ( .A(n_331), .B(n_319), .Y(n_395) );
NOR2x1_ASAP7_75t_SL g396 ( .A(n_356), .B(n_304), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_343), .A2(n_308), .B1(n_304), .B2(n_319), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_338), .B(n_305), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_338), .B(n_304), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_327), .Y(n_400) );
AND2x4_ASAP7_75t_SL g401 ( .A(n_330), .B(n_290), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_323), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_336), .B(n_300), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_324), .B(n_304), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_336), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_348), .Y(n_406) );
INVx5_ASAP7_75t_L g407 ( .A(n_354), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_348), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_338), .B(n_303), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_340), .B(n_306), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_343), .B(n_306), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_345), .B(n_303), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_353), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_353), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_327), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_345), .B(n_303), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_344), .A2(n_298), .B1(n_290), .B2(n_299), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_345), .B(n_297), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_341), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_327), .Y(n_420) );
OA21x2_ASAP7_75t_L g421 ( .A1(n_332), .A2(n_298), .B(n_306), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_342), .B(n_297), .Y(n_422) );
BUFx2_ASAP7_75t_L g423 ( .A(n_329), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_341), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_342), .B(n_306), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_349), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_349), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_329), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_347), .B(n_306), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_329), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_405), .B(n_354), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_405), .B(n_360), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_425), .B(n_360), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_369), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_369), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_425), .B(n_360), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_370), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_370), .Y(n_438) );
AND2x4_ASAP7_75t_SL g439 ( .A(n_363), .B(n_330), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_365), .B(n_347), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_406), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_365), .B(n_344), .Y(n_442) );
BUFx2_ASAP7_75t_L g443 ( .A(n_372), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_422), .B(n_360), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_367), .B(n_361), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_385), .B(n_354), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_422), .B(n_357), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_366), .B(n_357), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_373), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_373), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_379), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_366), .B(n_357), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_406), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_406), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_407), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_371), .A2(n_330), .B1(n_328), .B2(n_352), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_371), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_379), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_386), .Y(n_459) );
BUFx2_ASAP7_75t_L g460 ( .A(n_371), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_408), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_419), .B(n_352), .Y(n_462) );
AND2x4_ASAP7_75t_SL g463 ( .A(n_363), .B(n_330), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_418), .B(n_332), .Y(n_464) );
INVxp67_ASAP7_75t_L g465 ( .A(n_376), .Y(n_465) );
INVx3_ASAP7_75t_R g466 ( .A(n_415), .Y(n_466) );
BUFx3_ASAP7_75t_L g467 ( .A(n_375), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_376), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_419), .B(n_352), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_385), .B(n_354), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_386), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_408), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_374), .B(n_350), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_402), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_424), .B(n_350), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_402), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_424), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_426), .B(n_326), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_374), .B(n_361), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_408), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_367), .B(n_328), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_375), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_426), .B(n_339), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_418), .B(n_332), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_385), .B(n_354), .Y(n_485) );
NOR2xp67_ASAP7_75t_L g486 ( .A(n_407), .B(n_339), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_382), .B(n_339), .Y(n_487) );
INVxp67_ASAP7_75t_SL g488 ( .A(n_393), .Y(n_488) );
NOR2x1p5_ASAP7_75t_L g489 ( .A(n_375), .B(n_339), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_393), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_400), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_400), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_420), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_382), .B(n_385), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_427), .B(n_358), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_420), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_413), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_415), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_427), .B(n_346), .Y(n_499) );
INVx1_ASAP7_75t_SL g500 ( .A(n_401), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_401), .B(n_346), .Y(n_501) );
INVxp67_ASAP7_75t_L g502 ( .A(n_423), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_401), .B(n_298), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_423), .Y(n_504) );
INVx4_ASAP7_75t_L g505 ( .A(n_377), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_413), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_430), .B(n_306), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_412), .B(n_306), .Y(n_508) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_407), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_403), .B(n_53), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_403), .B(n_56), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_403), .B(n_298), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_403), .B(n_298), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_368), .Y(n_514) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_428), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_414), .B(n_58), .Y(n_516) );
BUFx2_ASAP7_75t_L g517 ( .A(n_377), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_412), .B(n_59), .Y(n_518) );
NAND3xp33_ASAP7_75t_L g519 ( .A(n_397), .B(n_60), .C(n_61), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_416), .B(n_63), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_377), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_430), .B(n_64), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_416), .B(n_69), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_414), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_428), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_494), .B(n_409), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_481), .B(n_428), .Y(n_527) );
INVx1_ASAP7_75t_SL g528 ( .A(n_439), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_494), .B(n_409), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_432), .B(n_411), .Y(n_530) );
OAI21xp33_ASAP7_75t_SL g531 ( .A1(n_489), .A2(n_395), .B(n_378), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_439), .A2(n_388), .B1(n_364), .B2(n_396), .Y(n_532) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_468), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_473), .B(n_398), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_434), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_479), .B(n_398), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_435), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_487), .B(n_384), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_432), .B(n_411), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_487), .B(n_384), .Y(n_540) );
INVxp67_ASAP7_75t_L g541 ( .A(n_468), .Y(n_541) );
AND2x4_ASAP7_75t_SL g542 ( .A(n_501), .B(n_394), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_433), .B(n_436), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_437), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_490), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_438), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_457), .B(n_387), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_460), .B(n_387), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_433), .B(n_410), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_449), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_463), .B(n_389), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_450), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_451), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_458), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_490), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_445), .B(n_429), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_459), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_463), .B(n_389), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_471), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_448), .B(n_399), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_436), .B(n_410), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_515), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_444), .B(n_429), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_474), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_448), .B(n_399), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_515), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_476), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_452), .B(n_378), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_504), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_455), .B(n_407), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_444), .B(n_404), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_504), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_497), .B(n_404), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_477), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_478), .B(n_391), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_465), .B(n_391), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_506), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_462), .B(n_390), .Y(n_578) );
INVx2_ASAP7_75t_SL g579 ( .A(n_443), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_469), .B(n_488), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_452), .B(n_396), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_524), .B(n_421), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_475), .B(n_390), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_495), .B(n_390), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_442), .B(n_364), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_491), .B(n_492), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_517), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_493), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_498), .Y(n_589) );
NOR2xp67_ASAP7_75t_L g590 ( .A(n_455), .B(n_407), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_455), .B(n_407), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_464), .B(n_394), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_500), .B(n_407), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_456), .A2(n_388), .B1(n_395), .B2(n_394), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_496), .Y(n_595) );
NOR2xp67_ASAP7_75t_L g596 ( .A(n_505), .B(n_394), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_483), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_441), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_464), .B(n_421), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_456), .A2(n_417), .B1(n_392), .B2(n_383), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_442), .B(n_421), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_484), .B(n_421), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_484), .B(n_392), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_447), .B(n_392), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_447), .B(n_383), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_441), .Y(n_606) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_502), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_499), .B(n_383), .Y(n_608) );
AND2x4_ASAP7_75t_L g609 ( .A(n_505), .B(n_381), .Y(n_609) );
AND2x4_ASAP7_75t_L g610 ( .A(n_505), .B(n_381), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_498), .B(n_381), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_453), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_453), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_508), .B(n_421), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_507), .B(n_380), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_454), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_440), .B(n_380), .Y(n_617) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_466), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_454), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_461), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_512), .B(n_380), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_461), .Y(n_622) );
INVx1_ASAP7_75t_SL g623 ( .A(n_618), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_618), .A2(n_511), .B1(n_510), .B2(n_521), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_543), .B(n_513), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_601), .B(n_472), .Y(n_626) );
INVx2_ASAP7_75t_SL g627 ( .A(n_579), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_585), .A2(n_601), .B1(n_594), .B2(n_581), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_586), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_526), .B(n_512), .Y(n_630) );
NOR2x1_ASAP7_75t_L g631 ( .A(n_590), .B(n_486), .Y(n_631) );
NAND3xp33_ASAP7_75t_L g632 ( .A(n_607), .B(n_519), .C(n_431), .Y(n_632) );
INVx3_ASAP7_75t_L g633 ( .A(n_570), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_543), .B(n_513), .Y(n_634) );
NAND2x1p5_ASAP7_75t_L g635 ( .A(n_528), .B(n_510), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_609), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_529), .B(n_485), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_530), .B(n_480), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_549), .B(n_472), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_530), .B(n_480), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_588), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_609), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_568), .A2(n_446), .B1(n_470), .B2(n_485), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_595), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_534), .B(n_446), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_535), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_560), .B(n_446), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_537), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_610), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_544), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_546), .Y(n_651) );
INVxp67_ASAP7_75t_L g652 ( .A(n_533), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_550), .Y(n_653) );
AND2x4_ASAP7_75t_L g654 ( .A(n_596), .B(n_467), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_552), .Y(n_655) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_533), .Y(n_656) );
OAI21xp5_ASAP7_75t_L g657 ( .A1(n_531), .A2(n_516), .B(n_510), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_545), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_565), .B(n_470), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_610), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_553), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_549), .B(n_525), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_561), .B(n_431), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_607), .B(n_431), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_561), .B(n_514), .Y(n_665) );
AND2x2_ASAP7_75t_SL g666 ( .A(n_570), .B(n_511), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_539), .B(n_467), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_538), .B(n_470), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_554), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_612), .Y(n_670) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_545), .Y(n_671) );
INVx2_ASAP7_75t_SL g672 ( .A(n_528), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_540), .B(n_485), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_536), .B(n_482), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_557), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_539), .B(n_482), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_559), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_547), .B(n_503), .Y(n_678) );
OR2x2_ASAP7_75t_L g679 ( .A(n_571), .B(n_514), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_564), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_563), .B(n_368), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_562), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_548), .B(n_511), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_567), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_574), .Y(n_685) );
OR2x2_ASAP7_75t_L g686 ( .A(n_571), .B(n_368), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_577), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_551), .B(n_520), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_580), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_563), .B(n_520), .Y(n_690) );
INVx2_ASAP7_75t_SL g691 ( .A(n_527), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_597), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_617), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_666), .A2(n_532), .B1(n_587), .B2(n_602), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_692), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_666), .A2(n_532), .B1(n_587), .B2(n_602), .Y(n_696) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_656), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_628), .B(n_541), .C(n_555), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_689), .A2(n_600), .B1(n_599), .B2(n_541), .C(n_614), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_646), .Y(n_700) );
AOI21xp33_ASAP7_75t_L g701 ( .A1(n_623), .A2(n_614), .B(n_576), .Y(n_701) );
OAI22xp5_ASAP7_75t_SL g702 ( .A1(n_623), .A2(n_657), .B1(n_627), .B2(n_635), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_629), .B(n_573), .Y(n_703) );
INVx3_ASAP7_75t_L g704 ( .A(n_654), .Y(n_704) );
OAI322xp33_ASAP7_75t_L g705 ( .A1(n_626), .A2(n_599), .A3(n_556), .B1(n_575), .B2(n_584), .C1(n_573), .C2(n_600), .Y(n_705) );
OR2x6_ASAP7_75t_L g706 ( .A(n_657), .B(n_593), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_656), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_626), .B(n_603), .Y(n_708) );
OAI31xp33_ASAP7_75t_SL g709 ( .A1(n_624), .A2(n_591), .A3(n_558), .B(n_592), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_658), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_693), .B(n_569), .Y(n_711) );
AOI311xp33_ASAP7_75t_L g712 ( .A1(n_664), .A2(n_598), .A3(n_620), .B(n_613), .C(n_606), .Y(n_712) );
AOI32xp33_ASAP7_75t_L g713 ( .A1(n_624), .A2(n_591), .A3(n_542), .B1(n_621), .B2(n_605), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_691), .B(n_572), .Y(n_714) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_658), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_647), .B(n_604), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_SL g717 ( .A1(n_664), .A2(n_518), .B(n_523), .C(n_566), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_674), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_635), .A2(n_509), .B1(n_583), .B2(n_608), .Y(n_719) );
OAI21xp5_ASAP7_75t_L g720 ( .A1(n_632), .A2(n_518), .B(n_516), .Y(n_720) );
OAI22xp33_ASAP7_75t_SL g721 ( .A1(n_633), .A2(n_578), .B1(n_582), .B2(n_615), .Y(n_721) );
OAI21xp33_ASAP7_75t_L g722 ( .A1(n_663), .A2(n_615), .B(n_582), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_672), .B(n_589), .Y(n_723) );
NAND3x2_ASAP7_75t_L g724 ( .A(n_667), .B(n_611), .C(n_516), .Y(n_724) );
INVxp33_ASAP7_75t_L g725 ( .A(n_631), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_654), .B(n_509), .Y(n_726) );
O2A1O1Ixp33_ASAP7_75t_L g727 ( .A1(n_671), .A2(n_622), .B(n_619), .C(n_616), .Y(n_727) );
AOI21xp33_ASAP7_75t_SL g728 ( .A1(n_633), .A2(n_522), .B(n_71), .Y(n_728) );
OAI21xp33_ASAP7_75t_L g729 ( .A1(n_652), .A2(n_509), .B(n_72), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_648), .Y(n_730) );
OR2x2_ASAP7_75t_L g731 ( .A(n_625), .B(n_509), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_650), .Y(n_732) );
OR2x2_ASAP7_75t_L g733 ( .A(n_634), .B(n_70), .Y(n_733) );
AOI32xp33_ASAP7_75t_L g734 ( .A1(n_688), .A2(n_87), .A3(n_74), .B1(n_75), .B2(n_77), .Y(n_734) );
INVx1_ASAP7_75t_SL g735 ( .A(n_718), .Y(n_735) );
O2A1O1Ixp33_ASAP7_75t_L g736 ( .A1(n_694), .A2(n_671), .B(n_652), .C(n_644), .Y(n_736) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_696), .A2(n_643), .B1(n_676), .B2(n_662), .C(n_639), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_700), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_730), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_699), .B(n_663), .Y(n_740) );
OAI321xp33_ASAP7_75t_L g741 ( .A1(n_702), .A2(n_690), .A3(n_641), .B1(n_662), .B2(n_639), .C(n_665), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_712), .B(n_660), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_732), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_722), .B(n_690), .Y(n_744) );
OR2x2_ASAP7_75t_L g745 ( .A(n_708), .B(n_640), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_695), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_724), .A2(n_683), .B1(n_649), .B2(n_642), .Y(n_747) );
INVxp67_ASAP7_75t_L g748 ( .A(n_697), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_706), .A2(n_636), .B1(n_665), .B2(n_681), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_706), .A2(n_630), .B1(n_638), .B2(n_678), .Y(n_750) );
AOI332xp33_ASAP7_75t_L g751 ( .A1(n_704), .A2(n_687), .A3(n_685), .B1(n_684), .B2(n_661), .B3(n_655), .C1(n_680), .C2(n_677), .Y(n_751) );
NAND2x1_ASAP7_75t_L g752 ( .A(n_706), .B(n_668), .Y(n_752) );
NAND2x1_ASAP7_75t_L g753 ( .A(n_704), .B(n_673), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_703), .B(n_651), .Y(n_754) );
AOI221xp5_ASAP7_75t_L g755 ( .A1(n_705), .A2(n_653), .B1(n_669), .B2(n_675), .C(n_681), .Y(n_755) );
AOI21xp33_ASAP7_75t_L g756 ( .A1(n_725), .A2(n_679), .B(n_686), .Y(n_756) );
NAND3xp33_ASAP7_75t_L g757 ( .A(n_736), .B(n_755), .C(n_742), .Y(n_757) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_741), .A2(n_721), .B1(n_701), .B2(n_698), .C(n_713), .Y(n_758) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_737), .B(n_709), .C(n_734), .Y(n_759) );
NOR2xp33_ASAP7_75t_SL g760 ( .A(n_735), .B(n_729), .Y(n_760) );
OAI21xp5_ASAP7_75t_SL g761 ( .A1(n_747), .A2(n_729), .B(n_720), .Y(n_761) );
NOR3xp33_ASAP7_75t_L g762 ( .A(n_741), .B(n_728), .C(n_719), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g763 ( .A(n_750), .B(n_727), .Y(n_763) );
AOI322xp5_ASAP7_75t_L g764 ( .A1(n_740), .A2(n_715), .A3(n_716), .B1(n_707), .B2(n_710), .C1(n_723), .C2(n_711), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_738), .Y(n_765) );
OAI221xp5_ASAP7_75t_L g766 ( .A1(n_752), .A2(n_717), .B1(n_726), .B2(n_714), .C(n_733), .Y(n_766) );
O2A1O1Ixp5_ASAP7_75t_L g767 ( .A1(n_753), .A2(n_682), .B(n_670), .C(n_731), .Y(n_767) );
NOR3xp33_ASAP7_75t_L g768 ( .A(n_757), .B(n_748), .C(n_744), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g769 ( .A1(n_760), .A2(n_756), .B(n_749), .Y(n_769) );
AOI21xp33_ASAP7_75t_L g770 ( .A1(n_759), .A2(n_743), .B(n_739), .Y(n_770) );
NOR2x1_ASAP7_75t_L g771 ( .A(n_761), .B(n_746), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g772 ( .A(n_767), .B(n_751), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_765), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_773), .Y(n_774) );
NAND2xp5_ASAP7_75t_SL g775 ( .A(n_768), .B(n_758), .Y(n_775) );
NOR3x1_ASAP7_75t_L g776 ( .A(n_772), .B(n_766), .C(n_763), .Y(n_776) );
NOR3xp33_ASAP7_75t_L g777 ( .A(n_775), .B(n_770), .C(n_771), .Y(n_777) );
OAI221xp5_ASAP7_75t_L g778 ( .A1(n_774), .A2(n_762), .B1(n_769), .B2(n_764), .C(n_754), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_778), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_777), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_780), .B(n_776), .Y(n_781) );
NOR2xp67_ASAP7_75t_L g782 ( .A(n_779), .B(n_745), .Y(n_782) );
OAI21xp33_ASAP7_75t_L g783 ( .A1(n_781), .A2(n_659), .B(n_645), .Y(n_783) );
AO21x2_ASAP7_75t_L g784 ( .A1(n_783), .A2(n_782), .B(n_637), .Y(n_784) );
NAND3xp33_ASAP7_75t_L g785 ( .A(n_784), .B(n_670), .C(n_78), .Y(n_785) );
OAI21xp5_ASAP7_75t_L g786 ( .A1(n_785), .A2(n_784), .B(n_79), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_786), .A2(n_73), .B1(n_80), .B2(n_82), .Y(n_787) );
OAI21xp5_ASAP7_75t_L g788 ( .A1(n_787), .A2(n_83), .B(n_84), .Y(n_788) );
endmodule