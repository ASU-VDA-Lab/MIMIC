module fake_jpeg_16856_n_246 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_246);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_246;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_149;
wire n_35;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_17),
.B1(n_19),
.B2(n_21),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_19),
.B1(n_13),
.B2(n_24),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_56),
.Y(n_78)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

OR2x2_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_19),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_59),
.Y(n_73)
);

AO22x2_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_62),
.B1(n_38),
.B2(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_13),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_21),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_19),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_13),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_19),
.Y(n_75)
);

XOR2x2_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_19),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_59),
.C(n_47),
.Y(n_87)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_59),
.B1(n_61),
.B2(n_57),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_77),
.B1(n_52),
.B2(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_76),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_43),
.B1(n_45),
.B2(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_52),
.Y(n_79)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_64),
.B(n_74),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_86),
.B(n_88),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_89),
.B1(n_96),
.B2(n_71),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_50),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_73),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_49),
.B(n_63),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_38),
.B1(n_41),
.B2(n_56),
.Y(n_89)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_58),
.B1(n_70),
.B2(n_48),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_97),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_60),
.B1(n_49),
.B2(n_58),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_51),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_77),
.B1(n_95),
.B2(n_82),
.Y(n_123)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_78),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_104),
.B(n_112),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_65),
.C(n_66),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_109),
.C(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_64),
.B(n_80),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_86),
.B(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_68),
.C(n_67),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_80),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_86),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_73),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_75),
.C(n_33),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_116),
.B(n_76),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_132),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_128),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_136),
.B(n_114),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_93),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_84),
.B1(n_95),
.B2(n_83),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_131),
.B1(n_58),
.B2(n_40),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_86),
.B1(n_82),
.B2(n_94),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_85),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_133),
.B(n_137),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_48),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_135),
.B(n_70),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_75),
.Y(n_136)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_115),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_141),
.B(n_148),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_110),
.B(n_109),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_152),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_137),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_0),
.Y(n_148)
);

NOR4xp25_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_17),
.C(n_20),
.D(n_40),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_35),
.C(n_22),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_130),
.C(n_136),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_151),
.B(n_157),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_20),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_155),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_0),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_20),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_122),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_152),
.A2(n_134),
.B1(n_125),
.B2(n_130),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_159),
.A2(n_176),
.B1(n_148),
.B2(n_143),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_122),
.Y(n_163)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_164),
.B(n_174),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_171),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_150),
.A2(n_134),
.B1(n_22),
.B2(n_16),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_169),
.B1(n_170),
.B2(n_18),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_158),
.A2(n_145),
.B1(n_146),
.B2(n_157),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_35),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_20),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_15),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_147),
.B(n_16),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_11),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_175),
.B(n_0),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_141),
.A2(n_55),
.B1(n_34),
.B2(n_16),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_172),
.A2(n_140),
.B1(n_155),
.B2(n_148),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_192),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_143),
.C(n_151),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_183),
.C(n_187),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_140),
.B1(n_155),
.B2(n_142),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_185),
.B1(n_190),
.B2(n_0),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_162),
.A2(n_24),
.B(n_22),
.Y(n_182)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_55),
.C(n_25),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_168),
.A2(n_55),
.B1(n_24),
.B2(n_18),
.Y(n_185)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_15),
.Y(n_187)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_18),
.B(n_11),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_11),
.B(n_10),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_176),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_177),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_181),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_180),
.B(n_159),
.CI(n_160),
.CON(n_194),
.SN(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_173),
.C(n_161),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_23),
.C(n_14),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_15),
.Y(n_198)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_15),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_23),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_204),
.A2(n_183),
.B1(n_190),
.B2(n_9),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_206),
.Y(n_219)
);

XNOR2x1_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_179),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_211),
.C(n_215),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_209),
.Y(n_223)
);

OAI321xp33_ASAP7_75t_L g209 ( 
.A1(n_195),
.A2(n_185),
.A3(n_187),
.B1(n_192),
.B2(n_184),
.C(n_23),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_23),
.C(n_14),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_214),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_201),
.B(n_10),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_199),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_221),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_202),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_200),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_224),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_205),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_207),
.B(n_194),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_219),
.B(n_194),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_227),
.B(n_228),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_196),
.C(n_197),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_232),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_215),
.B1(n_10),
.B2(n_3),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_218),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_14),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_234),
.B(n_236),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_217),
.B1(n_2),
.B2(n_3),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_14),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_1),
.C(n_3),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_233),
.A2(n_230),
.B(n_2),
.Y(n_238)
);

AOI322xp5_ASAP7_75t_L g241 ( 
.A1(n_238),
.A2(n_239),
.A3(n_1),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_240),
.C(n_235),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_1),
.C(n_4),
.Y(n_243)
);

OAI21x1_ASAP7_75t_L g244 ( 
.A1(n_243),
.A2(n_4),
.B(n_5),
.Y(n_244)
);

AOI221xp5_ASAP7_75t_L g245 ( 
.A1(n_244),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.C(n_239),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_245),
.A2(n_8),
.B(n_6),
.Y(n_246)
);


endmodule