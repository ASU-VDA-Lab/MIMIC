module fake_aes_8684_n_29 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_29);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
NOR2xp67_ASAP7_75t_L g10 ( .A(n_1), .B(n_2), .Y(n_10) );
BUFx10_ASAP7_75t_L g11 ( .A(n_3), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_1), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_2), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_6), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
BUFx6f_ASAP7_75t_L g16 ( .A(n_11), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_14), .B(n_0), .Y(n_17) );
OA21x2_ASAP7_75t_L g18 ( .A1(n_10), .A2(n_5), .B(n_7), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_15), .B(n_11), .Y(n_20) );
OR2x6_ASAP7_75t_L g21 ( .A(n_15), .B(n_12), .Y(n_21) );
NAND2x1p5_ASAP7_75t_L g22 ( .A(n_16), .B(n_13), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
AOI221xp5_ASAP7_75t_SL g25 ( .A1(n_24), .A2(n_17), .B1(n_16), .B2(n_22), .C(n_21), .Y(n_25) );
NAND4xp25_ASAP7_75t_L g26 ( .A(n_25), .B(n_17), .C(n_23), .D(n_21), .Y(n_26) );
NOR2xp67_ASAP7_75t_L g27 ( .A(n_26), .B(n_16), .Y(n_27) );
XNOR2xp5_ASAP7_75t_L g28 ( .A(n_27), .B(n_18), .Y(n_28) );
AOI22xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_4), .B1(n_8), .B2(n_9), .Y(n_29) );
endmodule