module fake_jpeg_21773_n_315 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_51),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_25),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_60),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_23),
.B1(n_20),
.B2(n_33),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_50),
.B1(n_23),
.B2(n_16),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_23),
.B1(n_20),
.B2(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_20),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_17),
.B(n_25),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_71),
.C(n_81),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_67),
.Y(n_112)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_17),
.B1(n_16),
.B2(n_25),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_17),
.B1(n_23),
.B2(n_16),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_90),
.B1(n_21),
.B2(n_22),
.Y(n_104)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_41),
.B(n_26),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_73),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_78),
.Y(n_122)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_47),
.B(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_29),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_83),
.Y(n_124)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_85),
.A2(n_87),
.B1(n_89),
.B2(n_91),
.Y(n_125)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_21),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_98),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_44),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_51),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_33),
.B1(n_16),
.B2(n_32),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_59),
.B(n_41),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_49),
.A2(n_33),
.B1(n_31),
.B2(n_22),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_94),
.A2(n_97),
.B1(n_35),
.B2(n_42),
.Y(n_128)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_95),
.A2(n_67),
.B1(n_84),
.B2(n_82),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_61),
.A2(n_26),
.B(n_28),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_19),
.C(n_27),
.Y(n_126)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_29),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_21),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_28),
.Y(n_114)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_114),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_104),
.A2(n_121),
.B1(n_32),
.B2(n_31),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_68),
.B1(n_76),
.B2(n_88),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_107),
.B1(n_86),
.B2(n_95),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_42),
.B1(n_35),
.B2(n_21),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_0),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_126),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_43),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_37),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_79),
.A2(n_30),
.B1(n_22),
.B2(n_31),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_99),
.B1(n_64),
.B2(n_77),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_69),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_37),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_132),
.A2(n_161),
.B(n_104),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_133),
.A2(n_139),
.B1(n_146),
.B2(n_151),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_135),
.B(n_141),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_106),
.B(n_30),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_137),
.B(n_138),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_63),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_84),
.B1(n_79),
.B2(n_80),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_101),
.B1(n_70),
.B2(n_74),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_140),
.A2(n_147),
.B1(n_110),
.B2(n_113),
.Y(n_178)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_118),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_143),
.B(n_145),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_63),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_149),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_130),
.B(n_127),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_119),
.B1(n_129),
.B2(n_131),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_115),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_148),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_109),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_97),
.B1(n_73),
.B2(n_75),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_140),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_65),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_158),
.B1(n_110),
.B2(n_34),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_103),
.B(n_64),
.C(n_43),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_159),
.C(n_122),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_107),
.Y(n_156)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_130),
.B(n_32),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_157),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_30),
.B1(n_27),
.B2(n_34),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_43),
.C(n_37),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_78),
.Y(n_160)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_114),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_169),
.C(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_151),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_146),
.A2(n_126),
.B(n_124),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_167),
.A2(n_168),
.B(n_175),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_124),
.B(n_116),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_159),
.C(n_132),
.Y(n_171)
);

A2O1A1O1Ixp25_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_116),
.B(n_37),
.C(n_28),
.D(n_24),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_24),
.C(n_162),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_122),
.B(n_113),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_190),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_161),
.A2(n_111),
.B(n_117),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_182),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_188),
.B1(n_174),
.B2(n_176),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_19),
.B(n_27),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_28),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_187),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_134),
.A2(n_19),
.B(n_28),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_139),
.A2(n_117),
.B(n_110),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_136),
.A2(n_28),
.B(n_18),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_29),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_136),
.B(n_28),
.Y(n_192)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_136),
.A2(n_18),
.B(n_24),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_193),
.A2(n_142),
.B1(n_147),
.B2(n_141),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_195),
.A2(n_210),
.B(n_214),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_198),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_170),
.B(n_148),
.Y(n_198)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_185),
.B(n_149),
.CI(n_143),
.CON(n_199),
.SN(n_199)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_199),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_200),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_164),
.A2(n_162),
.B1(n_18),
.B2(n_24),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_201),
.A2(n_213),
.B1(n_222),
.B2(n_182),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_173),
.B(n_9),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_205),
.Y(n_237)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_194),
.Y(n_206)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_165),
.Y(n_207)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

NOR2x1p5_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_18),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_208),
.A2(n_212),
.B1(n_215),
.B2(n_218),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_211),
.C(n_221),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_183),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_24),
.C(n_29),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_188),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_173),
.B(n_8),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_195),
.B1(n_217),
.B2(n_179),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_166),
.B(n_0),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_167),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_222)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_169),
.C(n_192),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_231),
.C(n_235),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_191),
.C(n_193),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_178),
.B1(n_170),
.B2(n_177),
.Y(n_233)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_168),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_220),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_172),
.C(n_163),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_163),
.C(n_189),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_238),
.C(n_240),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_189),
.C(n_184),
.Y(n_238)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_177),
.C(n_187),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_221),
.A2(n_194),
.B1(n_3),
.B2(n_4),
.Y(n_241)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_208),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_243)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_4),
.C(n_14),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_222),
.C(n_202),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_199),
.B(n_208),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_245),
.A2(n_239),
.B(n_213),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_251),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_227),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_205),
.Y(n_255)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_220),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_263),
.Y(n_275)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_259),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_226),
.A2(n_232),
.B1(n_240),
.B2(n_235),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_224),
.B1(n_241),
.B2(n_201),
.Y(n_267)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_202),
.Y(n_260)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_261),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_209),
.C(n_196),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_228),
.C(n_6),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_199),
.Y(n_263)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_264),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_276),
.C(n_262),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_247),
.B(n_248),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

NAND3xp33_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_254),
.C(n_260),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_272),
.Y(n_288)
);

OA21x2_ASAP7_75t_L g272 ( 
.A1(n_246),
.A2(n_243),
.B(n_206),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_258),
.A2(n_229),
.B1(n_206),
.B2(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_263),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_278),
.Y(n_282)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_279),
.B(n_286),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_253),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_290),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_252),
.C(n_251),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_283),
.C(n_269),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_252),
.C(n_253),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_265),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_256),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_250),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_289),
.A2(n_268),
.B1(n_264),
.B2(n_270),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_291),
.A2(n_296),
.B1(n_285),
.B2(n_287),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_275),
.Y(n_292)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_275),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_297),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_294),
.A2(n_283),
.B(n_284),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_288),
.A2(n_272),
.B1(n_276),
.B2(n_7),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_272),
.B1(n_6),
.B2(n_7),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_298),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_300),
.A2(n_299),
.B(n_295),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_303),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_298),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_302),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_307),
.Y(n_310)
);

OA21x2_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_292),
.B(n_304),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_310),
.B1(n_308),
.B2(n_305),
.Y(n_312)
);

AO21x1_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_293),
.B(n_12),
.Y(n_313)
);

MAJx2_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_14),
.C(n_11),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g315 ( 
.A(n_314),
.Y(n_315)
);


endmodule