module real_jpeg_23692_n_30 (n_17, n_8, n_0, n_21, n_168, n_2, n_29, n_10, n_9, n_12, n_24, n_165, n_166, n_170, n_6, n_28, n_161, n_162, n_169, n_167, n_23, n_11, n_14, n_160, n_25, n_163, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_164, n_16, n_15, n_13, n_30);

input n_17;
input n_8;
input n_0;
input n_21;
input n_168;
input n_2;
input n_29;
input n_10;
input n_9;
input n_12;
input n_24;
input n_165;
input n_166;
input n_170;
input n_6;
input n_28;
input n_161;
input n_162;
input n_169;
input n_167;
input n_23;
input n_11;
input n_14;
input n_160;
input n_25;
input n_163;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_164;
input n_16;
input n_15;
input n_13;

output n_30;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_64;
wire n_131;
wire n_47;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_80;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_0),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_1),
.B(n_35),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_1),
.B(n_150),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_1),
.B(n_147),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_2),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_3),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_3),
.B(n_120),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_4),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_5),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_6),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_6),
.B(n_57),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_7),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_8),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_9),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_9),
.B(n_73),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_10),
.A2(n_31),
.B(n_158),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_10),
.B(n_38),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_11),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_12),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_13),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_13),
.B(n_117),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_14),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_14),
.B(n_92),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_15),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_16),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_16),
.B(n_107),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_18),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_20),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_20),
.B(n_64),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_21),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_22),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_23),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_25),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_25),
.B(n_135),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_26),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_27),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_28),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_29),
.B(n_62),
.C(n_131),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_40),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_39),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_36),
.B(n_74),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_36),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_36),
.B(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_36),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_36),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_36),
.B(n_151),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_37),
.B(n_93),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_37),
.B(n_98),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_145),
.B(n_152),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_55),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_51),
.B(n_54),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_44),
.B(n_54),
.Y(n_155)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_47),
.B(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_48),
.Y(n_133)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_49),
.B(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_51),
.B(n_54),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_54),
.A2(n_146),
.B(n_149),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_59),
.B(n_144),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_138),
.B(n_143),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_134),
.B(n_137),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_66),
.B(n_130),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_124),
.B(n_129),
.Y(n_66)
);

OAI321xp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_116),
.A3(n_119),
.B1(n_122),
.B2(n_123),
.C(n_160),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_110),
.B(n_115),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_106),
.B(n_109),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_101),
.B(n_105),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B(n_100),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_95),
.B(n_99),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_91),
.B(n_94),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_85),
.B(n_90),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_96),
.B(n_97),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_102),
.B(n_103),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_111),
.B(n_112),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_113),
.B(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_128),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_142),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_157),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_161),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_162),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_163),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_164),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_165),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_166),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_167),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_168),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_169),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_170),
.Y(n_121)
);


endmodule