module fake_jpeg_23508_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_26),
.B(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_49),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_22),
.B(n_0),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_21),
.Y(n_86)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_60),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_64),
.Y(n_112)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_72),
.Y(n_126)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_17),
.B1(n_31),
.B2(n_32),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_80),
.B1(n_87),
.B2(n_88),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_69),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_31),
.B1(n_17),
.B2(n_36),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_33),
.B1(n_38),
.B2(n_37),
.Y(n_101)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_36),
.C(n_21),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_20),
.C(n_23),
.Y(n_98)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_74),
.Y(n_124)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_43),
.B(n_22),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_77),
.A2(n_39),
.B(n_24),
.C(n_27),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_41),
.A2(n_21),
.B1(n_32),
.B2(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_90),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_11),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_42),
.A2(n_39),
.B1(n_29),
.B2(n_27),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_52),
.A2(n_31),
.B1(n_26),
.B2(n_23),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_91),
.B(n_92),
.Y(n_100)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

NOR2x1_ASAP7_75t_SL g141 ( 
.A(n_97),
.B(n_111),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_19),
.C(n_38),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_75),
.B(n_25),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_99),
.B(n_106),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_101),
.A2(n_122),
.B1(n_119),
.B2(n_19),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_22),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_107),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_79),
.B(n_33),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_61),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_58),
.B(n_25),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_22),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_120),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_0),
.Y(n_111)
);

OR2x2_ASAP7_75t_SL g117 ( 
.A(n_59),
.B(n_15),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_119),
.B(n_18),
.Y(n_129)
);

FAx1_ASAP7_75t_SL g118 ( 
.A(n_91),
.B(n_22),
.CI(n_29),
.CON(n_118),
.SN(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_58),
.B(n_39),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_87),
.B1(n_68),
.B2(n_80),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_57),
.B(n_39),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_127),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_54),
.B(n_27),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_129),
.A2(n_150),
.B(n_141),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_134),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_133),
.B(n_152),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_115),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_91),
.B(n_34),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_135),
.A2(n_141),
.B(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_136),
.B(n_138),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_71),
.B1(n_55),
.B2(n_65),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_110),
.B(n_111),
.Y(n_170)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_142),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_54),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_140),
.B(n_155),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_149),
.A2(n_151),
.B1(n_162),
.B2(n_123),
.Y(n_191)
);

NAND2x1_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_78),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_98),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_100),
.B(n_56),
.C(n_65),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_128),
.C(n_94),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_154),
.A2(n_161),
.B1(n_108),
.B2(n_117),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_96),
.B(n_37),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_35),
.Y(n_156)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_97),
.A2(n_35),
.B1(n_34),
.B2(n_30),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_157),
.A2(n_111),
.B1(n_110),
.B2(n_103),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_103),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_159),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_160),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_101),
.A2(n_30),
.B1(n_24),
.B2(n_2),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_97),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_165),
.B(n_189),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_120),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_166),
.A2(n_170),
.B(n_171),
.Y(n_224)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_168),
.B(n_173),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_169),
.A2(n_138),
.B1(n_148),
.B2(n_149),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_118),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_175),
.C(n_190),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_150),
.A2(n_121),
.B1(n_124),
.B2(n_128),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_153),
.B1(n_144),
.B2(n_131),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_158),
.B(n_133),
.Y(n_208)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_185),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_121),
.B1(n_94),
.B2(n_24),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_184),
.A2(n_12),
.B1(n_7),
.B2(n_9),
.Y(n_227)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_187),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_123),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_135),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_191),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_129),
.B(n_8),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_14),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_136),
.A2(n_104),
.B(n_1),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_193),
.A2(n_143),
.B(n_3),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_194),
.A2(n_10),
.B1(n_5),
.B2(n_7),
.Y(n_225)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_157),
.B(n_9),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_197),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_1),
.Y(n_198)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_198),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_199),
.A2(n_211),
.B(n_220),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_162),
.B1(n_159),
.B2(n_147),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_200),
.A2(n_223),
.B1(n_194),
.B2(n_169),
.Y(n_231)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_206),
.B(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_210),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_171),
.A2(n_132),
.B(n_139),
.C(n_142),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_164),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_178),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_218),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_225),
.B1(n_227),
.B2(n_173),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_179),
.A2(n_134),
.B(n_2),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_178),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_226),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_222),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_175),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_181),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_202),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_229),
.Y(n_269)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_231),
.Y(n_252)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_242),
.Y(n_262)
);

AO22x2_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_193),
.B1(n_189),
.B2(n_184),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_233),
.A2(n_243),
.B1(n_200),
.B2(n_220),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_168),
.Y(n_235)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_235),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_180),
.Y(n_240)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_204),
.B1(n_217),
.B2(n_212),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_190),
.C(n_172),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_214),
.C(n_224),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_176),
.Y(n_247)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_247),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_224),
.A2(n_170),
.B1(n_165),
.B2(n_198),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_248),
.A2(n_211),
.B1(n_199),
.B2(n_166),
.Y(n_254)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_201),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_206),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_166),
.Y(n_250)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_235),
.C(n_240),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_254),
.A2(n_233),
.B1(n_243),
.B2(n_250),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_188),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_259),
.Y(n_271)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_188),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_233),
.B1(n_238),
.B2(n_261),
.Y(n_274)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_265),
.Y(n_272)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_248),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_233),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_234),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_268),
.Y(n_275)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_221),
.Y(n_270)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_273),
.B(n_281),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_274),
.A2(n_283),
.B1(n_254),
.B2(n_223),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_278),
.B(n_280),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_253),
.A2(n_236),
.B(n_233),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_285),
.B(n_256),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_236),
.C(n_208),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_238),
.C(n_210),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_282),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_262),
.A2(n_231),
.B1(n_249),
.B2(n_232),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_253),
.B(n_242),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_226),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_252),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_269),
.Y(n_288)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

NAND3xp33_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_263),
.C(n_203),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_290),
.A2(n_291),
.B(n_294),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_277),
.A2(n_260),
.B(n_197),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_256),
.B(n_245),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_274),
.C(n_255),
.Y(n_304)
);

BUFx12_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_296),
.B(n_298),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_297),
.A2(n_273),
.B1(n_279),
.B2(n_278),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_202),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_302),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_299),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_301),
.A2(n_304),
.B(n_307),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_292),
.A2(n_276),
.B1(n_282),
.B2(n_272),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_271),
.C(n_280),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_225),
.B1(n_227),
.B2(n_215),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_308),
.B(n_192),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_271),
.C(n_245),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_309),
.A2(n_216),
.B(n_167),
.Y(n_316)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_290),
.Y(n_311)
);

NOR2x1_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_167),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_266),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_312),
.A2(n_313),
.B(n_317),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_259),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_316),
.A2(n_303),
.B(n_306),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_296),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_319),
.B(n_320),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_296),
.B(n_187),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_322),
.B(n_314),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_317),
.B(n_177),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_321),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g327 ( 
.A1(n_325),
.A2(n_312),
.B(n_313),
.Y(n_327)
);

AOI31xp33_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_327),
.A3(n_323),
.B(n_195),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_195),
.C(n_196),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_185),
.C(n_3),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_7),
.Y(n_332)
);


endmodule