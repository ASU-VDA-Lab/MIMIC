module fake_netlist_6_1774_n_2045 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2045);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2045;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1971;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_35),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_182),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_136),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_32),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_50),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_100),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_34),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_106),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_13),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_91),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_144),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_28),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_127),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_3),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_14),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_198),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_80),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_175),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_27),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_22),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_147),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_60),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_200),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_206),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_131),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_113),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_150),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_185),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_184),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_22),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_156),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_153),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_142),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_178),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_112),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_81),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_4),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_164),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_151),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_114),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_192),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_86),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_34),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_103),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_32),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_195),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_48),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_89),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_37),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_90),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_190),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_199),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_191),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_141),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_18),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_204),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_19),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_37),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_27),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_58),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_13),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_92),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_30),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_122),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_138),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_181),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_157),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_5),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_132),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_115),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_177),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_73),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_56),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_139),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_123),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_62),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_168),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_68),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_39),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_165),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_39),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_158),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_107),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_28),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_183),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_135),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_94),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_33),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_56),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_167),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_126),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_17),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_66),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_60),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_12),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_65),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_83),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_174),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_97),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_12),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_77),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_99),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_205),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_143),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_49),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_4),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_203),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_152),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_50),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_202),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_64),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_52),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_155),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_52),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_70),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_104),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_134),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_44),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_9),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_2),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_110),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_101),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_146),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_64),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_6),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_96),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_9),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_170),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_63),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_161),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_57),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_68),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_75),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_19),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_140),
.Y(n_347)
);

BUFx5_ASAP7_75t_L g348 ( 
.A(n_197),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_7),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_11),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_36),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_154),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_130),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_7),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_162),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_54),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_3),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_176),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_71),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_5),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_63),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_119),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_65),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_82),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_163),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_87),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_76),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_128),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_41),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_72),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_20),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_29),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_121),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_20),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_55),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_48),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_24),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_116),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_23),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_42),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_207),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_74),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_193),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_102),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_15),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_73),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_188),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_2),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_44),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_61),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_95),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_145),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_201),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_46),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_166),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_25),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_189),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_18),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_171),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_120),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_66),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_71),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_149),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_25),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_74),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_55),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_0),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_1),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_196),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_248),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_209),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_248),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_352),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_248),
.Y(n_414)
);

INVxp33_ASAP7_75t_SL g415 ( 
.A(n_300),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_248),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_323),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_248),
.Y(n_418)
);

NOR2xp67_ASAP7_75t_L g419 ( 
.A(n_394),
.B(n_0),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_248),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_239),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_217),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_281),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_220),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_289),
.B(n_1),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_348),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_323),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_219),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_392),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_220),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_369),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_288),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_397),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_369),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_395),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_288),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_386),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_386),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_224),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_289),
.B(n_6),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_263),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_227),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_345),
.Y(n_443)
);

NOR2xp67_ASAP7_75t_L g444 ( 
.A(n_405),
.B(n_8),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_259),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_263),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_259),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_259),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_357),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_357),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_357),
.B(n_8),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_299),
.B(n_10),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_299),
.B(n_10),
.Y(n_453)
);

BUFx2_ASAP7_75t_SL g454 ( 
.A(n_303),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_216),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_229),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_212),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_212),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_377),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_377),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_377),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_388),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_232),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_336),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_336),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_234),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_216),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_388),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_381),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_246),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_303),
.B(n_11),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_348),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_341),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_381),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_388),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_235),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_251),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_396),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_253),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_256),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_322),
.B(n_14),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_258),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_240),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_396),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_353),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_396),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_264),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_225),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_265),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_266),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_348),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_268),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_276),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_322),
.B(n_400),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_225),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_278),
.Y(n_496)
);

NOR2xp67_ASAP7_75t_L g497 ( 
.A(n_383),
.B(n_15),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_231),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_279),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_286),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_231),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_348),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_280),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_280),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_290),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_292),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_290),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_291),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_297),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_341),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_208),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_291),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_211),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_302),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_246),
.B(n_16),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_214),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_348),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_218),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_293),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_293),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_211),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_301),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_301),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_317),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_317),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_309),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_489),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_411),
.Y(n_528)
);

AND3x2_ASAP7_75t_L g529 ( 
.A(n_425),
.B(n_383),
.C(n_238),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_515),
.B(n_246),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_410),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_515),
.B(n_283),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_445),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_447),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_447),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_410),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_412),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_R g538 ( 
.A(n_483),
.B(n_310),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_412),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_448),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_448),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_441),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_464),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_465),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_490),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_422),
.B(n_283),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_414),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_492),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_414),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_509),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_451),
.B(n_283),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_511),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_421),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_416),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_449),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_473),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_451),
.B(n_295),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_446),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_416),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_449),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_450),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_423),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_418),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_450),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_470),
.B(n_295),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_429),
.Y(n_566)
);

NAND2x1_ASAP7_75t_L g567 ( 
.A(n_457),
.B(n_400),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_485),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_SL g569 ( 
.A(n_440),
.B(n_233),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_418),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_459),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_420),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_433),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_516),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_469),
.Y(n_575)
);

AND2x6_ASAP7_75t_L g576 ( 
.A(n_494),
.B(n_383),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_R g577 ( 
.A(n_428),
.B(n_313),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_439),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_459),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_518),
.Y(n_580)
);

CKINVDCx16_ASAP7_75t_R g581 ( 
.A(n_513),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_460),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_442),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_420),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_456),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_463),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_458),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_454),
.B(n_221),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_474),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_426),
.Y(n_590)
);

CKINVDCx6p67_ASAP7_75t_R g591 ( 
.A(n_521),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_466),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_460),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_510),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_426),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_476),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_477),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_472),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_479),
.B(n_480),
.Y(n_599)
);

OAI21x1_ASAP7_75t_L g600 ( 
.A1(n_472),
.A2(n_238),
.B(n_210),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_482),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_461),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_415),
.A2(n_354),
.B1(n_356),
.B2(n_273),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_497),
.B(n_295),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_462),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_487),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_488),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_468),
.B(n_316),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_493),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_496),
.B(n_211),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_510),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_499),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_R g613 ( 
.A(n_500),
.B(n_315),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_506),
.B(n_316),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_488),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_468),
.B(n_316),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_546),
.B(n_514),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_536),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_528),
.B(n_417),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_536),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_569),
.A2(n_413),
.B1(n_435),
.B2(n_452),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_537),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_588),
.B(n_526),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_587),
.Y(n_624)
);

INVx4_ASAP7_75t_SL g625 ( 
.A(n_576),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_576),
.A2(n_453),
.B1(n_481),
.B2(n_471),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_533),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_570),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_565),
.B(n_431),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_587),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_594),
.B(n_431),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_576),
.A2(n_434),
.B1(n_454),
.B2(n_332),
.Y(n_632)
);

NOR2x1p5_ASAP7_75t_L g633 ( 
.A(n_591),
.B(n_401),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_537),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_530),
.B(n_210),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_611),
.B(n_543),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_551),
.B(n_366),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_530),
.B(n_532),
.Y(n_638)
);

AND2x6_ASAP7_75t_L g639 ( 
.A(n_530),
.B(n_366),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_587),
.Y(n_640)
);

OAI22xp33_ASAP7_75t_L g641 ( 
.A1(n_552),
.A2(n_406),
.B1(n_443),
.B2(n_332),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_534),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_582),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_537),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_570),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_584),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_532),
.B(n_366),
.Y(n_647)
);

OR2x6_ASAP7_75t_L g648 ( 
.A(n_556),
.B(n_427),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_535),
.Y(n_649)
);

NAND2xp33_ASAP7_75t_R g650 ( 
.A(n_578),
.B(n_223),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_532),
.B(n_282),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_576),
.A2(n_337),
.B1(n_360),
.B2(n_318),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_587),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_574),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_540),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_544),
.B(n_475),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_578),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_537),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_551),
.B(n_557),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_541),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_555),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_560),
.Y(n_662)
);

BUFx4f_ASAP7_75t_L g663 ( 
.A(n_591),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_537),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_584),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_575),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_580),
.A2(n_610),
.B1(n_585),
.B2(n_586),
.Y(n_667)
);

INVxp67_ASAP7_75t_SL g668 ( 
.A(n_590),
.Y(n_668)
);

INVxp33_ASAP7_75t_L g669 ( 
.A(n_603),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_551),
.B(n_228),
.Y(n_670)
);

NOR2x1p5_ASAP7_75t_L g671 ( 
.A(n_583),
.B(n_475),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_561),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_564),
.Y(n_673)
);

OR2x2_ASAP7_75t_L g674 ( 
.A(n_614),
.B(n_478),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_590),
.Y(n_675)
);

BUFx4f_ASAP7_75t_L g676 ( 
.A(n_576),
.Y(n_676)
);

INVx5_ASAP7_75t_L g677 ( 
.A(n_576),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_557),
.B(n_478),
.Y(n_678)
);

INVx4_ASAP7_75t_SL g679 ( 
.A(n_576),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_604),
.B(n_378),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_595),
.Y(n_681)
);

INVx8_ASAP7_75t_L g682 ( 
.A(n_592),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_598),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_571),
.Y(n_684)
);

INVx5_ASAP7_75t_L g685 ( 
.A(n_539),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_579),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_593),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_602),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_582),
.Y(n_689)
);

BUFx10_ASAP7_75t_L g690 ( 
.A(n_583),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_L g691 ( 
.A1(n_605),
.A2(n_337),
.B1(n_360),
.B2(n_318),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_587),
.B(n_348),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_604),
.B(n_484),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_604),
.B(n_484),
.Y(n_694)
);

BUFx8_ASAP7_75t_SL g695 ( 
.A(n_553),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_539),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_547),
.Y(n_697)
);

BUFx10_ASAP7_75t_L g698 ( 
.A(n_585),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_547),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_589),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_608),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_608),
.B(n_282),
.Y(n_702)
);

INVx5_ASAP7_75t_L g703 ( 
.A(n_539),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_599),
.B(n_486),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_542),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_616),
.B(n_486),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_538),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_586),
.B(n_455),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_572),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_600),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_608),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_539),
.Y(n_712)
);

BUFx4f_ASAP7_75t_L g713 ( 
.A(n_616),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_616),
.B(n_581),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_568),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_596),
.B(n_467),
.C(n_444),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_607),
.Y(n_717)
);

INVx6_ASAP7_75t_L g718 ( 
.A(n_554),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_577),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_531),
.B(n_549),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_554),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_SL g722 ( 
.A(n_596),
.B(n_211),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_607),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_615),
.A2(n_372),
.B1(n_376),
.B2(n_371),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_531),
.B(n_319),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_597),
.B(n_495),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_615),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_531),
.B(n_334),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_549),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_597),
.B(n_298),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_613),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_554),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_549),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_554),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_601),
.B(n_298),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_559),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_559),
.Y(n_737)
);

OR2x6_ASAP7_75t_L g738 ( 
.A(n_542),
.B(n_419),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_601),
.A2(n_609),
.B1(n_612),
.B2(n_606),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_529),
.B(n_340),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_554),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_606),
.B(n_495),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_563),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_558),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_563),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_L g746 ( 
.A(n_563),
.B(n_348),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_609),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_612),
.B(n_498),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_558),
.B(n_498),
.Y(n_749)
);

INVxp67_ASAP7_75t_SL g750 ( 
.A(n_563),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_563),
.Y(n_751)
);

AND2x6_ASAP7_75t_L g752 ( 
.A(n_600),
.B(n_213),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_527),
.B(n_311),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_SL g754 ( 
.A(n_567),
.B(n_226),
.Y(n_754)
);

OAI22xp33_ASAP7_75t_L g755 ( 
.A1(n_567),
.A2(n_372),
.B1(n_376),
.B2(n_371),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_527),
.B(n_311),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_562),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_545),
.Y(n_758)
);

INVx4_ASAP7_75t_L g759 ( 
.A(n_548),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_548),
.B(n_342),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_550),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_550),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_568),
.A2(n_379),
.B1(n_404),
.B2(n_402),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_726),
.B(n_241),
.C(n_230),
.Y(n_764)
);

NOR3xp33_ASAP7_75t_L g765 ( 
.A(n_641),
.B(n_257),
.C(n_255),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_704),
.B(n_261),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_704),
.B(n_213),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_659),
.B(n_501),
.Y(n_768)
);

AO22x1_ASAP7_75t_L g769 ( 
.A1(n_726),
.A2(n_379),
.B1(n_402),
.B2(n_404),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_676),
.B(n_348),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_638),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_617),
.B(n_215),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_675),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_629),
.B(n_501),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_617),
.B(n_215),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_666),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_659),
.B(n_711),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_659),
.B(n_222),
.Y(n_778)
);

AO22x2_ASAP7_75t_L g779 ( 
.A1(n_753),
.A2(n_314),
.B1(n_320),
.B2(n_325),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_677),
.B(n_367),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_643),
.B(n_503),
.Y(n_781)
);

NOR2x1p5_ASAP7_75t_L g782 ( 
.A(n_707),
.B(n_714),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_708),
.B(n_504),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_701),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_706),
.B(n_236),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_706),
.B(n_236),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_626),
.B(n_237),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_749),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_R g789 ( 
.A(n_707),
.B(n_566),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_742),
.B(n_267),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_678),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_677),
.B(n_367),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_L g793 ( 
.A(n_641),
.B(n_654),
.C(n_716),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_656),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_675),
.Y(n_795)
);

AND2x6_ASAP7_75t_SL g796 ( 
.A(n_648),
.B(n_504),
.Y(n_796)
);

OAI22xp33_ASAP7_75t_L g797 ( 
.A1(n_722),
.A2(n_347),
.B1(n_338),
.B2(n_335),
.Y(n_797)
);

INVx5_ASAP7_75t_L g798 ( 
.A(n_752),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_748),
.B(n_269),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_626),
.B(n_237),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_678),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_678),
.B(n_242),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_632),
.A2(n_347),
.B(n_362),
.C(n_358),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_757),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_717),
.B(n_242),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_681),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_723),
.B(n_244),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_727),
.Y(n_808)
);

INVx8_ASAP7_75t_L g809 ( 
.A(n_682),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_681),
.Y(n_810)
);

A2O1A1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_632),
.A2(n_358),
.B(n_362),
.C(n_368),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_677),
.B(n_387),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_674),
.B(n_244),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_623),
.B(n_245),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_748),
.B(n_270),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_677),
.B(n_387),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_713),
.B(n_625),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_652),
.A2(n_338),
.B1(n_368),
.B2(n_245),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_693),
.B(n_247),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_694),
.B(n_247),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_652),
.A2(n_335),
.B1(n_249),
.B2(n_250),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_627),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_642),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_710),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_619),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_R g826 ( 
.A(n_715),
.B(n_573),
.Y(n_826)
);

BUFx5_ASAP7_75t_L g827 ( 
.A(n_752),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_649),
.B(n_249),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_655),
.B(n_250),
.Y(n_829)
);

INVxp33_ASAP7_75t_L g830 ( 
.A(n_631),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_660),
.B(n_252),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_724),
.A2(n_333),
.B1(n_252),
.B2(n_254),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_661),
.B(n_254),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_662),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_672),
.Y(n_835)
);

OR2x2_ASAP7_75t_L g836 ( 
.A(n_636),
.B(n_505),
.Y(n_836)
);

INVx8_ASAP7_75t_L g837 ( 
.A(n_682),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_713),
.B(n_399),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_730),
.B(n_271),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_650),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_724),
.A2(n_260),
.B(n_262),
.C(n_274),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_673),
.Y(n_842)
);

AND2x2_ASAP7_75t_SL g843 ( 
.A(n_763),
.B(n_399),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_752),
.A2(n_333),
.B1(n_260),
.B2(n_262),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_SL g845 ( 
.A1(n_747),
.A2(n_373),
.B1(n_243),
.B2(n_409),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_670),
.A2(n_355),
.B1(n_364),
.B2(n_365),
.Y(n_846)
);

BUFx12f_ASAP7_75t_L g847 ( 
.A(n_657),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_648),
.B(n_505),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_684),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_719),
.B(n_507),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_686),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_650),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_683),
.Y(n_853)
);

INVxp67_ASAP7_75t_L g854 ( 
.A(n_705),
.Y(n_854)
);

AOI221xp5_ASAP7_75t_L g855 ( 
.A1(n_763),
.A2(n_305),
.B1(n_408),
.B2(n_407),
.C(n_398),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_687),
.B(n_274),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_647),
.A2(n_287),
.B(n_277),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_744),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_688),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_680),
.A2(n_277),
.B1(n_287),
.B2(n_294),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_668),
.B(n_294),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_753),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_637),
.B(n_314),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_637),
.B(n_320),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_637),
.B(n_325),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_621),
.A2(n_651),
.B1(n_635),
.B2(n_731),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_635),
.B(n_328),
.Y(n_867)
);

NAND3xp33_ASAP7_75t_L g868 ( 
.A(n_730),
.B(n_275),
.C(n_272),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_697),
.Y(n_869)
);

NOR3xp33_ASAP7_75t_L g870 ( 
.A(n_756),
.B(n_285),
.C(n_284),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_651),
.B(n_328),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_699),
.Y(n_872)
);

O2A1O1Ixp5_ASAP7_75t_L g873 ( 
.A1(n_702),
.A2(n_329),
.B(n_403),
.C(n_409),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_729),
.B(n_329),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_757),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_733),
.B(n_403),
.Y(n_876)
);

INVxp33_ASAP7_75t_L g877 ( 
.A(n_695),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_702),
.A2(n_517),
.B(n_502),
.C(n_491),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_735),
.B(n_296),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_618),
.Y(n_880)
);

NOR3x1_ASAP7_75t_L g881 ( 
.A(n_756),
.B(n_525),
.C(n_524),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_618),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_737),
.B(n_384),
.Y(n_883)
);

INVx4_ASAP7_75t_L g884 ( 
.A(n_624),
.Y(n_884)
);

NAND2xp33_ASAP7_75t_L g885 ( 
.A(n_639),
.B(n_391),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_679),
.B(n_393),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_735),
.B(n_304),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_710),
.B(n_491),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_710),
.B(n_502),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_709),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_643),
.B(n_507),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_620),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_689),
.B(n_508),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_628),
.Y(n_894)
);

INVx8_ASAP7_75t_L g895 ( 
.A(n_682),
.Y(n_895)
);

OR2x6_ASAP7_75t_L g896 ( 
.A(n_762),
.B(n_508),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_628),
.Y(n_897)
);

NOR2x1p5_ASAP7_75t_L g898 ( 
.A(n_760),
.B(n_306),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_648),
.B(n_512),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_709),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_689),
.B(n_307),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_740),
.B(n_308),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_695),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_725),
.B(n_312),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_728),
.B(n_321),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_671),
.B(n_512),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_SL g907 ( 
.A(n_663),
.B(n_243),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_645),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_750),
.A2(n_517),
.B(n_424),
.Y(n_909)
);

AND2x4_ASAP7_75t_SL g910 ( 
.A(n_657),
.B(n_243),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_667),
.A2(n_374),
.B1(n_327),
.B2(n_330),
.Y(n_911)
);

NOR2xp67_ASAP7_75t_L g912 ( 
.A(n_739),
.B(n_78),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_787),
.A2(n_800),
.B1(n_771),
.B2(n_766),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_766),
.B(n_639),
.Y(n_914)
);

O2A1O1Ixp5_ASAP7_75t_L g915 ( 
.A1(n_772),
.A2(n_736),
.B(n_720),
.C(n_645),
.Y(n_915)
);

O2A1O1Ixp5_ASAP7_75t_L g916 ( 
.A1(n_775),
.A2(n_736),
.B(n_665),
.C(n_646),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_789),
.Y(n_917)
);

BUFx4f_ASAP7_75t_L g918 ( 
.A(n_809),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_888),
.A2(n_710),
.B(n_630),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_888),
.A2(n_889),
.B(n_824),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_889),
.A2(n_630),
.B(n_622),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_824),
.A2(n_664),
.B(n_622),
.Y(n_922)
);

NOR2x1p5_ASAP7_75t_SL g923 ( 
.A(n_827),
.B(n_745),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_773),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_824),
.Y(n_925)
);

NOR3xp33_ASAP7_75t_L g926 ( 
.A(n_790),
.B(n_815),
.C(n_799),
.Y(n_926)
);

O2A1O1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_803),
.A2(n_755),
.B(n_691),
.C(n_692),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_799),
.B(n_634),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_798),
.B(n_657),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_783),
.B(n_690),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_824),
.A2(n_664),
.B(n_622),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_795),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_840),
.B(n_669),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_806),
.Y(n_934)
);

AO32x1_ASAP7_75t_L g935 ( 
.A1(n_860),
.A2(n_665),
.A3(n_646),
.B1(n_520),
.B2(n_522),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_777),
.A2(n_743),
.B(n_721),
.Y(n_936)
);

OAI21xp33_ASAP7_75t_L g937 ( 
.A1(n_815),
.A2(n_669),
.B(n_738),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_843),
.A2(n_752),
.B1(n_691),
.B2(n_755),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_803),
.A2(n_811),
.B(n_767),
.C(n_797),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_839),
.A2(n_754),
.B(n_663),
.C(n_758),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_804),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_810),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_SL g943 ( 
.A(n_776),
.B(n_759),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_814),
.B(n_634),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_904),
.B(n_644),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_884),
.A2(n_743),
.B(n_624),
.Y(n_946)
);

OAI321xp33_ASAP7_75t_L g947 ( 
.A1(n_797),
.A2(n_738),
.A3(n_761),
.B1(n_519),
.B2(n_520),
.C(n_525),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_852),
.B(n_690),
.Y(n_948)
);

NOR3xp33_ASAP7_75t_L g949 ( 
.A(n_793),
.B(n_759),
.C(n_754),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_884),
.A2(n_743),
.B(n_624),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_770),
.A2(n_741),
.B(n_751),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_827),
.B(n_690),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_SL g953 ( 
.A(n_847),
.B(n_759),
.Y(n_953)
);

AOI21x1_ASAP7_75t_L g954 ( 
.A1(n_780),
.A2(n_738),
.B(n_430),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_904),
.B(n_644),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_778),
.A2(n_696),
.B(n_734),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_768),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_789),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_905),
.B(n_658),
.Y(n_959)
);

BUFx12f_ASAP7_75t_L g960 ( 
.A(n_796),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_862),
.B(n_788),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_839),
.A2(n_692),
.B(n_633),
.C(n_746),
.Y(n_962)
);

BUFx4f_ASAP7_75t_L g963 ( 
.A(n_809),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_866),
.A2(n_712),
.B1(n_734),
.B2(n_732),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_774),
.B(n_698),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_844),
.A2(n_715),
.B1(n_653),
.B2(n_640),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_817),
.A2(n_640),
.B(n_653),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_858),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_843),
.B(n_696),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_850),
.B(n_808),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_863),
.A2(n_732),
.B(n_703),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_864),
.A2(n_703),
.B(n_685),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_768),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_788),
.B(n_698),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_891),
.B(n_640),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_848),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_893),
.B(n_653),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_844),
.B(n_718),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_791),
.B(n_718),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_869),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_801),
.B(n_718),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_853),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_817),
.A2(n_703),
.B(n_685),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_818),
.A2(n_375),
.B1(n_331),
.B2(n_339),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_827),
.B(n_685),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_836),
.Y(n_986)
);

OAI21xp33_ASAP7_75t_L g987 ( 
.A1(n_855),
.A2(n_380),
.B(n_343),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_885),
.A2(n_523),
.B(n_522),
.Y(n_988)
);

AOI21xp33_ASAP7_75t_L g989 ( 
.A1(n_879),
.A2(n_359),
.B(n_390),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_794),
.B(n_324),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_841),
.A2(n_523),
.B(n_438),
.C(n_437),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_822),
.B(n_326),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_827),
.B(n_243),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_838),
.A2(n_438),
.B(n_437),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_838),
.A2(n_865),
.B(n_883),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_823),
.B(n_344),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_802),
.A2(n_346),
.B(n_349),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_834),
.B(n_835),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_842),
.B(n_350),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_849),
.B(n_851),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_830),
.B(n_351),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_859),
.B(n_361),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_887),
.B(n_363),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_887),
.B(n_370),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_784),
.Y(n_1005)
);

AO22x1_ASAP7_75t_L g1006 ( 
.A1(n_765),
.A2(n_389),
.B1(n_382),
.B2(n_385),
.Y(n_1006)
);

OAI22x1_ASAP7_75t_L g1007 ( 
.A1(n_825),
.A2(n_436),
.B1(n_432),
.B2(n_430),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_854),
.B(n_424),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_899),
.B(n_16),
.Y(n_1009)
);

BUFx4f_ASAP7_75t_L g1010 ( 
.A(n_809),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_872),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_781),
.B(n_373),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_886),
.A2(n_125),
.B(n_187),
.Y(n_1013)
);

OAI321xp33_ASAP7_75t_L g1014 ( 
.A1(n_911),
.A2(n_373),
.A3(n_21),
.B1(n_23),
.B2(n_24),
.C(n_26),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_781),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_818),
.A2(n_373),
.B1(n_186),
.B2(n_179),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_896),
.B(n_17),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_902),
.A2(n_912),
.B1(n_898),
.B2(n_901),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_813),
.B(n_21),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_785),
.B(n_26),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_902),
.A2(n_173),
.B1(n_172),
.B2(n_160),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_906),
.B(n_159),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_786),
.B(n_29),
.Y(n_1023)
);

AOI21x1_ASAP7_75t_L g1024 ( 
.A1(n_792),
.A2(n_148),
.B(n_137),
.Y(n_1024)
);

AOI21x1_ASAP7_75t_L g1025 ( 
.A1(n_792),
.A2(n_133),
.B(n_124),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_841),
.A2(n_30),
.B(n_31),
.C(n_33),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_812),
.A2(n_118),
.B(n_117),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_890),
.A2(n_111),
.B(n_108),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_900),
.Y(n_1029)
);

BUFx4f_ASAP7_75t_L g1030 ( 
.A(n_837),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_901),
.A2(n_820),
.B1(n_819),
.B2(n_906),
.Y(n_1031)
);

BUFx12f_ASAP7_75t_L g1032 ( 
.A(n_782),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_867),
.A2(n_105),
.B1(n_98),
.B2(n_93),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_812),
.A2(n_88),
.B(n_85),
.Y(n_1034)
);

OAI321xp33_ASAP7_75t_L g1035 ( 
.A1(n_832),
.A2(n_36),
.A3(n_38),
.B1(n_40),
.B2(n_41),
.C(n_43),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_816),
.A2(n_84),
.B(n_79),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_857),
.A2(n_40),
.B(n_43),
.C(n_45),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_821),
.B(n_861),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_821),
.B(n_45),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_871),
.B(n_46),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_832),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_816),
.A2(n_47),
.B(n_51),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_880),
.A2(n_53),
.B(n_54),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_868),
.A2(n_764),
.B1(n_896),
.B2(n_870),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_896),
.A2(n_53),
.B1(n_57),
.B2(n_59),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_846),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_805),
.B(n_67),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_827),
.B(n_67),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_907),
.B(n_910),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_874),
.A2(n_69),
.B(n_70),
.C(n_72),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_882),
.A2(n_69),
.B(n_75),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_807),
.B(n_779),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_779),
.B(n_897),
.Y(n_1053)
);

AOI21x1_ASAP7_75t_L g1054 ( 
.A1(n_876),
.A2(n_908),
.B(n_894),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_873),
.A2(n_892),
.B(n_856),
.C(n_828),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_878),
.A2(n_909),
.B(n_833),
.Y(n_1056)
);

AOI33xp33_ASAP7_75t_L g1057 ( 
.A1(n_845),
.A2(n_769),
.A3(n_881),
.B1(n_779),
.B2(n_826),
.B3(n_877),
.Y(n_1057)
);

AOI21x1_ASAP7_75t_L g1058 ( 
.A1(n_829),
.A2(n_831),
.B(n_875),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_837),
.B(n_895),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_837),
.A2(n_895),
.B(n_903),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_826),
.B(n_895),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_776),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_888),
.A2(n_676),
.B(n_713),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_766),
.B(n_704),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_766),
.B(n_704),
.Y(n_1065)
);

BUFx4f_ASAP7_75t_L g1066 ( 
.A(n_809),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_888),
.A2(n_676),
.B(n_713),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_SL g1068 ( 
.A(n_903),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_840),
.B(n_852),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_776),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_930),
.B(n_965),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_980),
.Y(n_1073)
);

NAND2x1_ASAP7_75t_L g1074 ( 
.A(n_925),
.B(n_924),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_926),
.B(n_913),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_920),
.A2(n_1054),
.B(n_919),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_926),
.A2(n_969),
.B(n_914),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_932),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_922),
.A2(n_931),
.B(n_967),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_1063),
.A2(n_1067),
.B(n_921),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_970),
.B(n_1003),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_934),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_1070),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1004),
.B(n_1031),
.Y(n_1084)
);

AO21x1_ASAP7_75t_L g1085 ( 
.A1(n_1048),
.A2(n_1037),
.B(n_1052),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_916),
.A2(n_936),
.B(n_915),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_938),
.A2(n_939),
.B(n_1035),
.C(n_1014),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_986),
.B(n_1062),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_938),
.A2(n_1038),
.B1(n_1018),
.B2(n_928),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_915),
.A2(n_995),
.B(n_1056),
.Y(n_1090)
);

AO31x2_ASAP7_75t_L g1091 ( 
.A1(n_1053),
.A2(n_1055),
.A3(n_1050),
.B(n_1020),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_951),
.A2(n_950),
.B(n_946),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_985),
.A2(n_983),
.B(n_956),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_942),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_978),
.A2(n_964),
.B(n_962),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_975),
.A2(n_977),
.B(n_944),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_1058),
.A2(n_979),
.B(n_981),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_998),
.B(n_1000),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_947),
.B(n_937),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_971),
.A2(n_972),
.B(n_993),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_961),
.B(n_1019),
.Y(n_1101)
);

OAI21xp33_ASAP7_75t_L g1102 ( 
.A1(n_989),
.A2(n_987),
.B(n_990),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_961),
.B(n_1069),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1024),
.A2(n_1025),
.B(n_954),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_1011),
.A2(n_1029),
.B(n_1013),
.Y(n_1105)
);

INVxp67_ASAP7_75t_SL g1106 ( 
.A(n_925),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_933),
.B(n_949),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_949),
.B(n_1023),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_925),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_952),
.A2(n_966),
.B(n_1028),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_973),
.B(n_1044),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_927),
.A2(n_1039),
.B(n_1046),
.C(n_1009),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1048),
.A2(n_1040),
.B(n_1047),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1022),
.A2(n_929),
.B(n_988),
.Y(n_1114)
);

BUFx12f_ASAP7_75t_L g1115 ( 
.A(n_1032),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1062),
.B(n_976),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1009),
.B(n_1005),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_982),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_968),
.Y(n_1119)
);

OR2x6_ASAP7_75t_L g1120 ( 
.A(n_1060),
.B(n_941),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1005),
.B(n_957),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1005),
.B(n_997),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_SL g1123 ( 
.A1(n_1026),
.A2(n_1041),
.B(n_1042),
.Y(n_1123)
);

OA22x2_ASAP7_75t_L g1124 ( 
.A1(n_976),
.A2(n_974),
.B1(n_1007),
.B2(n_1045),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1012),
.A2(n_973),
.B(n_940),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_973),
.B(n_1005),
.Y(n_1126)
);

BUFx5_ASAP7_75t_L g1127 ( 
.A(n_923),
.Y(n_1127)
);

OA22x2_ASAP7_75t_L g1128 ( 
.A1(n_948),
.A2(n_958),
.B1(n_984),
.B2(n_1061),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_918),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1015),
.B(n_1057),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_917),
.Y(n_1131)
);

AOI21xp33_ASAP7_75t_L g1132 ( 
.A1(n_1001),
.A2(n_990),
.B(n_1002),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1017),
.A2(n_1016),
.B(n_1021),
.C(n_1049),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_SL g1134 ( 
.A1(n_1043),
.A2(n_1051),
.B(n_1034),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_1017),
.A2(n_1049),
.B(n_991),
.C(n_1033),
.Y(n_1135)
);

INVxp67_ASAP7_75t_L g1136 ( 
.A(n_1008),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1001),
.B(n_943),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_992),
.A2(n_996),
.B(n_999),
.C(n_994),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1027),
.A2(n_1036),
.B(n_1059),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_SL g1140 ( 
.A1(n_935),
.A2(n_918),
.B(n_1066),
.Y(n_1140)
);

INVx3_ASAP7_75t_SL g1141 ( 
.A(n_1015),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_973),
.A2(n_1010),
.B(n_1066),
.C(n_963),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_963),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_935),
.A2(n_1015),
.B(n_1010),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1015),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1030),
.A2(n_953),
.B(n_935),
.C(n_1006),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1030),
.A2(n_1068),
.B(n_960),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1068),
.B(n_930),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1064),
.A2(n_1065),
.B(n_926),
.C(n_766),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_958),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_924),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_958),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1064),
.A2(n_1065),
.B1(n_926),
.B2(n_913),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1064),
.A2(n_1065),
.B(n_926),
.C(n_766),
.Y(n_1157)
);

AOI21x1_ASAP7_75t_L g1158 ( 
.A1(n_945),
.A2(n_959),
.B(n_955),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_913),
.A2(n_1052),
.A3(n_800),
.B(n_787),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1070),
.B(n_776),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_1062),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1064),
.A2(n_1065),
.B(n_926),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_SL g1165 ( 
.A1(n_1028),
.A2(n_927),
.B(n_1037),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_SL g1166 ( 
.A1(n_1028),
.A2(n_927),
.B(n_1037),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1064),
.A2(n_1065),
.B(n_926),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_913),
.A2(n_1052),
.A3(n_800),
.B(n_787),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_914),
.A2(n_676),
.B(n_798),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1064),
.A2(n_1065),
.B(n_926),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_924),
.Y(n_1173)
);

BUFx4f_ASAP7_75t_L g1174 ( 
.A(n_1032),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_1062),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_920),
.A2(n_919),
.B(n_1054),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_924),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_920),
.A2(n_919),
.B(n_1054),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1064),
.A2(n_1065),
.B1(n_926),
.B2(n_913),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1064),
.A2(n_1065),
.B(n_926),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_920),
.A2(n_1054),
.B(n_919),
.Y(n_1183)
);

AOI21x1_ASAP7_75t_L g1184 ( 
.A1(n_945),
.A2(n_959),
.B(n_955),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1064),
.A2(n_1065),
.B1(n_926),
.B2(n_913),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_1062),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1064),
.A2(n_1065),
.B(n_926),
.C(n_766),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_930),
.B(n_965),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_925),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_926),
.A2(n_1065),
.B1(n_1064),
.B2(n_766),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_973),
.B(n_791),
.Y(n_1192)
);

AOI221x1_ASAP7_75t_L g1193 ( 
.A1(n_926),
.A2(n_949),
.B1(n_1064),
.B2(n_1065),
.C(n_913),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_924),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1062),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_920),
.A2(n_919),
.B(n_1054),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_914),
.A2(n_676),
.B(n_798),
.Y(n_1199)
);

OA21x2_ASAP7_75t_L g1200 ( 
.A1(n_915),
.A2(n_916),
.B(n_956),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1064),
.A2(n_1065),
.B1(n_926),
.B2(n_913),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_920),
.A2(n_919),
.B(n_1054),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1062),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1064),
.A2(n_1065),
.B(n_926),
.C(n_766),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_980),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_925),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1161),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1196),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1072),
.B(n_1189),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_1083),
.Y(n_1212)
);

NAND3xp33_ASAP7_75t_L g1213 ( 
.A(n_1191),
.B(n_1157),
.C(n_1149),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1087),
.A2(n_1167),
.B1(n_1160),
.B2(n_1208),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1190),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1120),
.B(n_1129),
.Y(n_1216)
);

AND2x6_ASAP7_75t_L g1217 ( 
.A(n_1190),
.B(n_1192),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1203),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1116),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1131),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1102),
.A2(n_1075),
.B1(n_1163),
.B2(n_1172),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1149),
.A2(n_1157),
.B(n_1188),
.C(n_1204),
.Y(n_1222)
);

OR2x6_ASAP7_75t_L g1223 ( 
.A(n_1120),
.B(n_1147),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1073),
.Y(n_1224)
);

INVx5_ASAP7_75t_L g1225 ( 
.A(n_1190),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1160),
.B(n_1167),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1137),
.B(n_1088),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1120),
.B(n_1129),
.Y(n_1228)
);

CKINVDCx8_ASAP7_75t_R g1229 ( 
.A(n_1131),
.Y(n_1229)
);

NOR2xp67_ASAP7_75t_L g1230 ( 
.A(n_1150),
.B(n_1154),
.Y(n_1230)
);

AO21x2_ASAP7_75t_L g1231 ( 
.A1(n_1075),
.A2(n_1110),
.B(n_1100),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1190),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1119),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1071),
.B(n_1151),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1143),
.B(n_1142),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1084),
.A2(n_1095),
.B(n_1096),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1162),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1152),
.B(n_1155),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1109),
.Y(n_1239)
);

CKINVDCx11_ASAP7_75t_R g1240 ( 
.A(n_1115),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1156),
.A2(n_1201),
.B(n_1186),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1168),
.A2(n_1182),
.B1(n_1181),
.B2(n_1099),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1132),
.B(n_1164),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1177),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1187),
.Y(n_1245)
);

BUFx12f_ASAP7_75t_L g1246 ( 
.A(n_1115),
.Y(n_1246)
);

NOR4xp25_ASAP7_75t_L g1247 ( 
.A(n_1188),
.B(n_1204),
.C(n_1087),
.D(n_1133),
.Y(n_1247)
);

INVxp67_ASAP7_75t_SL g1248 ( 
.A(n_1106),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1107),
.A2(n_1175),
.B1(n_1205),
.B2(n_1197),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1109),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1098),
.A2(n_1089),
.B(n_1165),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1169),
.B(n_1176),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1185),
.B(n_1195),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1166),
.A2(n_1081),
.B(n_1077),
.Y(n_1254)
);

INVx5_ASAP7_75t_L g1255 ( 
.A(n_1207),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1143),
.B(n_1142),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1174),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1193),
.B(n_1101),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1192),
.B(n_1145),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1192),
.B(n_1148),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1136),
.B(n_1103),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1174),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1114),
.A2(n_1090),
.B(n_1199),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1099),
.A2(n_1128),
.B1(n_1124),
.B2(n_1111),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1130),
.B(n_1124),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1128),
.B(n_1117),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1108),
.B(n_1150),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1206),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1141),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1121),
.B(n_1111),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_SL g1271 ( 
.A1(n_1154),
.A2(n_1141),
.B1(n_1122),
.B2(n_1113),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1207),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1078),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1112),
.A2(n_1133),
.B(n_1135),
.C(n_1138),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1074),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1078),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1135),
.B(n_1173),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1082),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1082),
.Y(n_1279)
);

BUFx12f_ASAP7_75t_L g1280 ( 
.A(n_1125),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1094),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1094),
.B(n_1173),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1126),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1123),
.A2(n_1085),
.B1(n_1118),
.B2(n_1179),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1159),
.B(n_1170),
.Y(n_1285)
);

INVx3_ASAP7_75t_R g1286 ( 
.A(n_1153),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1153),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1159),
.B(n_1170),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1179),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1159),
.B(n_1170),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1194),
.B(n_1091),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1194),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1138),
.B(n_1126),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1140),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1159),
.B(n_1170),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1106),
.B(n_1105),
.Y(n_1296)
);

INVx5_ASAP7_75t_L g1297 ( 
.A(n_1127),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1091),
.B(n_1158),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1091),
.B(n_1139),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1171),
.A2(n_1080),
.B(n_1092),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1144),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1134),
.A2(n_1079),
.B(n_1200),
.Y(n_1302)
);

OR2x6_ASAP7_75t_L g1303 ( 
.A(n_1097),
.B(n_1093),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1184),
.B(n_1127),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1127),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1146),
.B(n_1076),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1146),
.A2(n_1200),
.B1(n_1086),
.B2(n_1183),
.Y(n_1307)
);

AND2x6_ASAP7_75t_L g1308 ( 
.A(n_1104),
.B(n_1178),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1180),
.B(n_1198),
.Y(n_1309)
);

O2A1O1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1202),
.A2(n_926),
.B(n_1065),
.C(n_1064),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1087),
.A2(n_1065),
.B1(n_1064),
.B2(n_1160),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1196),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1120),
.B(n_1129),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1072),
.B(n_930),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1160),
.B(n_1167),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1087),
.A2(n_1065),
.B1(n_1064),
.B2(n_1160),
.Y(n_1316)
);

CKINVDCx11_ASAP7_75t_R g1317 ( 
.A(n_1115),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1160),
.B(n_1167),
.Y(n_1318)
);

INVx4_ASAP7_75t_L g1319 ( 
.A(n_1141),
.Y(n_1319)
);

INVx4_ASAP7_75t_L g1320 ( 
.A(n_1141),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1073),
.Y(n_1321)
);

BUFx12f_ASAP7_75t_L g1322 ( 
.A(n_1115),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1160),
.A2(n_926),
.B(n_1065),
.C(n_1064),
.Y(n_1323)
);

BUFx3_ASAP7_75t_L g1324 ( 
.A(n_1196),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1190),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1196),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_SL g1327 ( 
.A(n_1150),
.B(n_776),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1196),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1160),
.B(n_1167),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1072),
.B(n_930),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1196),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1073),
.Y(n_1332)
);

NAND2x1p5_ASAP7_75t_L g1333 ( 
.A(n_1190),
.B(n_824),
.Y(n_1333)
);

CKINVDCx16_ASAP7_75t_R g1334 ( 
.A(n_1115),
.Y(n_1334)
);

AND2x6_ASAP7_75t_L g1335 ( 
.A(n_1190),
.B(n_1192),
.Y(n_1335)
);

INVx4_ASAP7_75t_L g1336 ( 
.A(n_1141),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1160),
.B(n_1167),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1160),
.B(n_1167),
.Y(n_1338)
);

INVx4_ASAP7_75t_L g1339 ( 
.A(n_1141),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1073),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1146),
.A2(n_1085),
.A3(n_1193),
.B(n_1089),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1150),
.Y(n_1342)
);

BUFx8_ASAP7_75t_SL g1343 ( 
.A(n_1115),
.Y(n_1343)
);

INVx1_ASAP7_75t_SL g1344 ( 
.A(n_1161),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1072),
.B(n_930),
.Y(n_1345)
);

OAI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1191),
.A2(n_1065),
.B1(n_1064),
.B2(n_722),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1161),
.B(n_700),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1129),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1160),
.B(n_1167),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1129),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1102),
.A2(n_926),
.B1(n_421),
.B2(n_423),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1087),
.A2(n_1065),
.B1(n_1064),
.B2(n_1160),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1160),
.B(n_1167),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1120),
.B(n_1129),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_1240),
.Y(n_1355)
);

BUFx10_ASAP7_75t_L g1356 ( 
.A(n_1342),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1243),
.A2(n_1213),
.B1(n_1311),
.B2(n_1352),
.Y(n_1357)
);

CKINVDCx11_ASAP7_75t_R g1358 ( 
.A(n_1317),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1225),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_SL g1360 ( 
.A1(n_1311),
.A2(n_1316),
.B1(n_1352),
.B2(n_1214),
.Y(n_1360)
);

INVx6_ASAP7_75t_L g1361 ( 
.A(n_1225),
.Y(n_1361)
);

INVxp67_ASAP7_75t_SL g1362 ( 
.A(n_1248),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1235),
.B(n_1256),
.Y(n_1363)
);

BUFx10_ASAP7_75t_L g1364 ( 
.A(n_1269),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1265),
.B(n_1249),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_1225),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1226),
.A2(n_1337),
.B1(n_1338),
.B2(n_1329),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1269),
.Y(n_1368)
);

AO21x2_ASAP7_75t_L g1369 ( 
.A1(n_1300),
.A2(n_1302),
.B(n_1263),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1297),
.Y(n_1370)
);

CKINVDCx8_ASAP7_75t_R g1371 ( 
.A(n_1269),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1282),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1270),
.Y(n_1373)
);

INVx6_ASAP7_75t_L g1374 ( 
.A(n_1348),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1268),
.Y(n_1375)
);

BUFx12f_ASAP7_75t_L g1376 ( 
.A(n_1246),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1312),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1321),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1348),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1332),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1346),
.A2(n_1242),
.B1(n_1221),
.B2(n_1316),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1214),
.A2(n_1241),
.B1(n_1267),
.B2(n_1266),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1241),
.A2(n_1280),
.B1(n_1271),
.B2(n_1211),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1270),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1226),
.B(n_1315),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1340),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1314),
.A2(n_1330),
.B1(n_1345),
.B2(n_1264),
.Y(n_1387)
);

AOI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1309),
.A2(n_1236),
.B(n_1307),
.Y(n_1388)
);

NAND2x1p5_ASAP7_75t_L g1389 ( 
.A(n_1297),
.B(n_1216),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1219),
.Y(n_1390)
);

AO21x1_ASAP7_75t_SL g1391 ( 
.A1(n_1285),
.A2(n_1290),
.B(n_1295),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1323),
.B(n_1234),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1278),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1279),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1281),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1289),
.Y(n_1396)
);

BUFx4f_ASAP7_75t_SL g1397 ( 
.A(n_1322),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1289),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1315),
.B(n_1318),
.Y(n_1399)
);

CKINVDCx11_ASAP7_75t_R g1400 ( 
.A(n_1229),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1234),
.B(n_1238),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1227),
.A2(n_1277),
.B1(n_1254),
.B2(n_1349),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_R g1403 ( 
.A(n_1220),
.B(n_1327),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1212),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1318),
.A2(n_1337),
.B1(n_1353),
.B2(n_1329),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1292),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1291),
.Y(n_1407)
);

NAND2x1_ASAP7_75t_L g1408 ( 
.A(n_1223),
.B(n_1216),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1348),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1326),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1247),
.B(n_1285),
.Y(n_1411)
);

INVx8_ASAP7_75t_L g1412 ( 
.A(n_1217),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1238),
.A2(n_1252),
.B1(n_1253),
.B2(n_1235),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1252),
.B(n_1253),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1276),
.A2(n_1287),
.B1(n_1209),
.B2(n_1344),
.Y(n_1415)
);

AO21x2_ASAP7_75t_L g1416 ( 
.A1(n_1304),
.A2(n_1293),
.B(n_1307),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1273),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1261),
.B(n_1258),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1347),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1350),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1258),
.B(n_1254),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1283),
.Y(n_1422)
);

OA21x2_ASAP7_75t_L g1423 ( 
.A1(n_1288),
.A2(n_1295),
.B(n_1290),
.Y(n_1423)
);

INVx2_ASAP7_75t_SL g1424 ( 
.A(n_1210),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1328),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1256),
.B(n_1259),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1228),
.A2(n_1354),
.B1(n_1313),
.B2(n_1260),
.Y(n_1427)
);

BUFx12f_ASAP7_75t_L g1428 ( 
.A(n_1350),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1350),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1283),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1259),
.B(n_1354),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1251),
.A2(n_1313),
.B1(n_1228),
.B2(n_1223),
.Y(n_1432)
);

INVx3_ASAP7_75t_SL g1433 ( 
.A(n_1334),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1239),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1239),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1260),
.A2(n_1223),
.B1(n_1230),
.B2(n_1218),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1297),
.Y(n_1437)
);

AOI21xp33_ASAP7_75t_L g1438 ( 
.A1(n_1274),
.A2(n_1310),
.B(n_1222),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1245),
.B(n_1233),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1250),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1250),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1272),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1272),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1324),
.B(n_1331),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1231),
.A2(n_1294),
.B1(n_1299),
.B2(n_1306),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1237),
.Y(n_1446)
);

NAND2x1p5_ASAP7_75t_L g1447 ( 
.A(n_1319),
.B(n_1339),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1231),
.A2(n_1299),
.B1(n_1244),
.B2(n_1284),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1255),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1286),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1215),
.Y(n_1451)
);

CKINVDCx12_ASAP7_75t_R g1452 ( 
.A(n_1343),
.Y(n_1452)
);

BUFx2_ASAP7_75t_R g1453 ( 
.A(n_1257),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1215),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1232),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1262),
.B(n_1319),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1341),
.B(n_1222),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1232),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1274),
.A2(n_1304),
.B(n_1298),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1296),
.A2(n_1217),
.B1(n_1335),
.B2(n_1320),
.Y(n_1460)
);

INVx6_ASAP7_75t_L g1461 ( 
.A(n_1320),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1325),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1217),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1217),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1296),
.A2(n_1217),
.B1(n_1335),
.B2(n_1339),
.Y(n_1465)
);

OR2x6_ASAP7_75t_L g1466 ( 
.A(n_1303),
.B(n_1305),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1335),
.A2(n_1336),
.B1(n_1301),
.B2(n_1275),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1325),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1336),
.B(n_1335),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1333),
.A2(n_1308),
.B(n_1303),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1335),
.Y(n_1471)
);

CKINVDCx11_ASAP7_75t_R g1472 ( 
.A(n_1275),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1303),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1255),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1308),
.A2(n_1255),
.B1(n_1333),
.B2(n_1341),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1255),
.Y(n_1476)
);

NAND2x1p5_ASAP7_75t_L g1477 ( 
.A(n_1308),
.B(n_1297),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1308),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_SL g1479 ( 
.A1(n_1308),
.A2(n_669),
.B1(n_1243),
.B2(n_1049),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1249),
.B(n_1243),
.Y(n_1480)
);

BUFx8_ASAP7_75t_SL g1481 ( 
.A(n_1343),
.Y(n_1481)
);

CKINVDCx11_ASAP7_75t_R g1482 ( 
.A(n_1240),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1224),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1243),
.A2(n_722),
.B1(n_1137),
.B2(n_421),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1224),
.Y(n_1485)
);

OAI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1351),
.A2(n_722),
.B1(n_1065),
.B2(n_1064),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1225),
.Y(n_1487)
);

CKINVDCx6p67_ASAP7_75t_R g1488 ( 
.A(n_1240),
.Y(n_1488)
);

BUFx2_ASAP7_75t_R g1489 ( 
.A(n_1343),
.Y(n_1489)
);

INVx6_ASAP7_75t_L g1490 ( 
.A(n_1225),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1247),
.B(n_1213),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1212),
.Y(n_1492)
);

NAND2x1p5_ASAP7_75t_L g1493 ( 
.A(n_1297),
.B(n_1225),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1243),
.A2(n_926),
.B1(n_1102),
.B2(n_1065),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1269),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1243),
.A2(n_926),
.B1(n_1102),
.B2(n_1065),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1243),
.A2(n_926),
.B1(n_1102),
.B2(n_1065),
.Y(n_1497)
);

OAI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1351),
.A2(n_722),
.B1(n_1065),
.B2(n_1064),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1312),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1390),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1390),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1372),
.Y(n_1502)
);

AOI21xp33_ASAP7_75t_L g1503 ( 
.A1(n_1486),
.A2(n_1498),
.B(n_1496),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1461),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1477),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1401),
.B(n_1414),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1407),
.Y(n_1507)
);

INVx3_ASAP7_75t_L g1508 ( 
.A(n_1477),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1389),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1461),
.Y(n_1510)
);

BUFx2_ASAP7_75t_SL g1511 ( 
.A(n_1371),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1407),
.B(n_1457),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1372),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1411),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1411),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1423),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1423),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1389),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1423),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1480),
.B(n_1404),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1421),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1421),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1457),
.B(n_1418),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_1377),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1470),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1481),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1408),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1418),
.B(n_1365),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1491),
.A2(n_1436),
.B1(n_1385),
.B2(n_1399),
.Y(n_1529)
);

AO21x2_ASAP7_75t_L g1530 ( 
.A1(n_1369),
.A2(n_1438),
.B(n_1388),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1459),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1492),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_1410),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1401),
.B(n_1414),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1466),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1466),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1473),
.B(n_1466),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1466),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1373),
.B(n_1384),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1473),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1363),
.B(n_1478),
.Y(n_1541)
);

BUFx8_ASAP7_75t_SL g1542 ( 
.A(n_1481),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1392),
.B(n_1367),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1461),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1416),
.Y(n_1545)
);

INVx3_ASAP7_75t_L g1546 ( 
.A(n_1470),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1461),
.Y(n_1547)
);

INVx1_ASAP7_75t_SL g1548 ( 
.A(n_1425),
.Y(n_1548)
);

OAI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1494),
.A2(n_1497),
.B(n_1357),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1416),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1384),
.B(n_1491),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1416),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1369),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1369),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1363),
.B(n_1432),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1463),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1360),
.B(n_1382),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1363),
.B(n_1391),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1395),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_1370),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1391),
.B(n_1402),
.Y(n_1561)
);

BUFx2_ASAP7_75t_L g1562 ( 
.A(n_1362),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1479),
.B(n_1445),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1406),
.Y(n_1564)
);

BUFx12f_ASAP7_75t_L g1565 ( 
.A(n_1358),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1405),
.B(n_1419),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1370),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1381),
.B(n_1393),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1387),
.B(n_1413),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1426),
.B(n_1375),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1394),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1499),
.Y(n_1572)
);

OAI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1484),
.A2(n_1383),
.B(n_1415),
.Y(n_1573)
);

OA21x2_ASAP7_75t_L g1574 ( 
.A1(n_1448),
.A2(n_1475),
.B(n_1380),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1426),
.B(n_1378),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1422),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1426),
.B(n_1437),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1386),
.B(n_1483),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1485),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1430),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1364),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1463),
.Y(n_1582)
);

INVx4_ASAP7_75t_L g1583 ( 
.A(n_1412),
.Y(n_1583)
);

INVx2_ASAP7_75t_SL g1584 ( 
.A(n_1364),
.Y(n_1584)
);

AO21x2_ASAP7_75t_L g1585 ( 
.A1(n_1437),
.A2(n_1474),
.B(n_1442),
.Y(n_1585)
);

NAND3xp33_ASAP7_75t_L g1586 ( 
.A(n_1450),
.B(n_1467),
.C(n_1427),
.Y(n_1586)
);

AO21x2_ASAP7_75t_L g1587 ( 
.A1(n_1434),
.A2(n_1441),
.B(n_1435),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1471),
.A2(n_1493),
.B(n_1465),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1471),
.B(n_1431),
.Y(n_1589)
);

OA21x2_ASAP7_75t_L g1590 ( 
.A1(n_1396),
.A2(n_1398),
.B(n_1443),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1431),
.B(n_1439),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1476),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1412),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1440),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1451),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1454),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1412),
.Y(n_1597)
);

INVxp67_ASAP7_75t_L g1598 ( 
.A(n_1446),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1455),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1458),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1462),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1468),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1431),
.B(n_1417),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1449),
.Y(n_1604)
);

INVx2_ASAP7_75t_SL g1605 ( 
.A(n_1364),
.Y(n_1605)
);

OR2x6_ASAP7_75t_L g1606 ( 
.A(n_1525),
.B(n_1412),
.Y(n_1606)
);

OAI33xp33_ASAP7_75t_L g1607 ( 
.A1(n_1566),
.A2(n_1444),
.A3(n_1469),
.B1(n_1464),
.B2(n_1371),
.B3(n_1488),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1514),
.B(n_1433),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1500),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1501),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1537),
.B(n_1460),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1506),
.B(n_1424),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1527),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1523),
.B(n_1512),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1523),
.B(n_1424),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1512),
.B(n_1495),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1532),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1562),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1521),
.B(n_1522),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1514),
.B(n_1433),
.Y(n_1620)
);

AOI222xp33_ASAP7_75t_L g1621 ( 
.A1(n_1549),
.A2(n_1358),
.B1(n_1482),
.B2(n_1397),
.C1(n_1376),
.C2(n_1400),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1521),
.B(n_1368),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1522),
.B(n_1368),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1534),
.B(n_1403),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1525),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1528),
.B(n_1515),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1562),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1528),
.B(n_1429),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1535),
.Y(n_1629)
);

OA21x2_ASAP7_75t_L g1630 ( 
.A1(n_1552),
.A2(n_1456),
.B(n_1493),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1533),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1515),
.B(n_1379),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1520),
.B(n_1453),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1559),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1592),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1559),
.Y(n_1636)
);

NAND3xp33_ASAP7_75t_L g1637 ( 
.A(n_1503),
.B(n_1472),
.C(n_1482),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1572),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1551),
.B(n_1420),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1502),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1564),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1564),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1531),
.B(n_1420),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1543),
.B(n_1409),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1513),
.Y(n_1645)
);

NOR2x1_ASAP7_75t_L g1646 ( 
.A(n_1585),
.B(n_1487),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1548),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1590),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1537),
.B(n_1409),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1590),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1531),
.B(n_1379),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1551),
.B(n_1429),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1557),
.A2(n_1488),
.B1(n_1376),
.B2(n_1400),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1590),
.Y(n_1654)
);

AOI221xp5_ASAP7_75t_L g1655 ( 
.A1(n_1573),
.A2(n_1447),
.B1(n_1355),
.B2(n_1359),
.C(n_1487),
.Y(n_1655)
);

CKINVDCx12_ASAP7_75t_R g1656 ( 
.A(n_1542),
.Y(n_1656)
);

INVxp67_ASAP7_75t_SL g1657 ( 
.A(n_1571),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1561),
.B(n_1374),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1561),
.B(n_1374),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1535),
.Y(n_1660)
);

INVxp67_ASAP7_75t_L g1661 ( 
.A(n_1591),
.Y(n_1661)
);

INVx1_ASAP7_75t_SL g1662 ( 
.A(n_1603),
.Y(n_1662)
);

BUFx2_ASAP7_75t_L g1663 ( 
.A(n_1536),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1536),
.B(n_1447),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1558),
.B(n_1366),
.Y(n_1665)
);

NAND2x1_ASAP7_75t_L g1666 ( 
.A(n_1505),
.B(n_1490),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1557),
.A2(n_1472),
.B1(n_1355),
.B2(n_1356),
.Y(n_1667)
);

INVxp33_ASAP7_75t_L g1668 ( 
.A(n_1603),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1563),
.A2(n_1569),
.B1(n_1555),
.B2(n_1529),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1570),
.B(n_1356),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1538),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1563),
.A2(n_1356),
.B1(n_1428),
.B2(n_1361),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1537),
.B(n_1546),
.Y(n_1673)
);

OAI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1637),
.A2(n_1586),
.B1(n_1568),
.B2(n_1583),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1637),
.A2(n_1511),
.B1(n_1568),
.B2(n_1555),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1614),
.B(n_1558),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1614),
.B(n_1537),
.Y(n_1677)
);

AOI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1607),
.A2(n_1524),
.B1(n_1598),
.B2(n_1570),
.C(n_1575),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1658),
.B(n_1539),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1661),
.B(n_1539),
.Y(n_1680)
);

NAND4xp25_ASAP7_75t_L g1681 ( 
.A(n_1669),
.B(n_1579),
.C(n_1578),
.D(n_1594),
.Y(n_1681)
);

OAI21xp5_ASAP7_75t_SL g1682 ( 
.A1(n_1621),
.A2(n_1555),
.B(n_1593),
.Y(n_1682)
);

OAI21xp5_ASAP7_75t_SL g1683 ( 
.A1(n_1655),
.A2(n_1555),
.B(n_1593),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1626),
.B(n_1540),
.Y(n_1684)
);

NAND3xp33_ASAP7_75t_L g1685 ( 
.A(n_1608),
.B(n_1540),
.C(n_1592),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1608),
.B(n_1574),
.C(n_1576),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1657),
.B(n_1578),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1638),
.B(n_1507),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1609),
.B(n_1507),
.Y(n_1689)
);

OAI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1633),
.A2(n_1588),
.B(n_1580),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1658),
.B(n_1541),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1624),
.A2(n_1565),
.B1(n_1574),
.B2(n_1511),
.Y(n_1692)
);

INVx2_ASAP7_75t_SL g1693 ( 
.A(n_1613),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1610),
.B(n_1594),
.Y(n_1694)
);

NAND3xp33_ASAP7_75t_L g1695 ( 
.A(n_1620),
.B(n_1574),
.C(n_1577),
.Y(n_1695)
);

OAI21xp33_ASAP7_75t_L g1696 ( 
.A1(n_1620),
.A2(n_1518),
.B(n_1509),
.Y(n_1696)
);

AND2x2_ASAP7_75t_SL g1697 ( 
.A(n_1630),
.B(n_1525),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1619),
.B(n_1546),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_SL g1699 ( 
.A1(n_1667),
.A2(n_1509),
.B1(n_1518),
.B2(n_1582),
.C(n_1556),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1619),
.B(n_1546),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1672),
.A2(n_1588),
.B(n_1577),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_SL g1702 ( 
.A1(n_1653),
.A2(n_1565),
.B1(n_1452),
.B2(n_1526),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1618),
.B(n_1627),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1615),
.B(n_1525),
.Y(n_1704)
);

NAND3xp33_ASAP7_75t_L g1705 ( 
.A(n_1644),
.B(n_1574),
.C(n_1577),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1640),
.B(n_1602),
.Y(n_1706)
);

OAI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1670),
.A2(n_1583),
.B1(n_1593),
.B2(n_1597),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1645),
.B(n_1587),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1612),
.B(n_1587),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1617),
.A2(n_1577),
.B1(n_1541),
.B2(n_1589),
.Y(n_1710)
);

OAI21xp33_ASAP7_75t_L g1711 ( 
.A1(n_1668),
.A2(n_1518),
.B(n_1509),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1631),
.A2(n_1541),
.B1(n_1589),
.B2(n_1583),
.Y(n_1712)
);

NOR3xp33_ASAP7_75t_L g1713 ( 
.A(n_1643),
.B(n_1508),
.C(n_1505),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1632),
.B(n_1647),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1632),
.B(n_1587),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1611),
.A2(n_1541),
.B1(n_1589),
.B2(n_1583),
.Y(n_1716)
);

OAI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1664),
.A2(n_1504),
.B1(n_1547),
.B2(n_1544),
.C(n_1510),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1611),
.A2(n_1597),
.B1(n_1582),
.B2(n_1556),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1611),
.A2(n_1597),
.B1(n_1582),
.B2(n_1556),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1659),
.B(n_1525),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1662),
.B(n_1596),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1622),
.B(n_1596),
.Y(n_1722)
);

OAI221xp5_ASAP7_75t_SL g1723 ( 
.A1(n_1643),
.A2(n_1599),
.B1(n_1545),
.B2(n_1550),
.C(n_1516),
.Y(n_1723)
);

NAND3xp33_ASAP7_75t_L g1724 ( 
.A(n_1651),
.B(n_1604),
.C(n_1567),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1622),
.B(n_1599),
.Y(n_1725)
);

OAI21xp5_ASAP7_75t_SL g1726 ( 
.A1(n_1611),
.A2(n_1593),
.B(n_1589),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1634),
.Y(n_1727)
);

OA21x2_ASAP7_75t_L g1728 ( 
.A1(n_1648),
.A2(n_1554),
.B(n_1553),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1664),
.B(n_1505),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1628),
.A2(n_1593),
.B1(n_1530),
.B2(n_1600),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1623),
.B(n_1595),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1616),
.B(n_1639),
.Y(n_1732)
);

NAND3xp33_ASAP7_75t_L g1733 ( 
.A(n_1646),
.B(n_1560),
.C(n_1567),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1616),
.B(n_1601),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1673),
.B(n_1517),
.Y(n_1735)
);

OA21x2_ASAP7_75t_L g1736 ( 
.A1(n_1648),
.A2(n_1654),
.B(n_1650),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1639),
.B(n_1585),
.Y(n_1737)
);

NOR3xp33_ASAP7_75t_L g1738 ( 
.A(n_1666),
.B(n_1508),
.C(n_1510),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1656),
.A2(n_1452),
.B1(n_1428),
.B2(n_1504),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1736),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1674),
.B(n_1649),
.Y(n_1741)
);

AND2x4_ASAP7_75t_SL g1742 ( 
.A(n_1738),
.B(n_1606),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1727),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1709),
.B(n_1636),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1736),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1715),
.B(n_1629),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1736),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1728),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1735),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1708),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1698),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1698),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1737),
.B(n_1629),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1697),
.B(n_1625),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1733),
.B(n_1625),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1700),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1703),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1697),
.B(n_1519),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1675),
.A2(n_1649),
.B1(n_1652),
.B2(n_1665),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1689),
.B(n_1687),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1700),
.B(n_1695),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1676),
.B(n_1630),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1688),
.B(n_1660),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1677),
.B(n_1630),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1731),
.B(n_1660),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1706),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1694),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1684),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1678),
.B(n_1649),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1685),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1677),
.B(n_1630),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1722),
.B(n_1663),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1684),
.B(n_1641),
.Y(n_1773)
);

AND2x4_ASAP7_75t_L g1774 ( 
.A(n_1720),
.B(n_1606),
.Y(n_1774)
);

CKINVDCx16_ASAP7_75t_R g1775 ( 
.A(n_1702),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1704),
.B(n_1730),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1730),
.B(n_1671),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1725),
.B(n_1635),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1721),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1734),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1680),
.B(n_1642),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1701),
.B(n_1606),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1743),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1743),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1745),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1762),
.B(n_1679),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1768),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1768),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1757),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1745),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1762),
.B(n_1691),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1769),
.A2(n_1682),
.B1(n_1683),
.B2(n_1681),
.Y(n_1792)
);

OAI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1775),
.A2(n_1699),
.B1(n_1692),
.B2(n_1716),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1740),
.Y(n_1794)
);

INVx3_ASAP7_75t_L g1795 ( 
.A(n_1755),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1773),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1773),
.Y(n_1797)
);

NOR3xp33_ASAP7_75t_L g1798 ( 
.A(n_1775),
.B(n_1717),
.C(n_1690),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1746),
.B(n_1705),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1740),
.Y(n_1800)
);

NOR2xp67_ASAP7_75t_L g1801 ( 
.A(n_1770),
.B(n_1686),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1747),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1770),
.B(n_1714),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1762),
.B(n_1764),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1746),
.B(n_1732),
.Y(n_1805)
);

NOR2xp67_ASAP7_75t_R g1806 ( 
.A(n_1767),
.B(n_1613),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1747),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1751),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1757),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1751),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1752),
.Y(n_1811)
);

INVxp67_ASAP7_75t_SL g1812 ( 
.A(n_1758),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1747),
.Y(n_1813)
);

NOR3xp33_ASAP7_75t_L g1814 ( 
.A(n_1741),
.B(n_1739),
.C(n_1696),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1752),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1782),
.A2(n_1726),
.B1(n_1692),
.B2(n_1711),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1764),
.B(n_1693),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1748),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1748),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1756),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1771),
.B(n_1693),
.Y(n_1821)
);

NOR2x1_ASAP7_75t_L g1822 ( 
.A(n_1767),
.B(n_1724),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1756),
.Y(n_1823)
);

BUFx2_ASAP7_75t_L g1824 ( 
.A(n_1755),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1742),
.B(n_1713),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1744),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1744),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1749),
.Y(n_1828)
);

AOI32xp33_ASAP7_75t_L g1829 ( 
.A1(n_1777),
.A2(n_1707),
.A3(n_1729),
.B1(n_1719),
.B2(n_1718),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1753),
.B(n_1723),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_SL g1831 ( 
.A(n_1782),
.B(n_1489),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1753),
.B(n_1750),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1783),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1802),
.Y(n_1834)
);

A2O1A1Ixp33_ASAP7_75t_L g1835 ( 
.A1(n_1792),
.A2(n_1782),
.B(n_1777),
.C(n_1742),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1783),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1784),
.Y(n_1837)
);

INVxp67_ASAP7_75t_L g1838 ( 
.A(n_1803),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1830),
.B(n_1750),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1830),
.B(n_1772),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1784),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1824),
.B(n_1771),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1832),
.B(n_1772),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1801),
.B(n_1776),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1802),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1789),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1798),
.B(n_1776),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1809),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1832),
.B(n_1765),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1828),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1828),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1807),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1787),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1787),
.Y(n_1854)
);

INVxp67_ASAP7_75t_SL g1855 ( 
.A(n_1822),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1788),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1814),
.B(n_1776),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1807),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1799),
.B(n_1765),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1799),
.B(n_1779),
.Y(n_1860)
);

INVx1_ASAP7_75t_SL g1861 ( 
.A(n_1824),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1788),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1808),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1813),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1813),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1796),
.B(n_1763),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1808),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1810),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1796),
.B(n_1763),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1797),
.B(n_1778),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1810),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1812),
.B(n_1771),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1811),
.Y(n_1873)
);

AOI21xp33_ASAP7_75t_L g1874 ( 
.A1(n_1793),
.A2(n_1782),
.B(n_1759),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1811),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1795),
.B(n_1761),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1815),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1794),
.Y(n_1878)
);

INVx2_ASAP7_75t_SL g1879 ( 
.A(n_1795),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1815),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1805),
.B(n_1779),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1805),
.B(n_1766),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1797),
.B(n_1766),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1820),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1826),
.B(n_1780),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_1795),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1855),
.B(n_1825),
.Y(n_1887)
);

INVxp67_ASAP7_75t_L g1888 ( 
.A(n_1857),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1879),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1879),
.Y(n_1890)
);

INVx3_ASAP7_75t_SL g1891 ( 
.A(n_1861),
.Y(n_1891)
);

INVxp67_ASAP7_75t_L g1892 ( 
.A(n_1844),
.Y(n_1892)
);

INVxp67_ASAP7_75t_L g1893 ( 
.A(n_1847),
.Y(n_1893)
);

INVx1_ASAP7_75t_SL g1894 ( 
.A(n_1840),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1868),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1833),
.Y(n_1896)
);

BUFx3_ASAP7_75t_L g1897 ( 
.A(n_1846),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1874),
.A2(n_1782),
.B1(n_1831),
.B2(n_1825),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1876),
.B(n_1825),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1886),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1838),
.B(n_1791),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1836),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1886),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1840),
.B(n_1791),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1839),
.B(n_1786),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1839),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1837),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1848),
.B(n_1786),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1859),
.B(n_1826),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1841),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1835),
.B(n_1656),
.Y(n_1911)
);

INVx1_ASAP7_75t_SL g1912 ( 
.A(n_1859),
.Y(n_1912)
);

INVxp67_ASAP7_75t_L g1913 ( 
.A(n_1860),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1850),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1835),
.B(n_1761),
.Y(n_1915)
);

INVx1_ASAP7_75t_SL g1916 ( 
.A(n_1876),
.Y(n_1916)
);

INVx1_ASAP7_75t_SL g1917 ( 
.A(n_1878),
.Y(n_1917)
);

INVx1_ASAP7_75t_SL g1918 ( 
.A(n_1843),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1881),
.B(n_1816),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1851),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1853),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1854),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1882),
.B(n_1760),
.Y(n_1923)
);

INVxp67_ASAP7_75t_L g1924 ( 
.A(n_1883),
.Y(n_1924)
);

INVx3_ASAP7_75t_L g1925 ( 
.A(n_1842),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1842),
.B(n_1804),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1896),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1891),
.B(n_1894),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1891),
.B(n_1843),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1896),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_L g1931 ( 
.A(n_1911),
.B(n_1885),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1912),
.B(n_1829),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1925),
.Y(n_1933)
);

AOI21xp33_ASAP7_75t_L g1934 ( 
.A1(n_1893),
.A2(n_1888),
.B(n_1892),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1902),
.Y(n_1935)
);

AOI31xp33_ASAP7_75t_L g1936 ( 
.A1(n_1906),
.A2(n_1849),
.A3(n_1872),
.B(n_1869),
.Y(n_1936)
);

OAI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1915),
.A2(n_1898),
.B1(n_1891),
.B2(n_1919),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1897),
.B(n_1849),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1887),
.B(n_1872),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1887),
.B(n_1817),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1918),
.B(n_1878),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1897),
.B(n_1870),
.Y(n_1942)
);

NOR3xp33_ASAP7_75t_L g1943 ( 
.A(n_1913),
.B(n_1845),
.C(n_1834),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_SL g1944 ( 
.A(n_1916),
.B(n_1777),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_L g1945 ( 
.A(n_1924),
.B(n_1870),
.Y(n_1945)
);

OAI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1916),
.A2(n_1761),
.B1(n_1742),
.B2(n_1866),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1923),
.B(n_1895),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1902),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1907),
.Y(n_1949)
);

INVx1_ASAP7_75t_SL g1950 ( 
.A(n_1899),
.Y(n_1950)
);

AOI32xp33_ASAP7_75t_L g1951 ( 
.A1(n_1899),
.A2(n_1761),
.A3(n_1804),
.B1(n_1754),
.B2(n_1821),
.Y(n_1951)
);

HB1xp67_ASAP7_75t_L g1952 ( 
.A(n_1925),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1895),
.B(n_1827),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1904),
.B(n_1827),
.Y(n_1954)
);

XNOR2x1_ASAP7_75t_L g1955 ( 
.A(n_1917),
.B(n_1760),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1939),
.B(n_1925),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1952),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1950),
.B(n_1901),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1942),
.B(n_1905),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1940),
.B(n_1889),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1942),
.B(n_1889),
.Y(n_1961)
);

OAI22xp5_ASAP7_75t_L g1962 ( 
.A1(n_1936),
.A2(n_1908),
.B1(n_1926),
.B2(n_1917),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1933),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1933),
.B(n_1890),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1928),
.B(n_1890),
.Y(n_1965)
);

NOR2x1_ASAP7_75t_L g1966 ( 
.A(n_1929),
.B(n_1900),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1955),
.B(n_1900),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1927),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1955),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1930),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1935),
.Y(n_1971)
);

HB1xp67_ASAP7_75t_L g1972 ( 
.A(n_1941),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1938),
.B(n_1903),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1947),
.B(n_1909),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1945),
.B(n_1903),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1945),
.B(n_1926),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1932),
.B(n_1907),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1941),
.B(n_1909),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1948),
.Y(n_1979)
);

AOI21xp33_ASAP7_75t_L g1980 ( 
.A1(n_1972),
.A2(n_1937),
.B(n_1932),
.Y(n_1980)
);

NAND3xp33_ASAP7_75t_L g1981 ( 
.A(n_1966),
.B(n_1934),
.C(n_1943),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1957),
.Y(n_1982)
);

AOI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1969),
.A2(n_1944),
.B1(n_1931),
.B2(n_1946),
.Y(n_1983)
);

OAI32xp33_ASAP7_75t_L g1984 ( 
.A1(n_1969),
.A2(n_1977),
.A3(n_1962),
.B1(n_1967),
.B2(n_1978),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1956),
.Y(n_1985)
);

O2A1O1Ixp5_ASAP7_75t_SL g1986 ( 
.A1(n_1963),
.A2(n_1949),
.B(n_1914),
.C(n_1920),
.Y(n_1986)
);

AOI211xp5_ASAP7_75t_L g1987 ( 
.A1(n_1967),
.A2(n_1931),
.B(n_1953),
.C(n_1954),
.Y(n_1987)
);

NAND3xp33_ASAP7_75t_SL g1988 ( 
.A(n_1975),
.B(n_1951),
.C(n_1914),
.Y(n_1988)
);

AOI221xp5_ASAP7_75t_L g1989 ( 
.A1(n_1974),
.A2(n_1922),
.B1(n_1921),
.B2(n_1920),
.C(n_1910),
.Y(n_1989)
);

OAI211xp5_ASAP7_75t_L g1990 ( 
.A1(n_1978),
.A2(n_1921),
.B(n_1922),
.C(n_1910),
.Y(n_1990)
);

O2A1O1Ixp33_ASAP7_75t_L g1991 ( 
.A1(n_1965),
.A2(n_1800),
.B(n_1794),
.C(n_1834),
.Y(n_1991)
);

AOI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1959),
.A2(n_1806),
.B(n_1800),
.Y(n_1992)
);

AND2x4_ASAP7_75t_SL g1993 ( 
.A(n_1961),
.B(n_1774),
.Y(n_1993)
);

XNOR2xp5_ASAP7_75t_L g1994 ( 
.A(n_1976),
.B(n_1666),
.Y(n_1994)
);

NAND4xp25_ASAP7_75t_L g1995 ( 
.A(n_1980),
.B(n_1973),
.C(n_1958),
.D(n_1961),
.Y(n_1995)
);

OA22x2_ASAP7_75t_L g1996 ( 
.A1(n_1983),
.A2(n_1957),
.B1(n_1956),
.B2(n_1963),
.Y(n_1996)
);

NOR3xp33_ASAP7_75t_L g1997 ( 
.A(n_1981),
.B(n_1970),
.C(n_1968),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1985),
.B(n_1960),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1987),
.B(n_1960),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1982),
.Y(n_2000)
);

NAND3xp33_ASAP7_75t_L g2001 ( 
.A(n_1986),
.B(n_1964),
.C(n_1968),
.Y(n_2001)
);

NOR2x1p5_ASAP7_75t_L g2002 ( 
.A(n_1988),
.B(n_1971),
.Y(n_2002)
);

NAND4xp75_ASAP7_75t_L g2003 ( 
.A(n_1992),
.B(n_1964),
.C(n_1979),
.D(n_1971),
.Y(n_2003)
);

NOR2x1_ASAP7_75t_L g2004 ( 
.A(n_1990),
.B(n_1979),
.Y(n_2004)
);

AOI211x1_ASAP7_75t_L g2005 ( 
.A1(n_1984),
.A2(n_1862),
.B(n_1863),
.C(n_1856),
.Y(n_2005)
);

NOR3x1_ASAP7_75t_L g2006 ( 
.A(n_1994),
.B(n_1869),
.C(n_1866),
.Y(n_2006)
);

BUFx3_ASAP7_75t_L g2007 ( 
.A(n_1993),
.Y(n_2007)
);

OA211x2_ASAP7_75t_L g2008 ( 
.A1(n_1999),
.A2(n_1989),
.B(n_1991),
.C(n_1781),
.Y(n_2008)
);

AO21x1_ASAP7_75t_L g2009 ( 
.A1(n_1997),
.A2(n_1852),
.B(n_1845),
.Y(n_2009)
);

NOR4xp25_ASAP7_75t_L g2010 ( 
.A(n_2001),
.B(n_1995),
.C(n_2000),
.D(n_1998),
.Y(n_2010)
);

OA211x2_ASAP7_75t_L g2011 ( 
.A1(n_1996),
.A2(n_2002),
.B(n_2003),
.C(n_2004),
.Y(n_2011)
);

AOI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_2000),
.A2(n_1858),
.B(n_1852),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_SL g2013 ( 
.A(n_2007),
.B(n_1867),
.Y(n_2013)
);

NOR3xp33_ASAP7_75t_L g2014 ( 
.A(n_2006),
.B(n_1864),
.C(n_1858),
.Y(n_2014)
);

NOR2x1p5_ASAP7_75t_L g2015 ( 
.A(n_2011),
.B(n_2005),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_2009),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_2013),
.B(n_2010),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_2008),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_2014),
.B(n_1871),
.Y(n_2019)
);

AOI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_2012),
.A2(n_1864),
.B1(n_1865),
.B2(n_1880),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_2009),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2009),
.Y(n_2022)
);

AOI221xp5_ASAP7_75t_L g2023 ( 
.A1(n_2017),
.A2(n_1865),
.B1(n_1877),
.B2(n_1875),
.C(n_1873),
.Y(n_2023)
);

NAND4xp75_ASAP7_75t_L g2024 ( 
.A(n_2016),
.B(n_1884),
.C(n_1584),
.D(n_1605),
.Y(n_2024)
);

AOI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_2015),
.A2(n_2018),
.B1(n_2021),
.B2(n_2022),
.Y(n_2025)
);

INVx5_ASAP7_75t_L g2026 ( 
.A(n_2019),
.Y(n_2026)
);

OAI221xp5_ASAP7_75t_L g2027 ( 
.A1(n_2020),
.A2(n_1785),
.B1(n_1790),
.B2(n_1818),
.C(n_1819),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_2019),
.Y(n_2028)
);

AND3x2_ASAP7_75t_L g2029 ( 
.A(n_2016),
.B(n_1790),
.C(n_1785),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_2025),
.B(n_1818),
.Y(n_2030)
);

AND3x4_ASAP7_75t_L g2031 ( 
.A(n_2024),
.B(n_1774),
.C(n_1755),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2029),
.Y(n_2032)
);

NAND3xp33_ASAP7_75t_L g2033 ( 
.A(n_2026),
.B(n_1819),
.C(n_1820),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2032),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_2030),
.Y(n_2035)
);

HB1xp67_ASAP7_75t_L g2036 ( 
.A(n_2034),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_2036),
.Y(n_2037)
);

BUFx2_ASAP7_75t_L g2038 ( 
.A(n_2036),
.Y(n_2038)
);

OAI22x1_ASAP7_75t_L g2039 ( 
.A1(n_2038),
.A2(n_2026),
.B1(n_2028),
.B2(n_2035),
.Y(n_2039)
);

AOI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_2037),
.A2(n_2023),
.B(n_2033),
.Y(n_2040)
);

OAI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_2040),
.A2(n_2027),
.B(n_2031),
.Y(n_2041)
);

OAI21x1_ASAP7_75t_L g2042 ( 
.A1(n_2041),
.A2(n_2039),
.B(n_1821),
.Y(n_2042)
);

HB1xp67_ASAP7_75t_L g2043 ( 
.A(n_2042),
.Y(n_2043)
);

OAI221xp5_ASAP7_75t_R g2044 ( 
.A1(n_2043),
.A2(n_1712),
.B1(n_1716),
.B2(n_1710),
.C(n_1823),
.Y(n_2044)
);

AOI211xp5_ASAP7_75t_L g2045 ( 
.A1(n_2044),
.A2(n_1605),
.B(n_1584),
.C(n_1581),
.Y(n_2045)
);


endmodule