module fake_jpeg_2376_n_179 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_179);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_5),
.B(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_25),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_3),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g60 ( 
.A(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_51),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_19),
.B(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_69),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_1),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_54),
.B1(n_60),
.B2(n_59),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_73),
.A2(n_74),
.B1(n_66),
.B2(n_52),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_62),
.B1(n_61),
.B2(n_47),
.Y(n_74)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_45),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_81),
.B(n_62),
.Y(n_88)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_46),
.B1(n_49),
.B2(n_52),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_70),
.B(n_67),
.Y(n_87)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_84),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_101),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_92),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_71),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_48),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_48),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_98),
.Y(n_114)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_41),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_60),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_56),
.C(n_18),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_112),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_85),
.B1(n_78),
.B2(n_72),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_101),
.A2(n_76),
.B1(n_58),
.B2(n_55),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_94),
.B1(n_99),
.B2(n_5),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_50),
.B(n_22),
.Y(n_115)
);

AOI21x1_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_4),
.B(n_6),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_116),
.B(n_120),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_118),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_44),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_2),
.C(n_4),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_40),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_36),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_1),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_125),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_135),
.C(n_6),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_99),
.B1(n_39),
.B2(n_37),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_136),
.B(n_137),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_120),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_138),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

AOI322xp5_ASAP7_75t_SL g157 ( 
.A1(n_139),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_15),
.Y(n_157)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

OAI221xp5_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_141),
.B1(n_107),
.B2(n_110),
.C(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_137),
.B1(n_124),
.B2(n_13),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_31),
.B(n_26),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_148),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_151),
.C(n_152),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_132),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_24),
.C(n_23),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_7),
.C(n_8),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_7),
.C(n_8),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_154),
.B(n_9),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_131),
.B(n_16),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_156),
.B(n_11),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_157),
.A2(n_15),
.B1(n_142),
.B2(n_150),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_159),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_163),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_144),
.B1(n_154),
.B2(n_153),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_162),
.B(n_160),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_148),
.C(n_145),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_155),
.C(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_164),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_157),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_172),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_169),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_165),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_174),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_168),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_178),
.B(n_173),
.Y(n_179)
);


endmodule