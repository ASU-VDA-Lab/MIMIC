module fake_netlist_6_1307_n_37 (n_7, n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_9, n_8, n_37);

input n_7;
input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;
input n_9;
input n_8;

output n_37;

wire n_16;
wire n_34;
wire n_10;
wire n_18;
wire n_24;
wire n_21;
wire n_15;
wire n_33;
wire n_27;
wire n_14;
wire n_32;
wire n_36;
wire n_22;
wire n_26;
wire n_13;
wire n_35;
wire n_11;
wire n_28;
wire n_17;
wire n_23;
wire n_12;
wire n_20;
wire n_30;
wire n_19;
wire n_29;
wire n_31;
wire n_25;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx5p33_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx5p33_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

AND2x4_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_R g20 ( 
.A(n_14),
.B(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

OR2x6_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_16),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_R g23 ( 
.A(n_12),
.B(n_1),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_10),
.B1(n_13),
.B2(n_15),
.Y(n_24)
);

AOI221xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_10),
.B1(n_18),
.B2(n_2),
.C(n_4),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

OAI31xp33_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_19),
.A3(n_20),
.B(n_21),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_26),
.Y(n_29)
);

AND2x4_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

NOR2x1_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_30),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_31),
.Y(n_33)
);

NOR3xp33_ASAP7_75t_SL g34 ( 
.A(n_33),
.B(n_28),
.C(n_32),
.Y(n_34)
);

NOR5xp2_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_23),
.C(n_4),
.D(n_30),
.E(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_34),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_30),
.B1(n_29),
.B2(n_35),
.Y(n_37)
);


endmodule