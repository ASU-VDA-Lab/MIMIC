module fake_jpeg_13010_n_298 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_219;
wire n_70;
wire n_102;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_56),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_46),
.B(n_72),
.Y(n_111)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_R g48 ( 
.A(n_25),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_73),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_50),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_53),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_17),
.Y(n_54)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_63),
.Y(n_99)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_19),
.B(n_1),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_65),
.Y(n_126)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_68),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_20),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_69),
.B(n_74),
.Y(n_95)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_20),
.B(n_15),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_21),
.B(n_1),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_21),
.B(n_4),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_76),
.B(n_79),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_27),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_73),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_78),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_23),
.B(n_4),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_23),
.B(n_4),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_26),
.B(n_8),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_86),
.Y(n_104)
);

NAND2x1_ASAP7_75t_SL g83 ( 
.A(n_22),
.B(n_28),
.Y(n_83)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_83),
.B(n_39),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_26),
.B(n_15),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_84),
.B(n_85),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_33),
.B(n_8),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_33),
.B(n_9),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_88),
.B(n_49),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_48),
.B1(n_66),
.B2(n_64),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_90),
.A2(n_108),
.B(n_123),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_46),
.A2(n_28),
.B(n_24),
.C(n_22),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_93),
.A2(n_113),
.B(n_9),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_38),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_97),
.B(n_119),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_45),
.A2(n_31),
.B1(n_36),
.B2(n_35),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_101),
.A2(n_35),
.B1(n_67),
.B2(n_77),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_107),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_31),
.C(n_36),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_55),
.B(n_24),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_34),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_51),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_62),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_71),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_127),
.Y(n_158)
);

NAND2x1_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_41),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_65),
.B(n_41),
.C(n_36),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_14),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_50),
.A2(n_41),
.B1(n_35),
.B2(n_38),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_114),
.B1(n_129),
.B2(n_94),
.Y(n_176)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_39),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_137),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_34),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_148),
.C(n_167),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_139),
.Y(n_206)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_141),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_89),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_144),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_143),
.A2(n_146),
.B1(n_159),
.B2(n_162),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_101),
.A2(n_82),
.B1(n_78),
.B2(n_71),
.Y(n_146)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

NAND2xp33_ASAP7_75t_SL g190 ( 
.A(n_150),
.B(n_174),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_88),
.B(n_10),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_161),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_107),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_156),
.Y(n_188)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_98),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_127),
.A2(n_82),
.B1(n_78),
.B2(n_51),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_11),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_98),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_163),
.B(n_173),
.Y(n_196)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_95),
.B(n_14),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_94),
.Y(n_169)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_92),
.B(n_118),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_172),
.B(n_175),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_99),
.B(n_105),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_96),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_114),
.B1(n_126),
.B2(n_129),
.Y(n_181)
);

NOR3xp33_ASAP7_75t_SL g177 ( 
.A(n_137),
.B(n_152),
.C(n_136),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_SL g215 ( 
.A(n_177),
.B(n_123),
.C(n_132),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_181),
.A2(n_204),
.B1(n_207),
.B2(n_91),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_120),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_193),
.B(n_183),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_175),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_200),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_133),
.B1(n_108),
.B2(n_90),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_199),
.A2(n_116),
.B1(n_145),
.B2(n_91),
.Y(n_220)
);

NAND3xp33_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_104),
.C(n_132),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_161),
.B(n_106),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_201),
.B(n_157),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_147),
.A2(n_90),
.B1(n_124),
.B2(n_116),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_147),
.A2(n_158),
.B1(n_150),
.B2(n_176),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_146),
.B1(n_165),
.B2(n_168),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_208),
.A2(n_218),
.B1(n_185),
.B2(n_189),
.Y(n_243)
);

AND2x6_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_165),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_212),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_154),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_224),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_211),
.B(n_219),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_160),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_220),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_190),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_222),
.C(n_223),
.Y(n_233)
);

NOR4xp25_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_187),
.C(n_87),
.D(n_112),
.Y(n_239)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

CKINVDCx12_ASAP7_75t_R g221 ( 
.A(n_179),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_221),
.B(n_228),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_174),
.C(n_155),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_112),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_112),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_140),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_229),
.Y(n_244)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_230),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_186),
.B(n_140),
.C(n_164),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_185),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_196),
.B(n_117),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_198),
.A2(n_169),
.B1(n_149),
.B2(n_141),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_224),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_218),
.A2(n_198),
.B1(n_178),
.B2(n_192),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_235),
.B1(n_243),
.B2(n_248),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_210),
.A2(n_178),
.B1(n_192),
.B2(n_191),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_182),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_237),
.B(n_241),
.Y(n_251)
);

AOI221xp5_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_209),
.B1(n_229),
.B2(n_205),
.C(n_87),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_182),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_213),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_212),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_210),
.A2(n_195),
.B1(n_205),
.B2(n_189),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_252),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_245),
.B(n_246),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_258),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_216),
.B1(n_225),
.B2(n_215),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_254),
.Y(n_271)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_260),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_220),
.B(n_222),
.Y(n_256)
);

A2O1A1O1Ixp25_ASAP7_75t_L g270 ( 
.A1(n_256),
.A2(n_244),
.B(n_231),
.C(n_234),
.D(n_232),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_238),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_233),
.Y(n_267)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_227),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_262),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_269),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_233),
.C(n_241),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_251),
.C(n_231),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_251),
.B(n_237),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_270),
.A2(n_256),
.B1(n_261),
.B2(n_257),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_276),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_280),
.C(n_269),
.Y(n_282)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_257),
.A3(n_248),
.B1(n_255),
.B2(n_250),
.C1(n_203),
.C2(n_195),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_272),
.B(n_202),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_278),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_264),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_271),
.A2(n_202),
.B1(n_203),
.B2(n_206),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_170),
.B1(n_102),
.B2(n_103),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_206),
.C(n_139),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_278),
.A2(n_270),
.B1(n_266),
.B2(n_268),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_282),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_279),
.A2(n_266),
.B(n_171),
.Y(n_284)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_284),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_286),
.A2(n_102),
.B1(n_117),
.B2(n_179),
.Y(n_289)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_285),
.A2(n_280),
.B(n_274),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_282),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_289),
.A2(n_284),
.B1(n_286),
.B2(n_281),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_291),
.A2(n_290),
.B1(n_285),
.B2(n_288),
.Y(n_294)
);

AO21x1_ASAP7_75t_L g295 ( 
.A1(n_292),
.A2(n_293),
.B(n_275),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_283),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_294),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_293),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_295),
.B(n_275),
.Y(n_298)
);


endmodule