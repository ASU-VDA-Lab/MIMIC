module fake_aes_10889_n_45 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_45);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_2), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_1), .B(n_4), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_11), .Y(n_19) );
BUFx6f_ASAP7_75t_L g20 ( .A(n_6), .Y(n_20) );
NAND2xp5_ASAP7_75t_SL g21 ( .A(n_2), .B(n_9), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_14), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_1), .B(n_10), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_18), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_16), .B(n_0), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_18), .A2(n_0), .B1(n_3), .B2(n_4), .Y(n_26) );
OAI22xp5_ASAP7_75t_L g27 ( .A1(n_18), .A2(n_3), .B1(n_5), .B2(n_7), .Y(n_27) );
OAI21x1_ASAP7_75t_L g28 ( .A1(n_24), .A2(n_17), .B(n_19), .Y(n_28) );
AO31x2_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_22), .A3(n_17), .B(n_16), .Y(n_29) );
INVx1_ASAP7_75t_SL g30 ( .A(n_28), .Y(n_30) );
OAI221xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_26), .B1(n_25), .B2(n_21), .C(n_23), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_29), .Y(n_32) );
INVx3_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
INVx1_ASAP7_75t_SL g35 ( .A(n_32), .Y(n_35) );
NAND3xp33_ASAP7_75t_L g36 ( .A(n_34), .B(n_33), .C(n_26), .Y(n_36) );
NAND4xp75_ASAP7_75t_SL g37 ( .A(n_35), .B(n_29), .C(n_33), .D(n_21), .Y(n_37) );
AOI21xp5_ASAP7_75t_L g38 ( .A1(n_34), .A2(n_33), .B(n_20), .Y(n_38) );
NOR4xp75_ASAP7_75t_SL g39 ( .A(n_37), .B(n_29), .C(n_12), .D(n_13), .Y(n_39) );
NOR2x1_ASAP7_75t_L g40 ( .A(n_36), .B(n_20), .Y(n_40) );
HB1xp67_ASAP7_75t_L g41 ( .A(n_38), .Y(n_41) );
AOI21xp5_ASAP7_75t_L g42 ( .A1(n_40), .A2(n_20), .B(n_8), .Y(n_42) );
NOR3xp33_ASAP7_75t_SL g43 ( .A(n_39), .B(n_20), .C(n_41), .Y(n_43) );
XNOR2xp5_ASAP7_75t_L g44 ( .A(n_43), .B(n_42), .Y(n_44) );
INVx1_ASAP7_75t_L g45 ( .A(n_44), .Y(n_45) );
endmodule