module fake_jpeg_22441_n_119 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_119);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_26),
.B1(n_23),
.B2(n_22),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_25),
.B1(n_24),
.B2(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_50),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_28),
.B1(n_25),
.B2(n_24),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_21),
.B(n_20),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_53),
.Y(n_54)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_18),
.Y(n_50)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_23),
.Y(n_51)
);

OA21x2_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_22),
.B(n_16),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_33),
.B(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_70),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_37),
.B1(n_29),
.B2(n_20),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_63),
.A2(n_46),
.B1(n_40),
.B2(n_52),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_66),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_17),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_17),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_18),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_54),
.B(n_41),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_0),
.B(n_1),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_56),
.C(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_40),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_83),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_61),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_1),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_89),
.B(n_90),
.Y(n_99)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_66),
.B(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_85),
.B(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_58),
.B(n_65),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_74),
.B(n_84),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_80),
.C(n_85),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_86),
.C(n_87),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_77),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_104),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_73),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_18),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_102),
.Y(n_107)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_110),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_88),
.B1(n_90),
.B2(n_92),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_111),
.Y(n_113)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

AOI321xp33_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_99),
.A3(n_97),
.B1(n_96),
.B2(n_98),
.C(n_104),
.Y(n_112)
);

OAI21x1_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_107),
.B(n_3),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_113),
.A2(n_114),
.B1(n_107),
.B2(n_7),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_9),
.Y(n_117)
);

AOI322xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_2),
.A3(n_10),
.B1(n_11),
.B2(n_115),
.C1(n_108),
.C2(n_73),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_11),
.Y(n_119)
);


endmodule