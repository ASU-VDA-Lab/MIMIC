module fake_jpeg_21951_n_289 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_289);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_27),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_19),
.B1(n_35),
.B2(n_21),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_37),
.B1(n_18),
.B2(n_30),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_49),
.A2(n_83),
.B1(n_34),
.B2(n_26),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_50),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_31),
.B1(n_20),
.B2(n_28),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_51),
.A2(n_52),
.B1(n_69),
.B2(n_7),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_31),
.B1(n_28),
.B2(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_53),
.B(n_61),
.Y(n_118)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_30),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_33),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_77),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_33),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_67),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_32),
.B1(n_28),
.B2(n_18),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_68),
.A2(n_75),
.B1(n_87),
.B2(n_34),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_28),
.B1(n_35),
.B2(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_33),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_70),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_28),
.C(n_22),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_19),
.B1(n_22),
.B2(n_29),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_29),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_76),
.Y(n_110)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_86),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_43),
.B(n_27),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_80),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_23),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_81),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_43),
.A2(n_23),
.B1(n_36),
.B2(n_26),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_36),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_1),
.Y(n_96)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_41),
.A2(n_26),
.B1(n_25),
.B2(n_34),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_92),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_93),
.B1(n_66),
.B2(n_62),
.Y(n_138)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_94),
.B(n_98),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_9),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_101),
.Y(n_135)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_3),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_68),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_87),
.B1(n_78),
.B2(n_64),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_4),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_108),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_120),
.B1(n_103),
.B2(n_96),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_6),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_56),
.B(n_7),
.Y(n_115)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_11),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_58),
.B(n_86),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_121),
.A2(n_125),
.B(n_111),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_122),
.B(n_129),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_123),
.A2(n_128),
.B1(n_138),
.B2(n_109),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_117),
.A2(n_93),
.B1(n_108),
.B2(n_105),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_124),
.A2(n_132),
.B1(n_136),
.B2(n_146),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_110),
.A2(n_58),
.B(n_65),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_74),
.C(n_59),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_148),
.C(n_119),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_133),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_95),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_137),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_64),
.B1(n_77),
.B2(n_54),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_112),
.Y(n_133)
);

NAND3xp33_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_9),
.C(n_10),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_SL g163 ( 
.A(n_134),
.B(n_14),
.C(n_16),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_88),
.B1(n_91),
.B2(n_101),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_10),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_151),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_88),
.A2(n_62),
.B1(n_74),
.B2(n_72),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_143),
.B1(n_104),
.B2(n_100),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_72),
.B1(n_59),
.B2(n_82),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_149),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_56),
.B1(n_57),
.B2(n_13),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_12),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_119),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_104),
.B1(n_17),
.B2(n_16),
.Y(n_178)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_162),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_156),
.C(n_141),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_118),
.C(n_89),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_159),
.B(n_161),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_164),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_102),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_165),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_102),
.Y(n_166)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

FAx1_ASAP7_75t_SL g167 ( 
.A(n_124),
.B(n_90),
.CI(n_92),
.CON(n_167),
.SN(n_167)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_167),
.B(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_170),
.Y(n_206)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_136),
.B(n_16),
.CI(n_17),
.CON(n_171),
.SN(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_172),
.Y(n_204)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_145),
.Y(n_180)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_199),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_125),
.B1(n_123),
.B2(n_146),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_190),
.A2(n_194),
.B1(n_196),
.B2(n_165),
.Y(n_211)
);

AND2x4_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_151),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_191),
.A2(n_195),
.B(n_168),
.Y(n_224)
);

A2O1A1O1Ixp25_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_122),
.B(n_139),
.C(n_151),
.D(n_141),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_193),
.B(n_181),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_157),
.A2(n_144),
.B1(n_131),
.B2(n_149),
.Y(n_194)
);

NAND2xp33_ASAP7_75t_SL g195 ( 
.A(n_164),
.B(n_167),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_157),
.A2(n_170),
.B1(n_169),
.B2(n_180),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_198),
.B(n_202),
.Y(n_222)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_209),
.B(n_212),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_187),
.A2(n_178),
.B1(n_159),
.B2(n_182),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_211),
.B1(n_215),
.B2(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_154),
.Y(n_213)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_171),
.B1(n_173),
.B2(n_155),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_171),
.B1(n_156),
.B2(n_168),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_216),
.A2(n_225),
.B1(n_197),
.B2(n_201),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_191),
.A2(n_181),
.B(n_163),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_218),
.A2(n_205),
.B1(n_189),
.B2(n_193),
.Y(n_241)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_219),
.Y(n_231)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_181),
.B(n_131),
.Y(n_221)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_224),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_201),
.A2(n_191),
.B1(n_192),
.B2(n_200),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_172),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_226),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_186),
.B(n_122),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_139),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_185),
.C(n_186),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_213),
.C(n_223),
.Y(n_247)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_235),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_216),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_219),
.A2(n_189),
.B1(n_198),
.B2(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_222),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_238),
.B(n_212),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_243),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_257),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_248),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_240),
.C(n_229),
.Y(n_258)
);

AOI31xp67_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_225),
.A3(n_221),
.B(n_224),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_227),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_251),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_233),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_250),
.A2(n_254),
.B(n_256),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_211),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_237),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_230),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_221),
.B(n_214),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_234),
.A2(n_218),
.B(n_220),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_209),
.B(n_204),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_258),
.A2(n_264),
.B(n_267),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_236),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g269 ( 
.A(n_263),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_255),
.A2(n_244),
.B1(n_250),
.B2(n_230),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_239),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_229),
.C(n_256),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_241),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_268),
.Y(n_275)
);

AOI21x1_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_251),
.B(n_253),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_272),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_266),
.C(n_258),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_242),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_262),
.B(n_245),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_273),
.A2(n_267),
.B(n_232),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_278),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_261),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_249),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_281),
.A2(n_282),
.B(n_279),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_277),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_275),
.B(n_232),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_283),
.B(n_282),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_284),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_280),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_286),
.B(n_285),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_269),
.Y(n_289)
);


endmodule