module fake_jpeg_9075_n_313 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_6),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_26),
.Y(n_53)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_17),
.B1(n_33),
.B2(n_29),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_45),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_17),
.B1(n_33),
.B2(n_31),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_46),
.A2(n_56),
.B1(n_57),
.B2(n_61),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_17),
.B1(n_31),
.B2(n_29),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_31),
.B1(n_23),
.B2(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_65),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_23),
.B1(n_22),
.B2(n_18),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_32),
.C(n_23),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_63),
.C(n_27),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_22),
.B1(n_30),
.B2(n_34),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_27),
.B1(n_34),
.B2(n_19),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_64),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_42),
.B(n_25),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_25),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_39),
.A2(n_21),
.B1(n_24),
.B2(n_30),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_57),
.B1(n_21),
.B2(n_24),
.Y(n_71)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_44),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_0),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_68),
.A2(n_78),
.B(n_81),
.Y(n_111)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_71),
.A2(n_95),
.B1(n_24),
.B2(n_21),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_76),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_28),
.Y(n_73)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_75),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_28),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_32),
.B(n_39),
.C(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_77),
.B(n_84),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_64),
.B(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_47),
.B(n_40),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_47),
.B(n_65),
.Y(n_80)
);

AOI32xp33_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_43),
.A3(n_40),
.B1(n_41),
.B2(n_39),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_83),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_50),
.Y(n_83)
);

CKINVDCx6p67_ASAP7_75t_R g85 ( 
.A(n_59),
.Y(n_85)
);

CKINVDCx10_ASAP7_75t_R g128 ( 
.A(n_85),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_90),
.Y(n_122)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_19),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_52),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_92),
.B(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_98),
.Y(n_125)
);

NOR2x1_ASAP7_75t_R g95 ( 
.A(n_45),
.B(n_43),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_18),
.Y(n_96)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_99),
.A2(n_104),
.B1(n_74),
.B2(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_58),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_35),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_102),
.Y(n_124)
);

OR2x2_ASAP7_75t_SL g103 ( 
.A(n_49),
.B(n_43),
.Y(n_103)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_60),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_105),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_123),
.B1(n_88),
.B2(n_74),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_121),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_10),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_118),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_43),
.B1(n_41),
.B2(n_44),
.Y(n_123)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_131),
.A2(n_87),
.B1(n_69),
.B2(n_98),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_93),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_141),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_84),
.Y(n_135)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_93),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_41),
.C(n_42),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_96),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_138),
.B(n_144),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_95),
.B(n_80),
.C(n_86),
.Y(n_139)
);

A2O1A1O1Ixp25_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_118),
.B(n_123),
.C(n_126),
.D(n_115),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_92),
.B(n_68),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_140),
.A2(n_150),
.B(n_162),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_68),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_105),
.B1(n_131),
.B2(n_113),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_81),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_89),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_94),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_127),
.B(n_77),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_146),
.B(n_148),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_125),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_153),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_102),
.Y(n_148)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_101),
.B(n_103),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_164),
.B(n_162),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_130),
.A2(n_79),
.B(n_71),
.C(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_151),
.B(n_155),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_125),
.B(n_100),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_119),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_114),
.B(n_104),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_159),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_132),
.B(n_91),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_158),
.B(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_71),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_161),
.Y(n_193)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_114),
.A2(n_71),
.B(n_42),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_42),
.B(n_44),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_166),
.A2(n_190),
.B(n_146),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_169),
.A2(n_180),
.B1(n_185),
.B2(n_154),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_126),
.Y(n_171)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_171),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_153),
.Y(n_172)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_108),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_175),
.C(n_184),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_108),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_177),
.B(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_115),
.B1(n_119),
.B2(n_112),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_181),
.B(n_196),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_110),
.Y(n_182)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_110),
.Y(n_183)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_152),
.A2(n_41),
.B1(n_8),
.B2(n_2),
.Y(n_185)
);

NOR3xp33_ASAP7_75t_SL g186 ( 
.A(n_137),
.B(n_42),
.C(n_44),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_160),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_42),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_184),
.C(n_190),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_192),
.B(n_150),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_42),
.Y(n_194)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_151),
.B(n_44),
.Y(n_195)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_163),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_158),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_199),
.C(n_204),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_181),
.A2(n_137),
.B1(n_149),
.B2(n_142),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_198),
.A2(n_178),
.B1(n_166),
.B2(n_175),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_141),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_211),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_173),
.A2(n_139),
.B1(n_149),
.B2(n_150),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_183),
.B1(n_173),
.B2(n_222),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_209),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_210),
.B(n_212),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_149),
.C(n_161),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_193),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_214),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_150),
.C(n_163),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

XOR2x2_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_176),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_150),
.C(n_44),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_220),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_44),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_207),
.B(n_189),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_223),
.B(n_225),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_217),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_215),
.B(n_179),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_202),
.A2(n_221),
.B1(n_203),
.B2(n_205),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_236),
.B1(n_241),
.B2(n_208),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_232),
.B(n_11),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_170),
.B(n_186),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_233),
.A2(n_242),
.B(n_244),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_234),
.A2(n_237),
.B1(n_10),
.B2(n_5),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_211),
.A2(n_170),
.B1(n_171),
.B2(n_165),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_198),
.A2(n_191),
.B1(n_165),
.B2(n_168),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_172),
.B1(n_168),
.B2(n_0),
.Y(n_238)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_200),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_204),
.A2(n_1),
.B(n_3),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_201),
.C(n_199),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_250),
.C(n_253),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_201),
.C(n_219),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_252),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_197),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_208),
.C(n_216),
.Y(n_253)
);

AOI321xp33_ASAP7_75t_L g254 ( 
.A1(n_232),
.A2(n_218),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_255),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_10),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_256),
.B(n_261),
.Y(n_271)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_259),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g258 ( 
.A(n_229),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_241),
.C(n_238),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_231),
.A2(n_234),
.B1(n_237),
.B2(n_229),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_275),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_227),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_271),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_251),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_245),
.A2(n_233),
.B1(n_242),
.B2(n_240),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_272),
.B(n_274),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_240),
.B(n_243),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_273),
.A2(n_254),
.B(n_260),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_238),
.B1(n_236),
.B2(n_244),
.Y(n_274)
);

NOR3xp33_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_238),
.C(n_6),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_277),
.B(n_283),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_252),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_270),
.Y(n_289)
);

NAND2xp33_ASAP7_75t_SL g294 ( 
.A(n_279),
.B(n_283),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_268),
.B(n_276),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_280),
.A2(n_286),
.B(n_279),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_282),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_246),
.C(n_250),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_255),
.C(n_266),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_284),
.B(n_285),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_11),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_11),
.C(n_7),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_14),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_291),
.C(n_15),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_288),
.A2(n_275),
.B1(n_1),
.B2(n_9),
.Y(n_290)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_294),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_8),
.B1(n_9),
.B2(n_13),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_296),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_14),
.Y(n_298)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_278),
.Y(n_299)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_304),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_292),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_294),
.B(n_295),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_300),
.C(n_302),
.Y(n_309)
);

AO21x1_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_310),
.B(n_308),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_306),
.B(n_301),
.Y(n_310)
);

OAI221xp5_ASAP7_75t_SL g312 ( 
.A1(n_311),
.A2(n_307),
.B1(n_289),
.B2(n_16),
.C(n_15),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_16),
.Y(n_313)
);


endmodule