module fake_jpeg_4571_n_99 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_31),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_61),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_0),
.Y(n_63)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_50),
.B1(n_55),
.B2(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_0),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_49),
.B1(n_43),
.B2(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_42),
.Y(n_75)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_69),
.B1(n_44),
.B2(n_58),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

OR2x2_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_1),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_59),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_2),
.B(n_3),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_83),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_80),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_76),
.A2(n_54),
.B1(n_51),
.B2(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_75),
.B(n_1),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_82),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_56),
.B1(n_53),
.B2(n_4),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_86),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_89),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_90),
.B(n_87),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_91),
.A2(n_85),
.B1(n_10),
.B2(n_15),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_9),
.C(n_16),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_19),
.B(n_21),
.C(n_23),
.Y(n_94)
);

NOR2xp67_ASAP7_75t_SL g95 ( 
.A(n_94),
.B(n_25),
.Y(n_95)
);

AOI221xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.C(n_32),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_37),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_38),
.Y(n_99)
);


endmodule