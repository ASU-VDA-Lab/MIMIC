module fake_jpeg_30357_n_141 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_19),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_23),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_35),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_66),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_47),
.C(n_53),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_76),
.Y(n_86)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_67),
.Y(n_74)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_61),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_88),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_78),
.B(n_47),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_72),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_93),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_66),
.C(n_59),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_5),
.B(n_6),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_74),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_50),
.C(n_59),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_3),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_68),
.B1(n_51),
.B2(n_58),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_92),
.B1(n_31),
.B2(n_9),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_52),
.B1(n_57),
.B2(n_49),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_2),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_3),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_97),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_107),
.B(n_15),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_26),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_102),
.C(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_4),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_56),
.B1(n_27),
.B2(n_30),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_22),
.B1(n_24),
.B2(n_32),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

AO22x1_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_106)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_7),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_113),
.B1(n_33),
.B2(n_34),
.Y(n_123)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_112),
.A2(n_83),
.B1(n_17),
.B2(n_18),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_8),
.B1(n_11),
.B2(n_13),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_121),
.Y(n_127)
);

NAND2x1_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_16),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_110),
.B(n_101),
.C(n_98),
.D(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_44),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_123),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_36),
.C(n_37),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_42),
.C(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_130),
.B1(n_124),
.B2(n_119),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_124),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_127),
.Y(n_132)
);

AOI321xp33_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_133),
.A3(n_114),
.B1(n_118),
.B2(n_129),
.C(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_132),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_134),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_138),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_129),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_114),
.Y(n_141)
);


endmodule