module fake_netlist_1_1278_n_684 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_684);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_684;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_621;
wire n_285;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_522;
wire n_264;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_49), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_5), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_59), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_73), .Y(n_81) );
INVxp33_ASAP7_75t_L g82 ( .A(n_37), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_27), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_39), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_41), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_65), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_25), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_8), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_30), .Y(n_89) );
BUFx2_ASAP7_75t_L g90 ( .A(n_14), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_66), .Y(n_91) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_54), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_1), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_29), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_7), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_28), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_15), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_24), .Y(n_98) );
INVxp67_ASAP7_75t_L g99 ( .A(n_23), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_13), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_50), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_76), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_21), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_63), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_72), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_57), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_22), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_32), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_35), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_64), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_4), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_13), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_3), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_77), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_43), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_19), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_34), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_14), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_61), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_62), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_20), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_67), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_70), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_11), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_1), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_83), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_83), .Y(n_127) );
INVx3_ASAP7_75t_L g128 ( .A(n_95), .Y(n_128) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_85), .A2(n_38), .B(n_74), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_85), .Y(n_130) );
XOR2xp5_ASAP7_75t_L g131 ( .A(n_93), .B(n_0), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_92), .B(n_0), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_89), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g136 ( .A1(n_93), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_89), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_91), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_91), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_106), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_106), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_95), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_78), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_80), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_81), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_96), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_102), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_103), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_104), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_105), .Y(n_150) );
INVxp67_ASAP7_75t_L g151 ( .A(n_90), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_109), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_88), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_110), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_115), .Y(n_155) );
BUFx2_ASAP7_75t_L g156 ( .A(n_90), .Y(n_156) );
AND2x6_ASAP7_75t_L g157 ( .A(n_116), .B(n_40), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_88), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_117), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_118), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_119), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_120), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_122), .Y(n_163) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_118), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_123), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_124), .Y(n_166) );
INVxp67_ASAP7_75t_L g167 ( .A(n_79), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_124), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_153), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_127), .A2(n_97), .B1(n_113), .B2(n_112), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_151), .B(n_82), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_156), .B(n_99), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_156), .B(n_121), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_127), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_160), .B(n_94), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_160), .B(n_94), .Y(n_177) );
INVx2_ASAP7_75t_SL g178 ( .A(n_164), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_143), .B(n_98), .Y(n_180) );
NOR3xp33_ASAP7_75t_L g181 ( .A(n_133), .B(n_125), .C(n_100), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_167), .B(n_111), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_129), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_144), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_144), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_153), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_126), .B(n_98), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_143), .B(n_145), .Y(n_188) );
OAI221xp5_ASAP7_75t_L g189 ( .A1(n_166), .A2(n_107), .B1(n_101), .B2(n_87), .C(n_108), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_145), .B(n_108), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_126), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_158), .Y(n_192) );
INVxp67_ASAP7_75t_L g193 ( .A(n_131), .Y(n_193) );
NOR3xp33_ASAP7_75t_L g194 ( .A(n_136), .B(n_114), .C(n_84), .Y(n_194) );
INVxp67_ASAP7_75t_L g195 ( .A(n_131), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_135), .B(n_114), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_135), .B(n_84), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_158), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_147), .B(n_42), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_147), .B(n_2), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_137), .B(n_44), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_137), .B(n_36), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_149), .B(n_5), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_141), .B(n_45), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_149), .B(n_46), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_158), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_154), .B(n_6), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_144), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_166), .B(n_6), .Y(n_209) );
O2A1O1Ixp5_ASAP7_75t_L g210 ( .A1(n_154), .A2(n_47), .B(n_71), .C(n_69), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_159), .B(n_7), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_158), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_141), .Y(n_213) );
AND2x6_ASAP7_75t_SL g214 ( .A(n_136), .B(n_8), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_159), .B(n_9), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_168), .B(n_9), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_168), .B(n_10), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_165), .B(n_10), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_157), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_165), .B(n_11), .Y(n_220) );
BUFx8_ASAP7_75t_L g221 ( .A(n_157), .Y(n_221) );
INVxp33_ASAP7_75t_L g222 ( .A(n_146), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_144), .B(n_51), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_130), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_146), .B(n_12), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_129), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_130), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_132), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_132), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_144), .B(n_48), .Y(n_230) );
NOR2xp33_ASAP7_75t_SL g231 ( .A(n_221), .B(n_157), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_169), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_213), .A2(n_157), .B1(n_148), .B2(n_161), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_175), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_216), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_179), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_222), .B(n_163), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_186), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_192), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_191), .B(n_163), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_181), .B(n_148), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_178), .A2(n_157), .B1(n_161), .B2(n_152), .Y(n_242) );
BUFx2_ASAP7_75t_L g243 ( .A(n_178), .Y(n_243) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_190), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_182), .B(n_152), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_171), .B(n_155), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_188), .A2(n_155), .B(n_134), .C(n_140), .Y(n_247) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_176), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_216), .A2(n_157), .B1(n_140), .B2(n_134), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_222), .B(n_139), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_224), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_180), .B(n_139), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_196), .Y(n_253) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_177), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_221), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_183), .Y(n_256) );
INVx3_ASAP7_75t_L g257 ( .A(n_227), .Y(n_257) );
BUFx4f_ASAP7_75t_L g258 ( .A(n_209), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_172), .A2(n_157), .B1(n_138), .B2(n_150), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_174), .B(n_138), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_174), .B(n_173), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_228), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_198), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_206), .Y(n_264) );
OAI22xp33_ASAP7_75t_L g265 ( .A1(n_189), .A2(n_142), .B1(n_128), .B2(n_162), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_212), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_184), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_193), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_221), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_229), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_217), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_196), .B(n_142), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_182), .B(n_142), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_187), .B(n_142), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_183), .Y(n_275) );
INVxp67_ASAP7_75t_SL g276 ( .A(n_200), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_225), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_187), .B(n_128), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_197), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_195), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_203), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_219), .B(n_150), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_207), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_211), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_184), .Y(n_285) );
INVx4_ASAP7_75t_L g286 ( .A(n_183), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_197), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_183), .A2(n_162), .B(n_150), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_170), .B(n_128), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_215), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_218), .B(n_128), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_185), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_226), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_220), .B(n_162), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_250), .B(n_194), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_258), .A2(n_226), .B1(n_199), .B2(n_205), .Y(n_296) );
AND2x6_ASAP7_75t_L g297 ( .A(n_255), .B(n_226), .Y(n_297) );
BUFx12f_ASAP7_75t_L g298 ( .A(n_268), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_250), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_237), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_243), .B(n_214), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_237), .B(n_226), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_273), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_243), .B(n_150), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_244), .B(n_150), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_248), .B(n_204), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_286), .Y(n_307) );
INVx5_ASAP7_75t_L g308 ( .A(n_255), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_235), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_265), .A2(n_204), .B(n_201), .C(n_202), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_257), .Y(n_311) );
INVx2_ASAP7_75t_SL g312 ( .A(n_258), .Y(n_312) );
NAND3xp33_ASAP7_75t_L g313 ( .A(n_233), .B(n_210), .C(n_202), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_256), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_269), .B(n_162), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_268), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_286), .Y(n_317) );
OAI31xp33_ASAP7_75t_L g318 ( .A1(n_254), .A2(n_230), .A3(n_223), .B(n_208), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_258), .A2(n_208), .B1(n_185), .B2(n_230), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_286), .Y(n_320) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_257), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_269), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_279), .B(n_12), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_280), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_245), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_246), .B(n_15), .Y(n_326) );
INVx5_ASAP7_75t_L g327 ( .A(n_257), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_245), .B(n_16), .Y(n_328) );
AOI21xp33_ASAP7_75t_SL g329 ( .A1(n_280), .A2(n_17), .B(n_18), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_245), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_281), .A2(n_283), .B(n_231), .Y(n_331) );
INVx3_ASAP7_75t_L g332 ( .A(n_262), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_232), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_262), .Y(n_334) );
INVx3_ASAP7_75t_SL g335 ( .A(n_274), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_281), .A2(n_26), .B(n_31), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_283), .A2(n_33), .B(n_52), .Y(n_337) );
INVx2_ASAP7_75t_SL g338 ( .A(n_272), .Y(n_338) );
INVx4_ASAP7_75t_L g339 ( .A(n_262), .Y(n_339) );
BUFx4_ASAP7_75t_SL g340 ( .A(n_253), .Y(n_340) );
OR2x6_ASAP7_75t_SL g341 ( .A(n_253), .B(n_53), .Y(n_341) );
NOR2xp67_ASAP7_75t_SL g342 ( .A(n_256), .B(n_55), .Y(n_342) );
OR2x6_ASAP7_75t_L g343 ( .A(n_287), .B(n_56), .Y(n_343) );
BUFx12f_ASAP7_75t_L g344 ( .A(n_272), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_333), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_333), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_321), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_303), .B(n_290), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_321), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_314), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_311), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_299), .B(n_284), .Y(n_352) );
OA21x2_ASAP7_75t_L g353 ( .A1(n_313), .A2(n_288), .B(n_247), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_311), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_339), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_300), .B(n_277), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_339), .Y(n_357) );
OA21x2_ASAP7_75t_L g358 ( .A1(n_331), .A2(n_337), .B(n_336), .Y(n_358) );
INVxp33_ASAP7_75t_L g359 ( .A(n_324), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_302), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_309), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_327), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_295), .B(n_277), .Y(n_363) );
INVx2_ASAP7_75t_SL g364 ( .A(n_327), .Y(n_364) );
XNOR2xp5_ASAP7_75t_L g365 ( .A(n_301), .B(n_241), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_327), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_332), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_344), .A2(n_241), .B1(n_274), .B2(n_289), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_314), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_338), .B(n_271), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_314), .Y(n_371) );
OAI22xp33_ASAP7_75t_L g372 ( .A1(n_341), .A2(n_271), .B1(n_270), .B2(n_252), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_325), .A2(n_274), .B1(n_241), .B2(n_270), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_332), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_334), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_334), .Y(n_376) );
BUFx12f_ASAP7_75t_L g377 ( .A(n_364), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_372), .B(n_330), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_348), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_348), .B(n_276), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_372), .A2(n_343), .B1(n_326), .B2(n_327), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_363), .B(n_323), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_355), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_345), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_345), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_346), .Y(n_386) );
INVx3_ASAP7_75t_L g387 ( .A(n_366), .Y(n_387) );
BUFx12f_ASAP7_75t_L g388 ( .A(n_364), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_352), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_346), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_352), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_356), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_363), .B(n_343), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_350), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_350), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_356), .B(n_343), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_361), .B(n_373), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_355), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_360), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_364), .B(n_320), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_361), .B(n_306), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_347), .B(n_335), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_350), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_350), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_394), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_384), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_394), .Y(n_407) );
OAI33xp33_ASAP7_75t_L g408 ( .A1(n_381), .A2(n_278), .A3(n_291), .B1(n_304), .B2(n_316), .B3(n_296), .Y(n_408) );
OAI211xp5_ASAP7_75t_L g409 ( .A1(n_381), .A2(n_368), .B(n_323), .C(n_316), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_384), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_385), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_379), .B(n_347), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_392), .B(n_349), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_389), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g415 ( .A1(n_382), .A2(n_365), .B1(n_373), .B2(n_261), .C(n_306), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_380), .B(n_370), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_393), .B(n_359), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_385), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_380), .B(n_370), .Y(n_419) );
OAI211xp5_ASAP7_75t_L g420 ( .A1(n_393), .A2(n_305), .B(n_329), .C(n_362), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_392), .B(n_349), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_398), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_386), .B(n_360), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_386), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_390), .B(n_351), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_390), .Y(n_426) );
NOR2x1_ASAP7_75t_L g427 ( .A(n_398), .B(n_366), .Y(n_427) );
OAI322xp33_ASAP7_75t_L g428 ( .A1(n_378), .A2(n_365), .A3(n_335), .B1(n_294), .B2(n_240), .C1(n_251), .C2(n_260), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_396), .A2(n_344), .B1(n_298), .B2(n_357), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_394), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_399), .Y(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_398), .B(n_366), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_395), .Y(n_433) );
BUFx2_ASAP7_75t_L g434 ( .A(n_383), .Y(n_434) );
BUFx3_ASAP7_75t_L g435 ( .A(n_377), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_391), .B(n_351), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_395), .Y(n_437) );
NAND4xp25_ASAP7_75t_L g438 ( .A(n_396), .B(n_249), .C(n_242), .D(n_322), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_399), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_377), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_406), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_406), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_415), .A2(n_397), .B1(n_378), .B2(n_401), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_414), .B(n_383), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_410), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_410), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_417), .B(n_402), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_423), .B(n_397), .Y(n_448) );
INVxp33_ASAP7_75t_L g449 ( .A(n_440), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_411), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_411), .Y(n_451) );
NAND4xp25_ASAP7_75t_SL g452 ( .A(n_429), .B(n_340), .C(n_298), .D(n_402), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_418), .Y(n_453) );
NOR2x1_ASAP7_75t_L g454 ( .A(n_435), .B(n_387), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_409), .B(n_420), .C(n_427), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_416), .B(n_377), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_419), .B(n_388), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_434), .B(n_387), .Y(n_458) );
OR2x6_ASAP7_75t_L g459 ( .A(n_435), .B(n_388), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_423), .B(n_401), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_418), .Y(n_461) );
OAI21xp33_ASAP7_75t_L g462 ( .A1(n_435), .A2(n_315), .B(n_400), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_424), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_436), .B(n_400), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_434), .B(n_387), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_424), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_428), .B(n_388), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_426), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_431), .B(n_400), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_422), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_412), .B(n_362), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_412), .B(n_387), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_431), .B(n_404), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_426), .Y(n_474) );
INVx3_ASAP7_75t_L g475 ( .A(n_432), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_425), .B(n_354), .Y(n_476) );
BUFx2_ASAP7_75t_L g477 ( .A(n_432), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_439), .B(n_404), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_439), .B(n_404), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_425), .B(n_354), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_413), .B(n_374), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_413), .B(n_374), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_438), .A2(n_310), .B(n_328), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_421), .B(n_367), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_421), .B(n_357), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_427), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_405), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_405), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_405), .B(n_403), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_470), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_441), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_444), .B(n_437), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_448), .B(n_437), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_447), .B(n_432), .Y(n_494) );
NOR3xp33_ASAP7_75t_L g495 ( .A(n_452), .B(n_408), .C(n_366), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_471), .B(n_432), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_442), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_445), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_446), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_475), .B(n_437), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_464), .B(n_469), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_485), .B(n_433), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_469), .B(n_433), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_450), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_449), .B(n_322), .Y(n_505) );
INVxp67_ASAP7_75t_SL g506 ( .A(n_489), .Y(n_506) );
AND2x2_ASAP7_75t_SL g507 ( .A(n_467), .B(n_340), .Y(n_507) );
NAND2x1p5_ASAP7_75t_L g508 ( .A(n_454), .B(n_308), .Y(n_508) );
NOR2xp33_ASAP7_75t_SL g509 ( .A(n_455), .B(n_407), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_456), .B(n_430), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_477), .B(n_430), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_443), .A2(n_315), .B1(n_312), .B2(n_367), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_451), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_472), .B(n_430), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_476), .B(n_407), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_460), .B(n_407), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_458), .B(n_403), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_453), .Y(n_518) );
NOR2xp67_ASAP7_75t_SL g519 ( .A(n_459), .B(n_308), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_457), .B(n_403), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_461), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_463), .B(n_395), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_466), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_468), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_465), .B(n_353), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_473), .B(n_479), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_474), .Y(n_527) );
INVx1_ASAP7_75t_SL g528 ( .A(n_459), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_487), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_488), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_459), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_473), .B(n_353), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_475), .B(n_376), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_478), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_489), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_480), .B(n_308), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_486), .B(n_358), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_484), .B(n_358), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_481), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_482), .B(n_308), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_483), .B(n_358), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_462), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_483), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_447), .B(n_376), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_543), .B(n_358), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_530), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_509), .B(n_350), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_501), .B(n_358), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_506), .B(n_371), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_509), .B(n_350), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_535), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_539), .B(n_315), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_515), .B(n_375), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_494), .B(n_58), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_492), .B(n_371), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_534), .B(n_375), .Y(n_556) );
INVx3_ASAP7_75t_L g557 ( .A(n_500), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_491), .B(n_318), .Y(n_558) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_529), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_513), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_490), .B(n_371), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_497), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_498), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_490), .B(n_369), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_499), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_504), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_518), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_526), .B(n_369), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_510), .B(n_369), .Y(n_569) );
NOR2x1_ASAP7_75t_L g570 ( .A(n_528), .B(n_317), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_521), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_529), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_523), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_524), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_527), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_516), .B(n_297), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_542), .B(n_60), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_496), .B(n_68), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_531), .B(n_314), .Y(n_579) );
NOR2x1_ASAP7_75t_L g580 ( .A(n_531), .B(n_307), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_506), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_502), .B(n_297), .Y(n_582) );
CKINVDCx14_ASAP7_75t_R g583 ( .A(n_520), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_493), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_493), .B(n_297), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_544), .B(n_297), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_511), .B(n_75), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_503), .B(n_297), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_522), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_514), .B(n_259), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_537), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_522), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_525), .B(n_319), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_517), .Y(n_594) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_581), .B(n_495), .C(n_541), .Y(n_595) );
OAI21xp33_ASAP7_75t_L g596 ( .A1(n_583), .A2(n_541), .B(n_495), .Y(n_596) );
NOR3xp33_ASAP7_75t_SL g597 ( .A(n_577), .B(n_505), .C(n_545), .Y(n_597) );
AOI211xp5_ASAP7_75t_L g598 ( .A1(n_581), .A2(n_519), .B(n_536), .C(n_540), .Y(n_598) );
NAND3xp33_ASAP7_75t_L g599 ( .A(n_570), .B(n_537), .C(n_538), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_547), .A2(n_538), .B(n_532), .Y(n_600) );
NOR2xp33_ASAP7_75t_SL g601 ( .A(n_580), .B(n_507), .Y(n_601) );
NAND5xp2_ASAP7_75t_L g602 ( .A(n_577), .B(n_512), .C(n_508), .D(n_533), .E(n_532), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_547), .A2(n_508), .B(n_320), .Y(n_603) );
NOR3x1_ASAP7_75t_L g604 ( .A(n_583), .B(n_312), .C(n_282), .Y(n_604) );
AOI211xp5_ASAP7_75t_SL g605 ( .A1(n_559), .A2(n_317), .B(n_307), .C(n_263), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_584), .B(n_293), .Y(n_606) );
NOR2xp33_ASAP7_75t_SL g607 ( .A(n_554), .B(n_342), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_594), .B(n_293), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_562), .B(n_293), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_563), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_589), .B(n_293), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_592), .B(n_293), .Y(n_612) );
NAND4xp25_ASAP7_75t_L g613 ( .A(n_545), .B(n_548), .C(n_553), .D(n_578), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_559), .B(n_275), .Y(n_614) );
NOR2xp33_ASAP7_75t_SL g615 ( .A(n_587), .B(n_275), .Y(n_615) );
INVx2_ASAP7_75t_SL g616 ( .A(n_561), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_565), .Y(n_617) );
AOI211xp5_ASAP7_75t_L g618 ( .A1(n_550), .A2(n_275), .B(n_256), .C(n_236), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_566), .Y(n_619) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_579), .A2(n_232), .B(n_234), .Y(n_620) );
OAI21xp5_ASAP7_75t_L g621 ( .A1(n_579), .A2(n_234), .B(n_238), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_567), .Y(n_622) );
NOR3xp33_ASAP7_75t_L g623 ( .A(n_552), .B(n_238), .C(n_239), .Y(n_623) );
XNOR2x1_ASAP7_75t_L g624 ( .A(n_568), .B(n_239), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_572), .B(n_256), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_572), .B(n_256), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_557), .A2(n_275), .B1(n_266), .B2(n_264), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_591), .B(n_275), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_591), .B(n_264), .Y(n_629) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_616), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_610), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_617), .B(n_571), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_602), .A2(n_573), .B1(n_574), .B2(n_575), .Y(n_633) );
OAI21xp33_ASAP7_75t_L g634 ( .A1(n_596), .A2(n_557), .B(n_551), .Y(n_634) );
OAI21xp5_ASAP7_75t_L g635 ( .A1(n_605), .A2(n_550), .B(n_558), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_595), .A2(n_551), .B1(n_560), .B2(n_556), .C(n_546), .Y(n_636) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_623), .A2(n_593), .B(n_576), .C(n_564), .Y(n_637) );
XNOR2xp5_ASAP7_75t_L g638 ( .A(n_624), .B(n_586), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_619), .B(n_560), .Y(n_639) );
BUFx2_ASAP7_75t_L g640 ( .A(n_599), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_622), .B(n_546), .Y(n_641) );
INVxp33_ASAP7_75t_L g642 ( .A(n_601), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_613), .B(n_549), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_597), .A2(n_557), .B1(n_588), .B2(n_549), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_600), .B(n_555), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_629), .Y(n_646) );
OAI21xp5_ASAP7_75t_SL g647 ( .A1(n_623), .A2(n_582), .B(n_569), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_606), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g649 ( .A1(n_598), .A2(n_585), .B(n_590), .Y(n_649) );
XNOR2x1_ASAP7_75t_L g650 ( .A(n_608), .B(n_266), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_615), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_645), .B(n_600), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_651), .B(n_604), .Y(n_653) );
NOR4xp75_ASAP7_75t_SL g654 ( .A(n_643), .B(n_614), .C(n_612), .D(n_611), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_639), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_640), .B(n_609), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_630), .B(n_626), .Y(n_657) );
NOR2x1_ASAP7_75t_L g658 ( .A(n_635), .B(n_621), .Y(n_658) );
OAI211xp5_ASAP7_75t_L g659 ( .A1(n_633), .A2(n_618), .B(n_603), .C(n_620), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_642), .A2(n_603), .B1(n_627), .B2(n_625), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_630), .B(n_628), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_641), .B(n_648), .Y(n_662) );
NAND4xp25_ASAP7_75t_L g663 ( .A(n_633), .B(n_607), .C(n_285), .D(n_292), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_636), .B(n_267), .C(n_642), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_644), .B(n_631), .Y(n_665) );
INVx3_ASAP7_75t_L g666 ( .A(n_657), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_661), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_662), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_658), .A2(n_647), .B1(n_634), .B2(n_638), .Y(n_669) );
INVx3_ASAP7_75t_L g670 ( .A(n_653), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_652), .B(n_646), .Y(n_671) );
NAND3xp33_ASAP7_75t_L g672 ( .A(n_664), .B(n_650), .C(n_637), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_655), .Y(n_673) );
NAND3xp33_ASAP7_75t_L g674 ( .A(n_669), .B(n_656), .C(n_660), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_669), .A2(n_653), .B1(n_665), .B2(n_659), .Y(n_675) );
NOR3xp33_ASAP7_75t_L g676 ( .A(n_670), .B(n_672), .C(n_666), .Y(n_676) );
INVx2_ASAP7_75t_SL g677 ( .A(n_670), .Y(n_677) );
INVxp67_ASAP7_75t_L g678 ( .A(n_677), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_676), .B(n_668), .Y(n_679) );
INVx2_ASAP7_75t_SL g680 ( .A(n_674), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_680), .A2(n_675), .B1(n_666), .B2(n_671), .Y(n_681) );
AOI22x1_ASAP7_75t_L g682 ( .A1(n_678), .A2(n_673), .B1(n_667), .B2(n_654), .Y(n_682) );
OR2x6_ASAP7_75t_L g683 ( .A(n_681), .B(n_679), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_683), .A2(n_663), .B1(n_682), .B2(n_649), .C(n_632), .Y(n_684) );
endmodule