module fake_jpeg_26106_n_272 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_35),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_35),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_48),
.B1(n_53),
.B2(n_58),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_27),
.B1(n_23),
.B2(n_28),
.Y(n_48)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_27),
.B1(n_23),
.B2(n_29),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_57),
.B(n_32),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_29),
.B1(n_26),
.B2(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_65),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_25),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_38),
.Y(n_79)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_37),
.B(n_39),
.C(n_29),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_68),
.A2(n_99),
.B1(n_102),
.B2(n_36),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_51),
.B(n_38),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_79),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_24),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_71),
.B(n_78),
.Y(n_118)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_73),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_26),
.B1(n_32),
.B2(n_39),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_74),
.A2(n_90),
.B1(n_42),
.B2(n_1),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_82),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_47),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_77),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_47),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_87),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_56),
.B(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_51),
.B(n_34),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_19),
.B(n_21),
.Y(n_89)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_89),
.A2(n_18),
.B(n_42),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_50),
.A2(n_32),
.B1(n_40),
.B2(n_34),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_49),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_31),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_95),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_97),
.Y(n_129)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_38),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_54),
.A2(n_33),
.B1(n_20),
.B2(n_31),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_38),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_42),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_30),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_46),
.A2(n_33),
.B1(n_20),
.B2(n_30),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_40),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_42),
.B1(n_22),
.B2(n_18),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_22),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_36),
.B1(n_40),
.B2(n_42),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_117),
.B1(n_68),
.B2(n_70),
.Y(n_135)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_126),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_72),
.A2(n_21),
.B1(n_17),
.B2(n_22),
.Y(n_117)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_21),
.C(n_17),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_70),
.C(n_69),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_123),
.B(n_128),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_131),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

CKINVDCx12_ASAP7_75t_R g126 ( 
.A(n_92),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_89),
.B(n_100),
.Y(n_148)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_86),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_133),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_127),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_134),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_146),
.B1(n_139),
.B2(n_142),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_128),
.B1(n_111),
.B2(n_131),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_136),
.A2(n_125),
.B1(n_109),
.B2(n_130),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_123),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_150),
.Y(n_168)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_69),
.CI(n_83),
.CON(n_140),
.SN(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_159),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_104),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_141),
.A2(n_107),
.B(n_113),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_129),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_150),
.B(n_139),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_151),
.C(n_160),
.Y(n_172)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_104),
.C(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_153),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_81),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_108),
.A2(n_76),
.B1(n_88),
.B2(n_96),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_132),
.B1(n_116),
.B2(n_107),
.Y(n_179)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_87),
.Y(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_97),
.C(n_85),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_73),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_42),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_167),
.B1(n_181),
.B2(n_164),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_142),
.A2(n_130),
.B1(n_120),
.B2(n_109),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_163),
.A2(n_166),
.B(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_164),
.B(n_173),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_121),
.B(n_106),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_109),
.B1(n_112),
.B2(n_120),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_141),
.B(n_147),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_156),
.B(n_113),
.Y(n_173)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_176),
.B(n_137),
.CI(n_153),
.CON(n_198),
.SN(n_198)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_179),
.A2(n_183),
.B1(n_143),
.B2(n_144),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_134),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_182),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_77),
.B1(n_78),
.B2(n_84),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_132),
.B1(n_116),
.B2(n_84),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_85),
.Y(n_185)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_0),
.B(n_1),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_186),
.A2(n_75),
.B1(n_91),
.B2(n_2),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_163),
.B1(n_184),
.B2(n_183),
.Y(n_211)
);

XOR2x2_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_140),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_189),
.A2(n_203),
.B(n_207),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_149),
.C(n_145),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_195),
.C(n_204),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_160),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_198),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_138),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_197),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_137),
.C(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_205),
.B(n_170),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_141),
.Y(n_201)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_167),
.B1(n_181),
.B2(n_177),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_158),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_140),
.C(n_159),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_143),
.B(n_95),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_214),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_203),
.B(n_205),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_203),
.B1(n_189),
.B2(n_199),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_175),
.Y(n_212)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_223),
.B1(n_188),
.B2(n_201),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_166),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_218),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_178),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_177),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_224),
.C(n_191),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_187),
.A2(n_165),
.B1(n_180),
.B2(n_175),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_165),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_226),
.A2(n_230),
.B(n_232),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_214),
.B(n_173),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_236),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_231),
.B1(n_233),
.B2(n_235),
.Y(n_245)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_221),
.A2(n_219),
.B1(n_209),
.B2(n_218),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_210),
.B1(n_208),
.B2(n_182),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_234),
.B(n_215),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_198),
.B1(n_194),
.B2(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_198),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_238),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_207),
.B1(n_179),
.B2(n_16),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_220),
.C(n_224),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_247),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_244),
.Y(n_251)
);

OR2x2_ASAP7_75t_SL g243 ( 
.A(n_226),
.B(n_233),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_243),
.A2(n_248),
.B(n_1),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_16),
.C(n_73),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_231),
.B(n_0),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_254),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_242),
.A2(n_235),
.B1(n_225),
.B2(n_73),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_252),
.A2(n_245),
.B1(n_241),
.B2(n_240),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_253),
.A2(n_8),
.B(n_9),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_225),
.B1(n_3),
.B2(n_4),
.Y(n_254)
);

OAI221xp5_ASAP7_75t_SL g255 ( 
.A1(n_246),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_255)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_255),
.A2(n_6),
.B(n_7),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_256),
.B(n_259),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_5),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_258),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_5),
.C(n_6),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_260),
.A2(n_252),
.B1(n_10),
.B2(n_12),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_261),
.A2(n_254),
.B(n_10),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_263),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_265),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_268),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_264),
.A2(n_257),
.B(n_259),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_251),
.B(n_10),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_9),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_269),
.Y(n_272)
);


endmodule