module real_jpeg_19685_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_0),
.A2(n_5),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_0),
.A2(n_10),
.B1(n_33),
.B2(n_45),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_1),
.A2(n_5),
.B1(n_44),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_2),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_22),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_2),
.A2(n_3),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_2),
.A2(n_22),
.B(n_27),
.C(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_3),
.A2(n_6),
.B1(n_25),
.B2(n_27),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_3),
.A2(n_10),
.B1(n_27),
.B2(n_33),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_3),
.A2(n_5),
.B1(n_27),
.B2(n_44),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_SL g86 ( 
.A1(n_3),
.A2(n_6),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_3),
.B(n_114),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_3),
.A2(n_5),
.B(n_9),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_3),
.B(n_31),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_3),
.A2(n_7),
.B(n_25),
.C(n_145),
.Y(n_144)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_5),
.B(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_5),
.A2(n_9),
.B1(n_44),
.B2(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_6),
.A2(n_8),
.B1(n_22),
.B2(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_6),
.A2(n_7),
.B1(n_25),
.B2(n_32),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_7),
.A2(n_10),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_9),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_9),
.A2(n_10),
.B1(n_33),
.B2(n_52),
.Y(n_54)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_10),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_10),
.A2(n_27),
.B(n_52),
.C(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_91),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_89),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_74),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_14),
.B(n_74),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

BUFx24_ASAP7_75t_SL g177 ( 
.A(n_15),
.Y(n_177)
);

FAx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_57),
.CI(n_66),
.CON(n_15),
.SN(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_39),
.B2(n_56),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_17),
.A2(n_18),
.B1(n_68),
.B2(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_17),
.A2(n_18),
.B1(n_83),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_29),
.B1(n_37),
.B2(n_38),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_19),
.B(n_38),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_19),
.A2(n_38),
.B(n_72),
.C(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_19),
.A2(n_37),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_26),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_24),
.Y(n_20)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_24),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_27),
.B(n_51),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_27),
.B(n_46),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_27),
.A2(n_32),
.B(n_33),
.Y(n_145)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_29),
.B(n_37),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_29),
.A2(n_38),
.B1(n_49),
.B2(n_80),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_29),
.B(n_88),
.C(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_29),
.A2(n_38),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_36),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_35),
.Y(n_34)
);

AOI211xp5_ASAP7_75t_SL g96 ( 
.A1(n_37),
.A2(n_49),
.B(n_73),
.C(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_38),
.B(n_80),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_38),
.A2(n_80),
.B(n_147),
.C(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_49),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_40),
.A2(n_49),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_40),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_42),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_43),
.B1(n_46),
.B2(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_44),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_69),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_49),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_49),
.A2(n_69),
.B1(n_80),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_49),
.A2(n_80),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_49),
.A2(n_80),
.B1(n_122),
.B2(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_49),
.B(n_88),
.C(n_126),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_49),
.A2(n_80),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_49),
.B(n_153),
.C(n_159),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_55),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_51),
.B(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_53),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_62),
.B2(n_65),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_71),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_62),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B(n_72),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_69),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.C(n_81),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_75),
.A2(n_76),
.B1(n_78),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_78),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_80),
.B(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_81),
.A2(n_82),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_85),
.B1(n_88),
.B2(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_88),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_88),
.A2(n_110),
.B1(n_125),
.B2(n_128),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_88),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_88),
.B(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_88),
.A2(n_110),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_88),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_156)
);

NAND2x1_ASAP7_75t_SL g160 ( 
.A(n_88),
.B(n_144),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_115),
.B(n_170),
.C(n_176),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_103),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_93),
.B(n_103),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_101),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_95),
.B(n_99),
.C(n_101),
.Y(n_171)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_97),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.C(n_111),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_104),
.A2(n_105),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_106),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_106),
.A2(n_107),
.B1(n_143),
.B2(n_147),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_111),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_169),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_162),
.B(n_168),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_149),
.B(n_161),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_140),
.B(n_148),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_129),
.B(n_139),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_124),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_122),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_125),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_136),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_142),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_143),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_144),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_150),
.B(n_152),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_163),
.B(n_164),
.Y(n_168)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_171),
.B(n_172),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);


endmodule