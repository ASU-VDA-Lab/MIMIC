module fake_netlist_6_2204_n_786 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_786);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_786;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_148;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_772;
wire n_656;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_118),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_101),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_46),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_74),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_106),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_38),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_50),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_138),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_43),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_31),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_103),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_14),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_53),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_93),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_81),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_112),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_1),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_8),
.Y(n_171)
);

BUFx2_ASAP7_75t_SL g172 ( 
.A(n_132),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_147),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_24),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_30),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_10),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_45),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_122),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_60),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_35),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_141),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_107),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_40),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_41),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_17),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_58),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_19),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_95),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_44),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_71),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_26),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_142),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_8),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_3),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_126),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_85),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_49),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_97),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_127),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_76),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_161),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_173),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_171),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_0),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_163),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_196),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_150),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_151),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_156),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_153),
.B(n_0),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_152),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_164),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

INVxp33_ASAP7_75t_SL g221 ( 
.A(n_193),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_160),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_155),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_167),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_168),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_169),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_177),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_157),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_158),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_R g233 ( 
.A(n_178),
.B(n_32),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_180),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_181),
.Y(n_236)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_165),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_166),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g242 ( 
.A(n_200),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_184),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_185),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_183),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_188),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_182),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_204),
.Y(n_248)
);

OAI21x1_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_215),
.B(n_214),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_208),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_202),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_182),
.Y(n_252)
);

AND2x4_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_202),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_211),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_219),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_215),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_224),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_216),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_225),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_227),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_206),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_205),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_236),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_206),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_243),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_218),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_229),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_209),
.Y(n_271)
);

AND2x6_ASAP7_75t_L g272 ( 
.A(n_207),
.B(n_191),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_209),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_229),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_203),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_210),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_231),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_223),
.B(n_148),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_231),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_234),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_234),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_244),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_246),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_238),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_235),
.Y(n_286)
);

AND2x4_ASAP7_75t_L g287 ( 
.A(n_238),
.B(n_198),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_212),
.B(n_148),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_241),
.B(n_149),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_241),
.B(n_149),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_245),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_245),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_217),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_220),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_240),
.B(n_154),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_249),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_237),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_221),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_240),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_232),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_257),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_172),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_222),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_257),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_249),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_288),
.B(n_232),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_257),
.Y(n_307)
);

OAI21xp33_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_174),
.B(n_176),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_259),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_292),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_295),
.B(n_233),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_251),
.B(n_230),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_292),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_276),
.Y(n_315)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_292),
.Y(n_316)
);

AND2x6_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_33),
.Y(n_317)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_292),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_248),
.B(n_154),
.Y(n_320)
);

AO21x2_ASAP7_75t_L g321 ( 
.A1(n_247),
.A2(n_201),
.B(n_199),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_259),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_250),
.B(n_159),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_287),
.B(n_253),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_292),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_291),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_291),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_276),
.B(n_189),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_289),
.Y(n_330)
);

BUFx6f_ASAP7_75t_SL g331 ( 
.A(n_289),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_290),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_269),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_256),
.Y(n_334)
);

AO21x2_ASAP7_75t_L g335 ( 
.A1(n_247),
.A2(n_201),
.B(n_199),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_289),
.A2(n_194),
.B1(n_192),
.B2(n_190),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_272),
.A2(n_187),
.B1(n_194),
.B2(n_192),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_272),
.A2(n_197),
.B1(n_190),
.B2(n_159),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_269),
.Y(n_339)
);

BUFx4f_ASAP7_75t_L g340 ( 
.A(n_272),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_287),
.B(n_197),
.Y(n_341)
);

BUFx6f_ASAP7_75t_SL g342 ( 
.A(n_289),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_291),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_272),
.B(n_34),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_290),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_287),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_287),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_269),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_253),
.B(n_36),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_286),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_270),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_272),
.B(n_37),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_L g354 ( 
.A1(n_258),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_270),
.Y(n_355)
);

AND2x6_ASAP7_75t_L g356 ( 
.A(n_253),
.B(n_39),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_278),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_270),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_274),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_260),
.B(n_2),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_272),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_346),
.B(n_272),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_333),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_340),
.B(n_261),
.Y(n_364)
);

OR2x6_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_253),
.Y(n_365)
);

AND2x6_ASAP7_75t_SL g366 ( 
.A(n_298),
.B(n_252),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_263),
.Y(n_367)
);

AND2x6_ASAP7_75t_SL g368 ( 
.A(n_297),
.B(n_252),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_324),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_327),
.B(n_266),
.Y(n_370)
);

NAND3xp33_ASAP7_75t_L g371 ( 
.A(n_315),
.B(n_284),
.C(n_283),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_337),
.A2(n_268),
.B1(n_279),
.B2(n_278),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_329),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_327),
.B(n_274),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_317),
.A2(n_281),
.B1(n_280),
.B2(n_274),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

NAND3xp33_ASAP7_75t_SL g377 ( 
.A(n_337),
.B(n_273),
.C(n_264),
.Y(n_377)
);

INVx8_ASAP7_75t_L g378 ( 
.A(n_331),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_340),
.B(n_280),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_310),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_317),
.A2(n_281),
.B1(n_280),
.B2(n_285),
.Y(n_381)
);

OAI22xp33_ASAP7_75t_L g382 ( 
.A1(n_330),
.A2(n_285),
.B1(n_282),
.B2(n_271),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_327),
.B(n_281),
.Y(n_383)
);

OAI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_360),
.A2(n_282),
.B1(n_277),
.B2(n_275),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_357),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_333),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_357),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_317),
.A2(n_277),
.B1(n_275),
.B2(n_273),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_327),
.B(n_254),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_324),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_299),
.B(n_264),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_324),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_324),
.B(n_347),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_299),
.B(n_267),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_347),
.B(n_254),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g396 ( 
.A(n_300),
.B(n_267),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_328),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_340),
.B(n_271),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_310),
.A2(n_262),
.B1(n_255),
.B2(n_82),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_347),
.B(n_255),
.Y(n_400)
);

NOR2x1_ASAP7_75t_R g401 ( 
.A(n_334),
.B(n_262),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_313),
.B(n_42),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_347),
.B(n_47),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_329),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_347),
.B(n_48),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_300),
.Y(n_406)
);

NAND2xp33_ASAP7_75t_L g407 ( 
.A(n_317),
.B(n_51),
.Y(n_407)
);

NOR2x1p5_ASAP7_75t_L g408 ( 
.A(n_313),
.B(n_4),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_323),
.B(n_4),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_332),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_350),
.B(n_52),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_350),
.B(n_54),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_339),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_350),
.B(n_55),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_350),
.B(n_348),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_348),
.B(n_56),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_361),
.B(n_57),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_312),
.B(n_5),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_339),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_317),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_348),
.B(n_59),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_348),
.B(n_61),
.Y(n_422)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_356),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_361),
.B(n_63),
.Y(n_424)
);

NOR3xp33_ASAP7_75t_L g425 ( 
.A(n_306),
.B(n_320),
.C(n_354),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_308),
.B(n_6),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_331),
.A2(n_342),
.B1(n_341),
.B2(n_321),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_328),
.B(n_64),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_343),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_345),
.B(n_353),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_385),
.B(n_341),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_372),
.B(n_341),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_387),
.B(n_341),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_321),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_363),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_391),
.B(n_321),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_369),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_394),
.B(n_335),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_373),
.B(n_351),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_394),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_369),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_402),
.B(n_335),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_363),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_376),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_376),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_390),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_380),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_402),
.B(n_335),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_370),
.B(n_338),
.Y(n_449)
);

A2O1A1Ixp33_ASAP7_75t_SL g450 ( 
.A1(n_409),
.A2(n_302),
.B(n_314),
.C(n_326),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_368),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_343),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_423),
.Y(n_453)
);

BUFx12f_ASAP7_75t_L g454 ( 
.A(n_408),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_366),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_392),
.Y(n_456)
);

NAND2xp33_ASAP7_75t_SL g457 ( 
.A(n_423),
.B(n_331),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_423),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_418),
.B(n_415),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_396),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_406),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_R g462 ( 
.A(n_377),
.B(n_342),
.Y(n_462)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_378),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_404),
.B(n_303),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_367),
.B(n_336),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_386),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_410),
.B(n_308),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_395),
.B(n_400),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_425),
.A2(n_317),
.B1(n_356),
.B2(n_342),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_386),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_397),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_429),
.Y(n_472)
);

NOR3xp33_ASAP7_75t_SL g473 ( 
.A(n_371),
.B(n_303),
.C(n_296),
.Y(n_473)
);

NOR3xp33_ASAP7_75t_SL g474 ( 
.A(n_382),
.B(n_417),
.C(n_364),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_R g475 ( 
.A(n_378),
.B(n_317),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_420),
.A2(n_356),
.B1(n_344),
.B2(n_358),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_374),
.Y(n_477)
);

NAND2x1p5_ASAP7_75t_L g478 ( 
.A(n_379),
.B(n_296),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_396),
.B(n_410),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_413),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_383),
.Y(n_481)
);

BUFx4_ASAP7_75t_SL g482 ( 
.A(n_365),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_413),
.Y(n_483)
);

CKINVDCx11_ASAP7_75t_R g484 ( 
.A(n_378),
.Y(n_484)
);

NOR3xp33_ASAP7_75t_SL g485 ( 
.A(n_417),
.B(n_305),
.C(n_311),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_389),
.Y(n_486)
);

OR2x6_ASAP7_75t_L g487 ( 
.A(n_378),
.B(n_305),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_365),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_478),
.A2(n_430),
.B(n_405),
.Y(n_489)
);

AOI211x1_ASAP7_75t_L g490 ( 
.A1(n_465),
.A2(n_398),
.B(n_364),
.C(n_414),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_484),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_365),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_435),
.Y(n_493)
);

OAI21x1_ASAP7_75t_L g494 ( 
.A1(n_478),
.A2(n_430),
.B(n_403),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_443),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_440),
.B(n_384),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_478),
.A2(n_411),
.B(n_412),
.Y(n_497)
);

AO31x2_ASAP7_75t_L g498 ( 
.A1(n_448),
.A2(n_362),
.A3(n_424),
.B(n_416),
.Y(n_498)
);

CKINVDCx11_ASAP7_75t_R g499 ( 
.A(n_484),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_453),
.A2(n_421),
.B(n_422),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_453),
.A2(n_428),
.B(n_379),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_432),
.A2(n_427),
.B1(n_365),
.B2(n_393),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_435),
.Y(n_503)
);

AO32x2_ASAP7_75t_L g504 ( 
.A1(n_440),
.A2(n_407),
.A3(n_316),
.B1(n_318),
.B2(n_375),
.Y(n_504)
);

OAI21xp33_ASAP7_75t_L g505 ( 
.A1(n_439),
.A2(n_399),
.B(n_388),
.Y(n_505)
);

A2O1A1Ixp33_ASAP7_75t_L g506 ( 
.A1(n_474),
.A2(n_407),
.B(n_381),
.C(n_398),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_461),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_453),
.A2(n_419),
.B(n_344),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_479),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_466),
.A2(n_419),
.B(n_326),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_449),
.A2(n_311),
.B(n_356),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_460),
.B(n_356),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_460),
.B(n_356),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_466),
.A2(n_326),
.B(n_314),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_447),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_466),
.A2(n_326),
.B(n_314),
.Y(n_516)
);

CKINVDCx6p67_ASAP7_75t_R g517 ( 
.A(n_454),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_468),
.A2(n_316),
.B(n_318),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_437),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_459),
.A2(n_359),
.B1(n_314),
.B2(n_358),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_458),
.A2(n_318),
.B(n_316),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_438),
.A2(n_356),
.B(n_349),
.Y(n_522)
);

AOI21x1_ASAP7_75t_L g523 ( 
.A1(n_452),
.A2(n_301),
.B(n_304),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_486),
.B(n_339),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_458),
.A2(n_316),
.B(n_318),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_483),
.A2(n_355),
.B(n_352),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_434),
.B(n_349),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_434),
.B(n_349),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_436),
.B(n_358),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_458),
.A2(n_319),
.B(n_359),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_436),
.B(n_352),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_431),
.A2(n_319),
.B(n_359),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_433),
.A2(n_319),
.B(n_359),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_476),
.A2(n_319),
.B(n_359),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_457),
.A2(n_319),
.B(n_358),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_477),
.B(n_352),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_495),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_505),
.A2(n_492),
.B1(n_442),
.B2(n_464),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_529),
.B(n_442),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_499),
.Y(n_540)
);

AOI22x1_ASAP7_75t_L g541 ( 
.A1(n_511),
.A2(n_481),
.B1(n_470),
.B2(n_445),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_509),
.A2(n_467),
.B1(n_488),
.B2(n_513),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_512),
.B(n_488),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_515),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_507),
.A2(n_455),
.B1(n_451),
.B2(n_454),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_509),
.A2(n_488),
.B1(n_437),
.B2(n_441),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_495),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_508),
.A2(n_483),
.B(n_445),
.Y(n_548)
);

AOI21x1_ASAP7_75t_L g549 ( 
.A1(n_523),
.A2(n_471),
.B(n_472),
.Y(n_549)
);

OAI21x1_ASAP7_75t_L g550 ( 
.A1(n_508),
.A2(n_483),
.B(n_470),
.Y(n_550)
);

OAI21x1_ASAP7_75t_SL g551 ( 
.A1(n_522),
.A2(n_502),
.B(n_527),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_506),
.A2(n_469),
.B1(n_485),
.B2(n_441),
.Y(n_552)
);

BUFx8_ASAP7_75t_SL g553 ( 
.A(n_491),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_514),
.A2(n_443),
.B(n_480),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_496),
.B(n_451),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_519),
.B(n_446),
.Y(n_556)
);

OAI21x1_ASAP7_75t_L g557 ( 
.A1(n_514),
.A2(n_480),
.B(n_444),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_493),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_506),
.A2(n_457),
.B(n_450),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_503),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g561 ( 
.A1(n_516),
.A2(n_444),
.B(n_456),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_519),
.A2(n_455),
.B1(n_473),
.B2(n_441),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_499),
.Y(n_563)
);

OAI21x1_ASAP7_75t_L g564 ( 
.A1(n_516),
.A2(n_355),
.B(n_307),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_517),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_528),
.B(n_437),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_491),
.Y(n_567)
);

BUFx10_ASAP7_75t_L g568 ( 
.A(n_490),
.Y(n_568)
);

OAI21x1_ASAP7_75t_L g569 ( 
.A1(n_510),
.A2(n_355),
.B(n_307),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_526),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_531),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_524),
.A2(n_441),
.B1(n_437),
.B2(n_462),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_536),
.B(n_437),
.Y(n_573)
);

AOI21xp33_ASAP7_75t_L g574 ( 
.A1(n_520),
.A2(n_401),
.B(n_441),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_L g575 ( 
.A1(n_534),
.A2(n_487),
.B(n_301),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_501),
.A2(n_307),
.B(n_309),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_497),
.B(n_463),
.Y(n_577)
);

OAI21x1_ASAP7_75t_L g578 ( 
.A1(n_501),
.A2(n_309),
.B(n_322),
.Y(n_578)
);

OAI22xp33_ASAP7_75t_L g579 ( 
.A1(n_571),
.A2(n_487),
.B1(n_463),
.B2(n_504),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_547),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_571),
.B(n_463),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_SL g582 ( 
.A1(n_555),
.A2(n_475),
.B1(n_504),
.B2(n_482),
.Y(n_582)
);

A2O1A1Ixp33_ASAP7_75t_L g583 ( 
.A1(n_552),
.A2(n_504),
.B(n_497),
.C(n_532),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_551),
.A2(n_518),
.B(n_500),
.Y(n_584)
);

OR2x6_ASAP7_75t_L g585 ( 
.A(n_543),
.B(n_487),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_538),
.A2(n_487),
.B1(n_533),
.B2(n_530),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_539),
.B(n_498),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_556),
.B(n_535),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_544),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_556),
.B(n_489),
.Y(n_590)
);

AND2x2_ASAP7_75t_SL g591 ( 
.A(n_577),
.B(n_504),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_558),
.Y(n_592)
);

NAND4xp25_ASAP7_75t_L g593 ( 
.A(n_562),
.B(n_7),
.C(n_9),
.D(n_10),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_544),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_539),
.A2(n_489),
.B1(n_494),
.B2(n_304),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_558),
.Y(n_596)
);

BUFx2_ASAP7_75t_SL g597 ( 
.A(n_567),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_566),
.B(n_498),
.Y(n_598)
);

INVxp67_ASAP7_75t_SL g599 ( 
.A(n_560),
.Y(n_599)
);

AOI221xp5_ASAP7_75t_L g600 ( 
.A1(n_551),
.A2(n_325),
.B1(n_322),
.B2(n_309),
.C(n_521),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_559),
.A2(n_500),
.B(n_525),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_566),
.B(n_560),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_574),
.A2(n_494),
.B1(n_325),
.B2(n_322),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_547),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_537),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_537),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_573),
.Y(n_607)
);

OAI22xp33_ASAP7_75t_L g608 ( 
.A1(n_540),
.A2(n_563),
.B1(n_565),
.B2(n_541),
.Y(n_608)
);

OAI21x1_ASAP7_75t_L g609 ( 
.A1(n_576),
.A2(n_498),
.B(n_98),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_545),
.A2(n_498),
.B1(n_11),
.B2(n_12),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_561),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_542),
.A2(n_572),
.B1(n_546),
.B2(n_543),
.Y(n_612)
);

NAND2x1_ASAP7_75t_L g613 ( 
.A(n_543),
.B(n_577),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_561),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_543),
.B(n_9),
.Y(n_615)
);

OAI21x1_ASAP7_75t_L g616 ( 
.A1(n_576),
.A2(n_96),
.B(n_145),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_557),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_549),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_568),
.B(n_11),
.Y(n_619)
);

AOI21xp33_ASAP7_75t_L g620 ( 
.A1(n_541),
.A2(n_12),
.B(n_13),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_549),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_568),
.B(n_13),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_568),
.B(n_14),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_553),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_565),
.B(n_540),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_575),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g627 ( 
.A1(n_577),
.A2(n_104),
.B(n_144),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_577),
.B(n_65),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_570),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_557),
.B(n_20),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_593),
.A2(n_570),
.B1(n_554),
.B2(n_550),
.Y(n_631)
);

BUFx12f_ASAP7_75t_L g632 ( 
.A(n_625),
.Y(n_632)
);

AOI221xp5_ASAP7_75t_L g633 ( 
.A1(n_626),
.A2(n_570),
.B1(n_22),
.B2(n_23),
.C(n_24),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_592),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_607),
.B(n_21),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_601),
.A2(n_550),
.B(n_548),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_602),
.B(n_21),
.Y(n_637)
);

NAND2x1_ASAP7_75t_L g638 ( 
.A(n_588),
.B(n_578),
.Y(n_638)
);

AOI222xp33_ASAP7_75t_L g639 ( 
.A1(n_624),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.C1(n_26),
.C2(n_27),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_584),
.A2(n_578),
.B(n_548),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_615),
.B(n_66),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_SL g642 ( 
.A1(n_629),
.A2(n_554),
.B1(n_564),
.B2(n_569),
.Y(n_642)
);

BUFx6f_ASAP7_75t_SL g643 ( 
.A(n_628),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_599),
.Y(n_644)
);

OAI211xp5_ASAP7_75t_SL g645 ( 
.A1(n_624),
.A2(n_25),
.B(n_27),
.C(n_28),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_596),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_599),
.Y(n_647)
);

OAI211xp5_ASAP7_75t_L g648 ( 
.A1(n_626),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_648)
);

OA21x2_ASAP7_75t_L g649 ( 
.A1(n_583),
.A2(n_564),
.B(n_569),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_610),
.A2(n_29),
.B1(n_67),
.B2(n_68),
.Y(n_650)
);

OAI211xp5_ASAP7_75t_SL g651 ( 
.A1(n_619),
.A2(n_69),
.B(n_70),
.C(n_72),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_SL g652 ( 
.A1(n_612),
.A2(n_73),
.B1(n_75),
.B2(n_77),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_620),
.A2(n_146),
.B1(n_79),
.B2(n_80),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_581),
.A2(n_78),
.B1(n_84),
.B2(n_86),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_589),
.B(n_87),
.Y(n_655)
);

AOI21xp33_ASAP7_75t_SL g656 ( 
.A1(n_608),
.A2(n_90),
.B(n_91),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_587),
.B(n_92),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_598),
.B(n_94),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_583),
.A2(n_99),
.B(n_100),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_594),
.B(n_102),
.Y(n_660)
);

OAI22xp33_ASAP7_75t_L g661 ( 
.A1(n_622),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_606),
.Y(n_662)
);

AOI221xp5_ASAP7_75t_L g663 ( 
.A1(n_623),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.C(n_115),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_630),
.A2(n_582),
.B1(n_597),
.B2(n_608),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_613),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_580),
.B(n_116),
.Y(n_666)
);

BUFx12f_ASAP7_75t_L g667 ( 
.A(n_628),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_605),
.B(n_117),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_644),
.B(n_621),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_665),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_634),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_665),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_634),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_646),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_646),
.B(n_591),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_662),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_647),
.B(n_591),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_658),
.B(n_590),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_657),
.B(n_590),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_664),
.B(n_582),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_649),
.Y(n_681)
);

INVx4_ASAP7_75t_R g682 ( 
.A(n_643),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_665),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_638),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_645),
.A2(n_588),
.B1(n_586),
.B2(n_630),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_632),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_640),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_640),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_649),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_664),
.B(n_618),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_649),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_668),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_637),
.B(n_579),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_667),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_692),
.B(n_631),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_671),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_692),
.B(n_631),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_669),
.B(n_611),
.Y(n_698)
);

INVx5_ASAP7_75t_L g699 ( 
.A(n_681),
.Y(n_699)
);

OAI211xp5_ASAP7_75t_L g700 ( 
.A1(n_680),
.A2(n_639),
.B(n_648),
.C(n_633),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_671),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_694),
.Y(n_702)
);

OAI31xp33_ASAP7_75t_L g703 ( 
.A1(n_680),
.A2(n_661),
.A3(n_650),
.B(n_651),
.Y(n_703)
);

AO21x2_ASAP7_75t_L g704 ( 
.A1(n_681),
.A2(n_636),
.B(n_659),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_670),
.B(n_614),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_675),
.B(n_611),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_670),
.B(n_617),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_693),
.A2(n_650),
.B1(n_652),
.B2(n_643),
.Y(n_708)
);

AOI33xp33_ASAP7_75t_L g709 ( 
.A1(n_676),
.A2(n_661),
.A3(n_653),
.B1(n_660),
.B2(n_655),
.B3(n_579),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_692),
.B(n_635),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_706),
.B(n_675),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_696),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_696),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_706),
.B(n_677),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_701),
.B(n_671),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_698),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_705),
.B(n_677),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_710),
.B(n_693),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_705),
.B(n_683),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_718),
.B(n_695),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_716),
.A2(n_700),
.B1(n_643),
.B2(n_708),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_717),
.B(n_699),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_712),
.Y(n_723)
);

NOR3x1_ASAP7_75t_L g724 ( 
.A(n_713),
.B(n_686),
.C(n_694),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_720),
.B(n_702),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_724),
.B(n_717),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_721),
.A2(n_703),
.B1(n_704),
.B2(n_667),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_726),
.Y(n_728)
);

AOI211xp5_ASAP7_75t_L g729 ( 
.A1(n_725),
.A2(n_703),
.B(n_656),
.C(n_654),
.Y(n_729)
);

OAI221xp5_ASAP7_75t_L g730 ( 
.A1(n_727),
.A2(n_686),
.B1(n_685),
.B2(n_723),
.C(n_697),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_728),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_730),
.Y(n_732)
);

OAI211xp5_ASAP7_75t_L g733 ( 
.A1(n_732),
.A2(n_729),
.B(n_685),
.C(n_663),
.Y(n_733)
);

NAND3xp33_ASAP7_75t_L g734 ( 
.A(n_731),
.B(n_709),
.C(n_653),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_731),
.Y(n_735)
);

NOR2x1_ASAP7_75t_L g736 ( 
.A(n_735),
.B(n_722),
.Y(n_736)
);

NAND4xp25_ASAP7_75t_SL g737 ( 
.A(n_733),
.B(n_722),
.C(n_719),
.D(n_682),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_734),
.B(n_714),
.Y(n_738)
);

OAI21x1_ASAP7_75t_L g739 ( 
.A1(n_735),
.A2(n_719),
.B(n_715),
.Y(n_739)
);

AOI211xp5_ASAP7_75t_L g740 ( 
.A1(n_733),
.A2(n_641),
.B(n_690),
.C(n_684),
.Y(n_740)
);

AOI221xp5_ASAP7_75t_L g741 ( 
.A1(n_733),
.A2(n_690),
.B1(n_704),
.B2(n_683),
.C(n_684),
.Y(n_741)
);

OAI21xp33_ASAP7_75t_L g742 ( 
.A1(n_737),
.A2(n_670),
.B(n_672),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_736),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_741),
.A2(n_699),
.B(n_672),
.C(n_714),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_740),
.B(n_666),
.C(n_699),
.Y(n_745)
);

AOI222xp33_ASAP7_75t_L g746 ( 
.A1(n_739),
.A2(n_632),
.B1(n_699),
.B2(n_711),
.C1(n_676),
.C2(n_705),
.Y(n_746)
);

O2A1O1Ixp33_ASAP7_75t_SL g747 ( 
.A1(n_738),
.A2(n_682),
.B(n_715),
.C(n_687),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_738),
.Y(n_748)
);

AO22x1_ASAP7_75t_L g749 ( 
.A1(n_743),
.A2(n_699),
.B1(n_711),
.B2(n_705),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_748),
.A2(n_704),
.B(n_687),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_742),
.B(n_707),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_745),
.Y(n_752)
);

OAI322xp33_ASAP7_75t_L g753 ( 
.A1(n_747),
.A2(n_698),
.A3(n_669),
.B1(n_691),
.B2(n_689),
.C1(n_681),
.C2(n_688),
.Y(n_753)
);

OAI221xp5_ASAP7_75t_L g754 ( 
.A1(n_744),
.A2(n_746),
.B1(n_699),
.B2(n_585),
.C(n_688),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_743),
.Y(n_755)
);

NOR2x1p5_ASAP7_75t_L g756 ( 
.A(n_755),
.B(n_627),
.Y(n_756)
);

NOR3xp33_ASAP7_75t_SL g757 ( 
.A(n_754),
.B(n_600),
.C(n_674),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_752),
.B(n_674),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_751),
.A2(n_707),
.B1(n_585),
.B2(n_679),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_749),
.B(n_678),
.Y(n_760)
);

NAND5xp2_ASAP7_75t_L g761 ( 
.A(n_750),
.B(n_679),
.C(n_678),
.D(n_603),
.E(n_595),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_753),
.B(n_707),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_755),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_755),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_763),
.Y(n_765)
);

NAND4xp75_ASAP7_75t_L g766 ( 
.A(n_764),
.B(n_758),
.C(n_760),
.D(n_762),
.Y(n_766)
);

AOI22x1_ASAP7_75t_L g767 ( 
.A1(n_756),
.A2(n_673),
.B1(n_707),
.B2(n_604),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_761),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_757),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_SL g770 ( 
.A1(n_759),
.A2(n_673),
.B1(n_585),
.B2(n_691),
.Y(n_770)
);

NOR3xp33_ASAP7_75t_L g771 ( 
.A(n_759),
.B(n_616),
.C(n_609),
.Y(n_771)
);

NAND5xp2_ASAP7_75t_L g772 ( 
.A(n_764),
.B(n_603),
.C(n_595),
.D(n_642),
.E(n_123),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_765),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_766),
.Y(n_774)
);

AO22x2_ASAP7_75t_L g775 ( 
.A1(n_769),
.A2(n_673),
.B1(n_691),
.B2(n_689),
.Y(n_775)
);

AOI221xp5_ASAP7_75t_L g776 ( 
.A1(n_768),
.A2(n_770),
.B1(n_772),
.B2(n_771),
.C(n_767),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_765),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_774),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_773),
.Y(n_779)
);

AOI21x1_ASAP7_75t_L g780 ( 
.A1(n_778),
.A2(n_779),
.B(n_777),
.Y(n_780)
);

XNOR2xp5_ASAP7_75t_L g781 ( 
.A(n_780),
.B(n_776),
.Y(n_781)
);

AOI221xp5_ASAP7_75t_L g782 ( 
.A1(n_781),
.A2(n_775),
.B1(n_689),
.B2(n_121),
.C(n_124),
.Y(n_782)
);

OAI221xp5_ASAP7_75t_SL g783 ( 
.A1(n_782),
.A2(n_119),
.B1(n_120),
.B2(n_125),
.C(n_129),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_783),
.Y(n_784)
);

OAI221xp5_ASAP7_75t_R g785 ( 
.A1(n_784),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.C(n_134),
.Y(n_785)
);

AOI211xp5_ASAP7_75t_L g786 ( 
.A1(n_785),
.A2(n_135),
.B(n_136),
.C(n_139),
.Y(n_786)
);


endmodule