module real_jpeg_3995_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_0),
.A2(n_45),
.B1(n_50),
.B2(n_55),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_0),
.A2(n_55),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_0),
.A2(n_55),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_0),
.A2(n_55),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_2),
.A2(n_87),
.B1(n_88),
.B2(n_90),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_2),
.A2(n_46),
.B1(n_87),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_2),
.A2(n_87),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_3),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_3),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_3),
.A2(n_193),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_3),
.A2(n_193),
.B1(n_334),
.B2(n_340),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_3),
.A2(n_193),
.B1(n_390),
.B2(n_406),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_4),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_4),
.B(n_300),
.C(n_302),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_L g304 ( 
.A1(n_4),
.A2(n_305),
.B1(n_306),
.B2(n_308),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_4),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_4),
.B(n_204),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_4),
.A2(n_26),
.B1(n_182),
.B2(n_351),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_4),
.B(n_156),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_4),
.A2(n_265),
.B(n_434),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_5),
.A2(n_283),
.B1(n_285),
.B2(n_286),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_5),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_5),
.A2(n_285),
.B1(n_308),
.B2(n_312),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_5),
.A2(n_285),
.B1(n_340),
.B2(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_5),
.A2(n_247),
.B1(n_285),
.B2(n_390),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_7),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_7),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_7),
.A2(n_64),
.B1(n_101),
.B2(n_105),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_7),
.A2(n_64),
.B1(n_271),
.B2(n_274),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_8),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_8),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_8),
.A2(n_148),
.B1(n_247),
.B2(n_249),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_8),
.A2(n_148),
.B1(n_328),
.B2(n_331),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_8),
.A2(n_148),
.B1(n_308),
.B2(n_393),
.Y(n_392)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_9),
.Y(n_98)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_10),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_10),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_10),
.Y(n_280)
);

BUFx5_ASAP7_75t_L g410 ( 
.A(n_10),
.Y(n_410)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_11),
.Y(n_135)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_11),
.Y(n_139)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_11),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_11),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_11),
.Y(n_263)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_12),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_13),
.Y(n_133)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_13),
.Y(n_136)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_13),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_13),
.Y(n_149)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_13),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_13),
.Y(n_192)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_13),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_13),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_13),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_14),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_14),
.A2(n_38),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_14),
.A2(n_38),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_14),
.A2(n_38),
.B1(n_147),
.B2(n_229),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_233),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_231),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_205),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_19),
.B(n_205),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_159),
.C(n_174),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_20),
.A2(n_21),
.B1(n_159),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_93),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_22),
.B(n_129),
.C(n_158),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_58),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_23),
.A2(n_58),
.B1(n_59),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_23),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_42),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_25),
.A2(n_270),
.B(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_34),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_26),
.A2(n_44),
.B(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_26),
.A2(n_178),
.B(n_180),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_26),
.A2(n_178),
.B1(n_269),
.B2(n_277),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_26),
.A2(n_42),
.B(n_327),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_26),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_26),
.A2(n_182),
.B1(n_339),
.B2(n_351),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_26),
.A2(n_44),
.B(n_180),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_29),
.Y(n_276)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_29),
.Y(n_334)
);

BUFx5_ASAP7_75t_L g340 ( 
.A(n_29),
.Y(n_340)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_33),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_33),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_34),
.Y(n_184)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_36),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_56),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_53),
.Y(n_353)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_54),
.Y(n_330)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_54),
.Y(n_364)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_68),
.B1(n_85),
.B2(n_86),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_61),
.A2(n_166),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_70),
.B1(n_73),
.B2(n_77),
.Y(n_69)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_62),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_63),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g307 ( 
.A(n_63),
.Y(n_307)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_89),
.B1(n_96),
.B2(n_99),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_67),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_68),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_68),
.A2(n_85),
.B1(n_304),
.B2(n_311),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_68),
.A2(n_85),
.B1(n_311),
.B2(n_321),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_68),
.A2(n_85),
.B1(n_321),
.B2(n_392),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_79),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_76),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_77),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_78),
.Y(n_219)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_78),
.Y(n_310)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_78),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_78),
.Y(n_375)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_82),
.Y(n_273)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_85),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_85),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_86),
.Y(n_165)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_89),
.Y(n_170)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_129),
.B1(n_130),
.B2(n_158),
.Y(n_93)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_100),
.B(n_109),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_95),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_95),
.B(n_198),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_95),
.A2(n_202),
.B1(n_404),
.B2(n_405),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_95),
.A2(n_202),
.B1(n_405),
.B2(n_430),
.Y(n_429)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_97),
.Y(n_382)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_100),
.Y(n_209)
);

OAI32xp33_ASAP7_75t_L g372 ( 
.A1(n_101),
.A2(n_373),
.A3(n_376),
.B1(n_379),
.B2(n_380),
.Y(n_372)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_SL g388 ( 
.A1(n_102),
.A2(n_305),
.B(n_379),
.Y(n_388)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_103),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_103),
.Y(n_257)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_108),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_123),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_110),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_110),
.A2(n_204),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_110),
.A2(n_246),
.B(n_253),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_110),
.A2(n_204),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_115),
.B1(n_118),
.B2(n_121),
.Y(n_111)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_114),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_114),
.Y(n_261)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_114),
.Y(n_406)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g378 ( 
.A(n_116),
.Y(n_378)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_140)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_123),
.B(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_126),
.B(n_305),
.Y(n_379)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_128),
.Y(n_211)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_146),
.B(n_150),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_131),
.A2(n_146),
.B1(n_157),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_131),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_131),
.A2(n_157),
.B1(n_433),
.B2(n_435),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_140),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_141),
.Y(n_390)
);

INVx6_ASAP7_75t_SL g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_145),
.Y(n_259)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_147),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_151),
.A2(n_226),
.B(n_227),
.Y(n_225)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_155),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_156),
.A2(n_226),
.B1(n_282),
.B2(n_288),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_157),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_159),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_164),
.B2(n_173),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_160),
.A2(n_161),
.B1(n_225),
.B2(n_230),
.Y(n_224)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_161),
.B(n_164),
.Y(n_223)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B(n_167),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_166),
.B(n_186),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_166),
.A2(n_417),
.B(n_418),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_166),
.A2(n_167),
.B(n_216),
.Y(n_431)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_174),
.B(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_188),
.C(n_196),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_176),
.B(n_241),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_185),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_177),
.B(n_185),
.Y(n_443)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_179),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

INVx3_ASAP7_75t_SL g181 ( 
.A(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_187),
.B(n_305),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_188),
.A2(n_189),
.B1(n_196),
.B2(n_197),
.Y(n_241)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_190),
.Y(n_288)
);

OAI32xp33_ASAP7_75t_L g255 ( 
.A1(n_191),
.A2(n_256),
.A3(n_258),
.B1(n_260),
.B2(n_264),
.Y(n_255)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_202),
.B(n_203),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g457 ( 
.A(n_205),
.Y(n_457)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_207),
.CI(n_222),
.CON(n_205),
.SN(n_205)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_214),
.B(n_221),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_208),
.B(n_214),
.Y(n_221)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_220),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_215),
.Y(n_418)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_218),
.Y(n_384)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_219),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_225),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_289),
.B(n_453),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_236),
.B(n_239),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.C(n_244),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_240),
.B(n_242),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_244),
.B(n_445),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_254),
.C(n_281),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_245),
.B(n_281),
.Y(n_441)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_246),
.Y(n_430)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_254),
.B(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_268),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_255),
.B(n_268),
.Y(n_426)
);

BUFx12f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_282),
.Y(n_435)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_283),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_437),
.B(n_450),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_422),
.B(n_436),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_398),
.B(n_421),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_368),
.B(n_397),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_335),
.B(n_367),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_316),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_296),
.B(n_316),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_303),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_297),
.B(n_303),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_305),
.B(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_SL g306 ( 
.A(n_307),
.Y(n_306)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_315),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_326),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_320),
.B2(n_325),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_318),
.B(n_325),
.C(n_326),
.Y(n_369)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_320),
.Y(n_325)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_327),
.Y(n_342)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx6_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_347),
.B(n_366),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_346),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_346),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_338),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_348),
.A2(n_354),
.B(n_365),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_349),
.B(n_350),
.Y(n_365)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_357),
.B(n_361),
.Y(n_356)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx8_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx4_ASAP7_75t_SL g362 ( 
.A(n_363),
.Y(n_362)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_369),
.B(n_370),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_386),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_387),
.C(n_391),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_385),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_372),
.B(n_385),
.Y(n_415)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx11_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_383),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_391),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_389),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_392),
.Y(n_417)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_399),
.B(n_400),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_401),
.A2(n_402),
.B1(n_413),
.B2(n_414),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_401),
.B(n_416),
.C(n_419),
.Y(n_423)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_407),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_403),
.B(n_408),
.C(n_412),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_408),
.A2(n_409),
.B1(n_411),
.B2(n_412),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_411),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_415),
.A2(n_416),
.B1(n_419),
.B2(n_420),
.Y(n_414)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_415),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_416),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_424),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_428),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_427),
.C(n_428),
.Y(n_447)
);

BUFx24_ASAP7_75t_SL g455 ( 
.A(n_428),
.Y(n_455)
);

FAx1_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_431),
.CI(n_432),
.CON(n_428),
.SN(n_428)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_431),
.C(n_432),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_438),
.B(n_446),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_438),
.A2(n_451),
.B(n_452),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_444),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_444),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_442),
.C(n_443),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_440),
.B(n_449),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_442),
.B(n_443),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_447),
.B(n_448),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);


endmodule