module fake_aes_10642_n_605 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_605);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_605;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_466;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g72 ( .A(n_63), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_26), .Y(n_73) );
CKINVDCx5p33_ASAP7_75t_R g74 ( .A(n_56), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_64), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_24), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_55), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_30), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_16), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_13), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_60), .Y(n_81) );
INVxp67_ASAP7_75t_L g82 ( .A(n_19), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_5), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_57), .Y(n_84) );
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_40), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_19), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_43), .Y(n_87) );
CKINVDCx16_ASAP7_75t_R g88 ( .A(n_32), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_35), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_46), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_59), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_8), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_29), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_5), .Y(n_94) );
CKINVDCx16_ASAP7_75t_R g95 ( .A(n_42), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_45), .Y(n_96) );
INVxp67_ASAP7_75t_L g97 ( .A(n_33), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_68), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_22), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_38), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_12), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_52), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_1), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_25), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_6), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_50), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_10), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_15), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_67), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_21), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_37), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_71), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_6), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_11), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_73), .Y(n_116) );
NOR2x1_ASAP7_75t_L g117 ( .A(n_75), .B(n_0), .Y(n_117) );
INVx3_ASAP7_75t_L g118 ( .A(n_73), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_81), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_81), .Y(n_120) );
OAI21x1_ASAP7_75t_L g121 ( .A1(n_84), .A2(n_28), .B(n_69), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_84), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_87), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_114), .B(n_0), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_88), .B(n_1), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_87), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_98), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_79), .B(n_2), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_72), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_113), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_79), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_85), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_98), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_95), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_113), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_74), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_76), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_77), .Y(n_138) );
AND2x6_ASAP7_75t_L g139 ( .A(n_78), .B(n_31), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_103), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_91), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_96), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_74), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_103), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_89), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_89), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_102), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_90), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_110), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_80), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_80), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_83), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_90), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_83), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_153), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_131), .B(n_105), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_143), .B(n_97), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
NOR2x1_ASAP7_75t_L g159 ( .A(n_154), .B(n_94), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_150), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_146), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_116), .B(n_86), .Y(n_162) );
NAND2x1p5_ASAP7_75t_L g163 ( .A(n_118), .B(n_105), .Y(n_163) );
INVx1_ASAP7_75t_SL g164 ( .A(n_136), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_131), .B(n_147), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_150), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_150), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_147), .B(n_112), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_150), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_151), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_151), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_151), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_151), .Y(n_173) );
INVxp67_ASAP7_75t_L g174 ( .A(n_125), .Y(n_174) );
OR2x2_ASAP7_75t_L g175 ( .A(n_124), .B(n_82), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_151), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_118), .Y(n_177) );
NOR2xp33_ASAP7_75t_R g178 ( .A(n_153), .B(n_99), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_122), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_149), .B(n_99), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_121), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_125), .B(n_86), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_139), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_139), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_149), .B(n_111), .Y(n_185) );
HB1xp67_ASAP7_75t_L g186 ( .A(n_145), .Y(n_186) );
AND2x6_ASAP7_75t_L g187 ( .A(n_125), .B(n_94), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_116), .B(n_115), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_119), .B(n_112), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_122), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_148), .A2(n_109), .B1(n_108), .B2(n_107), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_119), .B(n_106), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_122), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_124), .A2(n_101), .B1(n_92), .B2(n_106), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_118), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_120), .B(n_100), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_118), .Y(n_197) );
INVxp67_ASAP7_75t_L g198 ( .A(n_124), .Y(n_198) );
CKINVDCx11_ASAP7_75t_R g199 ( .A(n_138), .Y(n_199) );
OR2x6_ASAP7_75t_L g200 ( .A(n_128), .B(n_104), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_118), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_152), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_152), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_127), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_184), .B(n_134), .Y(n_205) );
OR2x2_ASAP7_75t_L g206 ( .A(n_198), .B(n_129), .Y(n_206) );
BUFx2_ASAP7_75t_L g207 ( .A(n_187), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_165), .B(n_135), .Y(n_208) );
BUFx2_ASAP7_75t_L g209 ( .A(n_187), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_167), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_192), .B(n_135), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_168), .B(n_120), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_167), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_200), .B(n_117), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_183), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_200), .B(n_117), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_187), .A2(n_130), .B1(n_126), .B2(n_123), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_167), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_180), .B(n_126), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_166), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_163), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_157), .B(n_154), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_163), .Y(n_223) );
NAND3xp33_ASAP7_75t_SL g224 ( .A(n_178), .B(n_132), .C(n_100), .Y(n_224) );
NAND3xp33_ASAP7_75t_SL g225 ( .A(n_164), .B(n_128), .C(n_130), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_161), .Y(n_226) );
BUFx12f_ASAP7_75t_L g227 ( .A(n_199), .Y(n_227) );
NOR3xp33_ASAP7_75t_SL g228 ( .A(n_155), .B(n_123), .C(n_93), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_166), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_187), .A2(n_137), .B1(n_141), .B2(n_139), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_184), .B(n_137), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_171), .Y(n_232) );
NAND3xp33_ASAP7_75t_L g233 ( .A(n_194), .B(n_137), .C(n_141), .Y(n_233) );
NOR3xp33_ASAP7_75t_SL g234 ( .A(n_155), .B(n_140), .C(n_144), .Y(n_234) );
NOR2xp33_ASAP7_75t_R g235 ( .A(n_161), .B(n_139), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_171), .Y(n_236) );
CKINVDCx14_ASAP7_75t_R g237 ( .A(n_186), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_202), .A2(n_141), .B(n_137), .C(n_142), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_200), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_172), .Y(n_240) );
OR2x6_ASAP7_75t_L g241 ( .A(n_200), .B(n_121), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_187), .Y(n_242) );
BUFx2_ASAP7_75t_L g243 ( .A(n_187), .Y(n_243) );
NOR3xp33_ASAP7_75t_SL g244 ( .A(n_191), .B(n_140), .C(n_144), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_200), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_172), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_163), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_156), .B(n_121), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_156), .B(n_152), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_182), .B(n_142), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_173), .Y(n_251) );
AND2x2_ASAP7_75t_SL g252 ( .A(n_184), .B(n_142), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_173), .Y(n_253) );
INVxp67_ASAP7_75t_SL g254 ( .A(n_174), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_179), .Y(n_255) );
NAND2x1p5_ASAP7_75t_L g256 ( .A(n_183), .B(n_141), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_175), .B(n_141), .Y(n_257) );
OR2x6_ASAP7_75t_L g258 ( .A(n_182), .B(n_138), .Y(n_258) );
INVx4_ASAP7_75t_L g259 ( .A(n_187), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_227), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_231), .A2(n_181), .B(n_177), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_220), .Y(n_262) );
INVx2_ASAP7_75t_SL g263 ( .A(n_221), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_259), .B(n_175), .Y(n_264) );
CKINVDCx8_ASAP7_75t_R g265 ( .A(n_239), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_259), .B(n_188), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_214), .A2(n_188), .B1(n_162), .B2(n_185), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_214), .A2(n_188), .B1(n_162), .B2(n_159), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_232), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_214), .B(n_194), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_241), .A2(n_181), .B(n_177), .Y(n_271) );
NAND2x1p5_ASAP7_75t_L g272 ( .A(n_221), .B(n_201), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_206), .B(n_189), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_258), .B(n_162), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_216), .B(n_188), .Y(n_275) );
AND2x2_ASAP7_75t_SL g276 ( .A(n_259), .B(n_207), .Y(n_276) );
BUFx12f_ASAP7_75t_L g277 ( .A(n_227), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_232), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_258), .B(n_162), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_223), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_237), .Y(n_281) );
NAND2x1p5_ASAP7_75t_L g282 ( .A(n_247), .B(n_195), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_258), .B(n_159), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_220), .Y(n_284) );
INVx1_ASAP7_75t_SL g285 ( .A(n_207), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_217), .A2(n_203), .B1(n_202), .B2(n_138), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_229), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_258), .B(n_203), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_241), .A2(n_181), .B(n_201), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_216), .A2(n_196), .B1(n_169), .B2(n_176), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_209), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_215), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_209), .Y(n_293) );
NOR2x1_ASAP7_75t_SL g294 ( .A(n_241), .B(n_197), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_216), .B(n_195), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_250), .B(n_204), .Y(n_296) );
NAND3xp33_ASAP7_75t_L g297 ( .A(n_244), .B(n_181), .C(n_193), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_242), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_235), .B(n_197), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_233), .A2(n_169), .B1(n_160), .B2(n_170), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_206), .B(n_170), .Y(n_301) );
INVx5_ASAP7_75t_L g302 ( .A(n_242), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_249), .B(n_160), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_272), .Y(n_304) );
OAI21x1_ASAP7_75t_SL g305 ( .A1(n_294), .A2(n_230), .B(n_211), .Y(n_305) );
CKINVDCx16_ASAP7_75t_R g306 ( .A(n_277), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_269), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_274), .B(n_249), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_269), .Y(n_309) );
BUFx4f_ASAP7_75t_SL g310 ( .A(n_277), .Y(n_310) );
BUFx4f_ASAP7_75t_SL g311 ( .A(n_277), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_270), .A2(n_279), .B1(n_274), .B2(n_245), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_262), .Y(n_313) );
OAI22xp33_ASAP7_75t_L g314 ( .A1(n_265), .A2(n_245), .B1(n_239), .B2(n_226), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_260), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_267), .B(n_248), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_271), .A2(n_241), .B(n_248), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_280), .B(n_243), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_280), .B(n_266), .Y(n_319) );
OR2x6_ASAP7_75t_L g320 ( .A(n_266), .B(n_243), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_292), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_281), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_301), .A2(n_222), .B1(n_257), .B2(n_225), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_262), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_265), .Y(n_325) );
INVxp67_ASAP7_75t_L g326 ( .A(n_279), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_L g327 ( .A1(n_286), .A2(n_219), .B(n_212), .C(n_238), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_273), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_262), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_288), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_296), .B(n_250), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g332 ( .A1(n_328), .A2(n_254), .B1(n_228), .B2(n_275), .C(n_268), .Y(n_332) );
INVxp67_ASAP7_75t_R g333 ( .A(n_310), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_323), .A2(n_272), .B1(n_276), .B2(n_288), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_317), .A2(n_289), .B(n_294), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_304), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_323), .A2(n_283), .B1(n_224), .B2(n_264), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_307), .Y(n_338) );
AOI211xp5_ASAP7_75t_L g339 ( .A1(n_314), .A2(n_283), .B(n_297), .C(n_208), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_307), .Y(n_340) );
AOI22xp33_ASAP7_75t_SL g341 ( .A1(n_311), .A2(n_276), .B1(n_266), .B2(n_263), .Y(n_341) );
OAI221xp5_ASAP7_75t_L g342 ( .A1(n_312), .A2(n_234), .B1(n_290), .B2(n_297), .C(n_295), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_316), .A2(n_318), .B1(n_319), .B2(n_304), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_321), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_331), .B(n_296), .Y(n_345) );
OAI21xp33_ASAP7_75t_SL g346 ( .A1(n_309), .A2(n_278), .B(n_276), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_313), .Y(n_347) );
AOI22xp33_ASAP7_75t_SL g348 ( .A1(n_306), .A2(n_266), .B1(n_263), .B2(n_298), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_331), .A2(n_248), .B1(n_291), .B2(n_298), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_306), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_316), .A2(n_298), .B1(n_291), .B2(n_278), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_315), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_319), .A2(n_285), .B1(n_293), .B2(n_252), .Y(n_353) );
AO21x2_ASAP7_75t_L g354 ( .A1(n_317), .A2(n_286), .B(n_261), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_308), .A2(n_291), .B1(n_293), .B2(n_252), .Y(n_355) );
AO31x2_ASAP7_75t_L g356 ( .A1(n_309), .A2(n_127), .A3(n_133), .B(n_284), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_347), .B(n_313), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_334), .A2(n_330), .B1(n_308), .B2(n_326), .Y(n_358) );
AOI21xp5_ASAP7_75t_L g359 ( .A1(n_335), .A2(n_329), .B(n_324), .Y(n_359) );
OAI211xp5_ASAP7_75t_L g360 ( .A1(n_332), .A2(n_346), .B(n_341), .C(n_337), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_347), .B(n_329), .Y(n_361) );
OAI31xp33_ASAP7_75t_L g362 ( .A1(n_343), .A2(n_319), .A3(n_327), .B(n_318), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_338), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_344), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_340), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_344), .Y(n_366) );
OAI21xp5_ASAP7_75t_L g367 ( .A1(n_342), .A2(n_327), .B(n_329), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_344), .Y(n_368) );
AOI221x1_ASAP7_75t_L g369 ( .A1(n_344), .A2(n_305), .B1(n_321), .B2(n_324), .C(n_313), .Y(n_369) );
NOR4xp25_ASAP7_75t_SL g370 ( .A(n_350), .B(n_325), .C(n_322), .D(n_305), .Y(n_370) );
OA21x2_ASAP7_75t_L g371 ( .A1(n_351), .A2(n_324), .B(n_127), .Y(n_371) );
AO21x2_ASAP7_75t_L g372 ( .A1(n_354), .A2(n_133), .B(n_303), .Y(n_372) );
NAND3xp33_ASAP7_75t_L g373 ( .A(n_339), .B(n_133), .C(n_304), .Y(n_373) );
OAI211xp5_ASAP7_75t_L g374 ( .A1(n_348), .A2(n_304), .B(n_326), .C(n_137), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_344), .Y(n_375) );
AO21x2_ASAP7_75t_L g376 ( .A1(n_354), .A2(n_284), .B(n_287), .Y(n_376) );
OAI21x1_ASAP7_75t_L g377 ( .A1(n_336), .A2(n_272), .B(n_300), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_356), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_356), .B(n_287), .Y(n_379) );
AOI222xp33_ASAP7_75t_L g380 ( .A1(n_345), .A2(n_319), .B1(n_318), .B2(n_139), .C1(n_285), .C2(n_190), .Y(n_380) );
NAND2xp33_ASAP7_75t_SL g381 ( .A(n_349), .B(n_318), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_356), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_356), .B(n_336), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_356), .B(n_321), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_336), .B(n_321), .Y(n_385) );
OR2x6_ASAP7_75t_L g386 ( .A(n_354), .B(n_321), .Y(n_386) );
AOI222xp33_ASAP7_75t_L g387 ( .A1(n_350), .A2(n_139), .B1(n_204), .B2(n_179), .C1(n_190), .C2(n_193), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_353), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_378), .Y(n_389) );
INVx5_ASAP7_75t_L g390 ( .A(n_384), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_378), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_357), .Y(n_392) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_360), .A2(n_352), .B1(n_355), .B2(n_158), .C(n_176), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_378), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_383), .B(n_321), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_378), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_382), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_382), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_382), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_384), .Y(n_400) );
OR2x6_ASAP7_75t_L g401 ( .A(n_383), .B(n_320), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_383), .B(n_3), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_363), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_384), .Y(n_404) );
NOR2x1_ASAP7_75t_SL g405 ( .A(n_374), .B(n_320), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_379), .B(n_3), .Y(n_406) );
NAND3xp33_ASAP7_75t_L g407 ( .A(n_360), .B(n_352), .C(n_181), .Y(n_407) );
OAI22xp33_ASAP7_75t_L g408 ( .A1(n_373), .A2(n_333), .B1(n_320), .B2(n_282), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_363), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_365), .Y(n_410) );
AND2x4_ASAP7_75t_SL g411 ( .A(n_357), .B(n_320), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_379), .B(n_58), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_388), .B(n_4), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_369), .A2(n_299), .B(n_292), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_388), .B(n_4), .Y(n_415) );
BUFx2_ASAP7_75t_L g416 ( .A(n_364), .Y(n_416) );
NAND3xp33_ASAP7_75t_L g417 ( .A(n_373), .B(n_205), .C(n_292), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_365), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_379), .B(n_7), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_357), .B(n_320), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_372), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_361), .B(n_7), .Y(n_422) );
AND2x2_ASAP7_75t_SL g423 ( .A(n_358), .B(n_333), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_372), .B(n_8), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_372), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_372), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_361), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_361), .B(n_9), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_376), .Y(n_429) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_374), .A2(n_282), .B1(n_213), .B2(n_218), .C(n_210), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_364), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g432 ( .A(n_367), .B(n_292), .C(n_158), .Y(n_432) );
OAI31xp33_ASAP7_75t_L g433 ( .A1(n_381), .A2(n_282), .A3(n_218), .B(n_213), .Y(n_433) );
INVx1_ASAP7_75t_SL g434 ( .A(n_390), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_403), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_392), .B(n_372), .Y(n_436) );
NOR2xp67_ASAP7_75t_SL g437 ( .A(n_424), .B(n_370), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_400), .B(n_376), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_403), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_400), .B(n_376), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_418), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_390), .B(n_386), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_404), .B(n_376), .Y(n_443) );
AOI32xp33_ASAP7_75t_L g444 ( .A1(n_406), .A2(n_381), .A3(n_358), .B1(n_370), .B2(n_12), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_406), .B(n_367), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_409), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_404), .B(n_376), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_390), .B(n_386), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_419), .B(n_362), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_413), .B(n_371), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_390), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_390), .B(n_386), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_427), .B(n_386), .Y(n_453) );
NAND2xp33_ASAP7_75t_R g454 ( .A(n_412), .B(n_371), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_395), .B(n_386), .Y(n_455) );
OR2x6_ASAP7_75t_L g456 ( .A(n_401), .B(n_386), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_419), .B(n_364), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_402), .B(n_385), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_402), .B(n_362), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_410), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_424), .Y(n_461) );
NAND2xp33_ASAP7_75t_SL g462 ( .A(n_412), .B(n_385), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_416), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_413), .B(n_415), .Y(n_464) );
BUFx2_ASAP7_75t_L g465 ( .A(n_431), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_395), .B(n_386), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_431), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_389), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_415), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_411), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_427), .B(n_371), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_401), .B(n_366), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_423), .B(n_371), .Y(n_473) );
OAI33xp33_ASAP7_75t_L g474 ( .A1(n_408), .A2(n_9), .A3(n_10), .B1(n_11), .B2(n_13), .B3(n_14), .Y(n_474) );
AND2x2_ASAP7_75t_SL g475 ( .A(n_412), .B(n_371), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_391), .Y(n_476) );
INVxp67_ASAP7_75t_SL g477 ( .A(n_391), .Y(n_477) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_393), .A2(n_359), .B1(n_366), .B2(n_368), .C(n_210), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_394), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_394), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_401), .B(n_371), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_422), .B(n_359), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_396), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_458), .B(n_401), .Y(n_484) );
OAI22xp33_ASAP7_75t_L g485 ( .A1(n_454), .A2(n_407), .B1(n_423), .B2(n_428), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_446), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_455), .B(n_411), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_464), .B(n_14), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_457), .B(n_396), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_460), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_464), .B(n_15), .Y(n_491) );
NAND4xp25_ASAP7_75t_SL g492 ( .A(n_444), .B(n_433), .C(n_405), .D(n_369), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_435), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_439), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_455), .B(n_425), .Y(n_495) );
OAI33xp33_ASAP7_75t_L g496 ( .A1(n_469), .A2(n_426), .A3(n_425), .B1(n_421), .B2(n_420), .B3(n_429), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_470), .B(n_16), .Y(n_497) );
XNOR2xp5_ASAP7_75t_L g498 ( .A(n_466), .B(n_17), .Y(n_498) );
INVx2_ASAP7_75t_SL g499 ( .A(n_451), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_441), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_449), .A2(n_474), .B1(n_473), .B2(n_459), .Y(n_501) );
OAI322xp33_ASAP7_75t_L g502 ( .A1(n_461), .A2(n_426), .A3(n_421), .B1(n_429), .B2(n_397), .C1(n_398), .C2(n_399), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_438), .B(n_398), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_438), .B(n_440), .Y(n_504) );
OAI211xp5_ASAP7_75t_SL g505 ( .A1(n_482), .A2(n_445), .B(n_436), .C(n_478), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_483), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_473), .A2(n_432), .B1(n_380), .B2(n_417), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_440), .B(n_397), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_466), .B(n_399), .Y(n_509) );
OAI211xp5_ASAP7_75t_L g510 ( .A1(n_462), .A2(n_380), .B(n_387), .C(n_405), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_462), .A2(n_414), .B(n_366), .Y(n_511) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_475), .A2(n_368), .B1(n_366), .B2(n_375), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_477), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_476), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_434), .B(n_17), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_454), .A2(n_387), .B1(n_430), .B2(n_368), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_465), .B(n_18), .Y(n_517) );
NAND2x1_ASAP7_75t_L g518 ( .A(n_456), .B(n_368), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_480), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_443), .B(n_375), .Y(n_520) );
OAI21xp33_ASAP7_75t_L g521 ( .A1(n_450), .A2(n_375), .B(n_377), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_463), .Y(n_522) );
AOI222xp33_ASAP7_75t_L g523 ( .A1(n_450), .A2(n_437), .B1(n_475), .B2(n_447), .C1(n_443), .C2(n_471), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_467), .B(n_377), .Y(n_524) );
OA22x2_ASAP7_75t_L g525 ( .A1(n_456), .A2(n_448), .B1(n_442), .B2(n_452), .Y(n_525) );
AOI21x1_ASAP7_75t_L g526 ( .A1(n_442), .A2(n_377), .B(n_253), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_468), .Y(n_527) );
AOI322xp5_ASAP7_75t_L g528 ( .A1(n_447), .A2(n_18), .A3(n_20), .B1(n_302), .B2(n_255), .C1(n_253), .C2(n_251), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_522), .B(n_472), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_501), .A2(n_456), .B1(n_442), .B2(n_448), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_506), .B(n_471), .Y(n_531) );
NOR3xp33_ASAP7_75t_L g532 ( .A(n_497), .B(n_481), .C(n_479), .Y(n_532) );
OAI21xp33_ASAP7_75t_L g533 ( .A1(n_525), .A2(n_481), .B(n_456), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_504), .B(n_453), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_486), .Y(n_535) );
NOR4xp25_ASAP7_75t_SL g536 ( .A(n_505), .B(n_448), .C(n_452), .D(n_20), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_495), .B(n_479), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_509), .B(n_453), .Y(n_538) );
OAI322xp33_ASAP7_75t_L g539 ( .A1(n_488), .A2(n_468), .A3(n_255), .B1(n_251), .B2(n_246), .C1(n_240), .C2(n_236), .Y(n_539) );
NOR4xp25_ASAP7_75t_SL g540 ( .A(n_513), .B(n_23), .C(n_27), .D(n_34), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_510), .A2(n_302), .B(n_255), .C(n_292), .Y(n_541) );
AOI21xp33_ASAP7_75t_L g542 ( .A1(n_515), .A2(n_36), .B(n_39), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_499), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_490), .Y(n_544) );
XOR2x2_ASAP7_75t_L g545 ( .A(n_498), .B(n_41), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_485), .B(n_292), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_493), .Y(n_547) );
XNOR2x1_ASAP7_75t_L g548 ( .A(n_525), .B(n_44), .Y(n_548) );
XOR2xp5_ASAP7_75t_L g549 ( .A(n_484), .B(n_47), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_514), .B(n_48), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_519), .B(n_49), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_489), .B(n_51), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_487), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_494), .B(n_53), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_527), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_500), .B(n_54), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_503), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_535), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_557), .B(n_523), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_544), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_547), .Y(n_561) );
NOR2xp33_ASAP7_75t_R g562 ( .A(n_543), .B(n_492), .Y(n_562) );
NAND5xp2_ASAP7_75t_L g563 ( .A(n_530), .B(n_528), .C(n_507), .D(n_516), .E(n_491), .Y(n_563) );
NOR2xp33_ASAP7_75t_SL g564 ( .A(n_533), .B(n_517), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_534), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_532), .B(n_508), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_537), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_553), .B(n_492), .Y(n_568) );
OAI22xp33_ASAP7_75t_L g569 ( .A1(n_546), .A2(n_518), .B1(n_503), .B2(n_508), .Y(n_569) );
AOI222xp33_ASAP7_75t_L g570 ( .A1(n_546), .A2(n_496), .B1(n_521), .B2(n_524), .C1(n_520), .C2(n_502), .Y(n_570) );
NOR2x1_ASAP7_75t_L g571 ( .A(n_548), .B(n_511), .Y(n_571) );
XNOR2xp5_ASAP7_75t_L g572 ( .A(n_545), .B(n_512), .Y(n_572) );
AOI222xp33_ASAP7_75t_L g573 ( .A1(n_531), .A2(n_541), .B1(n_529), .B2(n_520), .C1(n_552), .C2(n_555), .Y(n_573) );
AOI211xp5_ASAP7_75t_L g574 ( .A1(n_532), .A2(n_511), .B(n_526), .C(n_65), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_538), .B(n_61), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_555), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_576), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_566), .B(n_529), .Y(n_578) );
A2O1A1Ixp33_ASAP7_75t_L g579 ( .A1(n_568), .A2(n_541), .B(n_542), .C(n_548), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g580 ( .A1(n_568), .A2(n_539), .B1(n_549), .B2(n_551), .C(n_550), .Y(n_580) );
A2O1A1Ixp33_ASAP7_75t_L g581 ( .A1(n_571), .A2(n_536), .B(n_554), .C(n_556), .Y(n_581) );
OA22x2_ASAP7_75t_L g582 ( .A1(n_572), .A2(n_540), .B1(n_66), .B2(n_70), .Y(n_582) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_558), .Y(n_583) );
OR3x1_ASAP7_75t_L g584 ( .A(n_563), .B(n_62), .C(n_302), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_562), .Y(n_585) );
NAND2x1p5_ASAP7_75t_L g586 ( .A(n_575), .B(n_302), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_560), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_559), .A2(n_302), .B1(n_256), .B2(n_236), .Y(n_588) );
OAI211xp5_ASAP7_75t_L g589 ( .A1(n_562), .A2(n_302), .B(n_229), .C(n_240), .Y(n_589) );
NOR3x1_ASAP7_75t_L g590 ( .A(n_564), .B(n_256), .C(n_246), .Y(n_590) );
OAI211xp5_ASAP7_75t_L g591 ( .A1(n_570), .A2(n_215), .B(n_256), .C(n_573), .Y(n_591) );
NAND4xp25_ASAP7_75t_L g592 ( .A(n_574), .B(n_215), .C(n_559), .D(n_575), .Y(n_592) );
AOI211x1_ASAP7_75t_L g593 ( .A1(n_569), .A2(n_215), .B(n_565), .C(n_567), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g594 ( .A1(n_561), .A2(n_215), .B1(n_564), .B2(n_568), .C(n_570), .Y(n_594) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_594), .A2(n_591), .B1(n_585), .B2(n_593), .C(n_577), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_578), .B(n_583), .Y(n_596) );
NAND4xp25_ASAP7_75t_L g597 ( .A(n_581), .B(n_590), .C(n_579), .D(n_592), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_582), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_597), .A2(n_580), .B1(n_588), .B2(n_586), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_596), .Y(n_600) );
XNOR2xp5_ASAP7_75t_L g601 ( .A(n_599), .B(n_598), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_600), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_602), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_603), .A2(n_601), .B1(n_595), .B2(n_584), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_604), .A2(n_589), .B(n_587), .Y(n_605) );
endmodule