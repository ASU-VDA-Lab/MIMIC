module fake_netlist_6_3676_n_1793 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1793);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1793;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_43),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_12),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_72),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_84),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_53),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_63),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_109),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_66),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_37),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_128),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_108),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_5),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_92),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_133),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_44),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_61),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_83),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_54),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_20),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_56),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_65),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_115),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_13),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_95),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_36),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_135),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_80),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_0),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_12),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_14),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_149),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_88),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_59),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_136),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_31),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_55),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_52),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_101),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_90),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_125),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_33),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_26),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_17),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_120),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_36),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_103),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_106),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_37),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_146),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_13),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_153),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_81),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_97),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_9),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_150),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_70),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_7),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_127),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_104),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_25),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_75),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_110),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_152),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_58),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_139),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_86),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_74),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_38),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_32),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_27),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_143),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_99),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_154),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_94),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_26),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_112),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_73),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_130),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_60),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_132),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_14),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_50),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_44),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_121),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_82),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_131),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_67),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_8),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_64),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_45),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_155),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_35),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_51),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_27),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_116),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_77),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_78),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_134),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_32),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_8),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_41),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_15),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_89),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_5),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_54),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_30),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_124),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_85),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_46),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_148),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_9),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_18),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_122),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_102),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_33),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_71),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_43),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_76),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_34),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_40),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_79),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_7),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_38),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_47),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_23),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_137),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_140),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_42),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_19),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_118),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_50),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_69),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_24),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_119),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_0),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_48),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_57),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_19),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_100),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_55),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_113),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_145),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_30),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_46),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_96),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_41),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_98),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_28),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_159),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_163),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_262),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_262),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_1),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_262),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_262),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_262),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_262),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_160),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_170),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_162),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_257),
.B(n_1),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_164),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_167),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_169),
.Y(n_326)
);

INVxp33_ASAP7_75t_SL g327 ( 
.A(n_158),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_262),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_262),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_257),
.B(n_2),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_172),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_285),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_173),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_247),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_182),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_156),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_182),
.Y(n_337)
);

INVxp33_ASAP7_75t_SL g338 ( 
.A(n_168),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_156),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_178),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_245),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_285),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_161),
.B(n_2),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_184),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_190),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_156),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_156),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_156),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_179),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_185),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_179),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_247),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_192),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_157),
.B(n_3),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_198),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_R g356 ( 
.A(n_181),
.B(n_107),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_179),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_285),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_171),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_199),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_179),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_212),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_188),
.B(n_3),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_204),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_222),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_179),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_226),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_229),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_288),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_288),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_245),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_288),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_209),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_288),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_211),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_288),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_216),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_218),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_188),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_350),
.Y(n_380)
);

NAND2xp33_ASAP7_75t_L g381 ( 
.A(n_314),
.B(n_242),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_336),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_325),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_316),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_311),
.B(n_206),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_350),
.B(n_281),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_322),
.B(n_166),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_336),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_311),
.B(n_206),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_339),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_350),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_335),
.B(n_281),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_339),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_313),
.B(n_315),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_316),
.Y(n_395)
);

OAI21x1_ASAP7_75t_L g396 ( 
.A1(n_313),
.A2(n_234),
.B(n_223),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_337),
.B(n_157),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_346),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_346),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_341),
.B(n_177),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_334),
.B(n_175),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_315),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_350),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_347),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_371),
.B(n_177),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_347),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_317),
.Y(n_407)
);

OA21x2_ASAP7_75t_L g408 ( 
.A1(n_348),
.A2(n_277),
.B(n_242),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_348),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_317),
.B(n_223),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_350),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_349),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_318),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_349),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_351),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_318),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_350),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_359),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_351),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_328),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_328),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_368),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_329),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_329),
.B(n_234),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_357),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_332),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_357),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_361),
.B(n_180),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_310),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_354),
.A2(n_252),
.B1(n_228),
.B2(n_291),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_361),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_366),
.B(n_180),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_366),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_369),
.B(n_186),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_369),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_370),
.B(n_186),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_370),
.B(n_191),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_372),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_372),
.B(n_191),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_374),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_334),
.B(n_176),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_374),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_320),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_376),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_403),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g446 ( 
.A(n_383),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_408),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_384),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_408),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_408),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_403),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_429),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_384),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_403),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_408),
.Y(n_455)
);

BUFx4f_ASAP7_75t_L g456 ( 
.A(n_408),
.Y(n_456)
);

NAND3xp33_ASAP7_75t_L g457 ( 
.A(n_387),
.B(n_330),
.C(n_319),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_387),
.B(n_397),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_418),
.B(n_352),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_384),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_397),
.B(n_309),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_408),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_408),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_381),
.A2(n_363),
.B1(n_343),
.B2(n_277),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_418),
.B(n_327),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_381),
.A2(n_363),
.B1(n_343),
.B2(n_229),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_386),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_384),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_384),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_403),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_397),
.B(n_379),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_422),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_408),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_430),
.A2(n_295),
.B1(n_296),
.B2(n_201),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_420),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_397),
.A2(n_306),
.B1(n_260),
.B2(n_250),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_395),
.Y(n_477)
);

AND3x2_ASAP7_75t_L g478 ( 
.A(n_422),
.B(n_358),
.C(n_342),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_403),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_395),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_403),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_394),
.Y(n_482)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_420),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_403),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_400),
.B(n_379),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_392),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_395),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_403),
.Y(n_489)
);

INVxp33_ASAP7_75t_L g490 ( 
.A(n_383),
.Y(n_490)
);

BUFx4f_ASAP7_75t_L g491 ( 
.A(n_420),
.Y(n_491)
);

BUFx10_ASAP7_75t_L g492 ( 
.A(n_426),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_395),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_418),
.B(n_352),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_429),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_394),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_401),
.B(n_338),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_400),
.B(n_321),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_392),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_402),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_392),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_395),
.Y(n_502)
);

NOR3xp33_ASAP7_75t_L g503 ( 
.A(n_401),
.B(n_355),
.C(n_240),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_392),
.B(n_355),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_400),
.B(n_323),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_426),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_402),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_420),
.Y(n_509)
);

INVx8_ASAP7_75t_L g510 ( 
.A(n_400),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_405),
.Y(n_511)
);

INVx5_ASAP7_75t_L g512 ( 
.A(n_403),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_402),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_403),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_420),
.Y(n_515)
);

INVxp33_ASAP7_75t_SL g516 ( 
.A(n_430),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_402),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_407),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_405),
.B(n_324),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_441),
.B(n_326),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_407),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_429),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_407),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_407),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_405),
.B(n_331),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_405),
.B(n_376),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_420),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_420),
.Y(n_528)
);

INVxp67_ASAP7_75t_SL g529 ( 
.A(n_396),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_407),
.Y(n_530)
);

INVxp67_ASAP7_75t_SL g531 ( 
.A(n_396),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_441),
.B(n_340),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_413),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_420),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_430),
.B(n_344),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_443),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_386),
.B(n_345),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_413),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_420),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_413),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_413),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_386),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_427),
.B(n_353),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_385),
.A2(n_373),
.B1(n_367),
.B2(n_375),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_443),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_413),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_396),
.Y(n_547)
);

BUFx6f_ASAP7_75t_SL g548 ( 
.A(n_436),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_434),
.B(n_312),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_416),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_416),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_420),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_L g553 ( 
.A(n_434),
.B(n_356),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_443),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_386),
.B(n_360),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_396),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_434),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_386),
.B(n_364),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_416),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_416),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_427),
.B(n_377),
.Y(n_561)
);

AND2x6_ASAP7_75t_L g562 ( 
.A(n_434),
.B(n_185),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_386),
.B(n_378),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_386),
.B(n_312),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_436),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_439),
.B(n_227),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_428),
.B(n_432),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_439),
.B(n_219),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_436),
.B(n_312),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_416),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_421),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_421),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_439),
.Y(n_573)
);

OAI22xp33_ASAP7_75t_SL g574 ( 
.A1(n_385),
.A2(n_221),
.B1(n_232),
.B2(n_225),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_439),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_427),
.B(n_312),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_436),
.B(n_333),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_436),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_436),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_421),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_421),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_427),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_436),
.B(n_231),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_385),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_421),
.B(n_233),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_423),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_423),
.B(n_236),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_423),
.B(n_237),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_423),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_427),
.B(n_362),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_423),
.Y(n_591)
);

INVxp33_ASAP7_75t_SL g592 ( 
.A(n_428),
.Y(n_592)
);

AO22x2_ASAP7_75t_L g593 ( 
.A1(n_535),
.A2(n_458),
.B1(n_503),
.B2(n_457),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_447),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_579),
.Y(n_595)
);

NOR3xp33_ASAP7_75t_L g596 ( 
.A(n_497),
.B(n_187),
.C(n_183),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_482),
.B(n_389),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_486),
.A2(n_365),
.B1(n_193),
.B2(n_195),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_592),
.B(n_194),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_573),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_486),
.A2(n_389),
.B1(n_410),
.B2(n_424),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_592),
.B(n_196),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_573),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_487),
.B(n_238),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_465),
.B(n_197),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_487),
.B(n_499),
.Y(n_606)
);

OAI22xp33_ASAP7_75t_L g607 ( 
.A1(n_499),
.A2(n_273),
.B1(n_200),
.B2(n_195),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_501),
.B(n_239),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_501),
.B(n_244),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_496),
.B(n_389),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_496),
.B(n_410),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_511),
.B(n_549),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_511),
.B(n_246),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_549),
.B(n_249),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_584),
.B(n_410),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_584),
.B(n_424),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_578),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_456),
.A2(n_424),
.B(n_428),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_471),
.B(n_432),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_567),
.B(n_427),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_L g621 ( 
.A(n_510),
.B(n_185),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_447),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_545),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_449),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_520),
.A2(n_251),
.B1(n_255),
.B2(n_256),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_461),
.B(n_202),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_510),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_567),
.B(n_427),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_510),
.A2(n_307),
.B1(n_267),
.B2(n_263),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_498),
.B(n_203),
.Y(n_630)
);

AND2x4_ASAP7_75t_SL g631 ( 
.A(n_492),
.B(n_193),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_510),
.A2(n_207),
.B1(n_213),
.B2(n_200),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_510),
.B(n_382),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_471),
.B(n_432),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_578),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_526),
.B(n_382),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_449),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_526),
.B(n_382),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_579),
.A2(n_290),
.B1(n_299),
.B2(n_207),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_467),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_467),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_542),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_542),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_450),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_450),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_557),
.A2(n_299),
.B1(n_290),
.B2(n_213),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_455),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_557),
.B(n_258),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_553),
.B(n_388),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_505),
.B(n_208),
.C(n_205),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_455),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_462),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_575),
.B(n_388),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_575),
.B(n_388),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_485),
.B(n_215),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_462),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_463),
.Y(n_657)
);

NOR3xp33_ASAP7_75t_SL g658 ( 
.A(n_459),
.B(n_217),
.C(n_210),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_463),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_525),
.A2(n_294),
.B1(n_274),
.B2(n_305),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_485),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_543),
.B(n_390),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_473),
.A2(n_270),
.B1(n_286),
.B2(n_215),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_561),
.B(n_390),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_576),
.B(n_268),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_544),
.B(n_287),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_590),
.B(n_302),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_556),
.B(n_473),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_566),
.B(n_390),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_529),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_568),
.B(n_393),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_513),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_545),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_492),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_531),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_547),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_582),
.B(n_393),
.Y(n_677)
);

AO22x2_ASAP7_75t_L g678 ( 
.A1(n_516),
.A2(n_221),
.B1(n_225),
.B2(n_232),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_582),
.B(n_393),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_L g680 ( 
.A(n_556),
.B(n_185),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_582),
.B(n_398),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_519),
.B(n_185),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_513),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_523),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_495),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_585),
.B(n_398),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_523),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_506),
.B(n_437),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_533),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_555),
.B(n_270),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_565),
.A2(n_273),
.B1(n_276),
.B2(n_278),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_492),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_565),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_446),
.B(n_220),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_556),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_490),
.B(n_224),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_533),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_565),
.A2(n_276),
.B1(n_278),
.B2(n_286),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_540),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_500),
.Y(n_700)
);

OAI21xp5_ASAP7_75t_L g701 ( 
.A1(n_456),
.A2(n_491),
.B(n_537),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_587),
.B(n_398),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_504),
.B(n_292),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_558),
.B(n_161),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_506),
.B(n_437),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_588),
.B(n_399),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_540),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_563),
.B(n_292),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_556),
.Y(n_709)
);

INVx4_ASAP7_75t_L g710 ( 
.A(n_556),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_500),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_464),
.B(n_437),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_551),
.Y(n_713)
);

NOR2xp67_ASAP7_75t_L g714 ( 
.A(n_577),
.B(n_399),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_551),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_476),
.B(n_292),
.Y(n_716)
);

OAI22xp33_ASAP7_75t_L g717 ( 
.A1(n_474),
.A2(n_235),
.B1(n_308),
.B2(n_174),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_534),
.B(n_399),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_534),
.B(n_539),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_560),
.Y(n_720)
);

INVx8_ASAP7_75t_L g721 ( 
.A(n_548),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_560),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_570),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_565),
.A2(n_292),
.B1(n_306),
.B2(n_308),
.Y(n_724)
);

NAND2xp33_ASAP7_75t_L g725 ( 
.A(n_562),
.B(n_292),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_534),
.B(n_404),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_570),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_466),
.B(n_404),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_456),
.Y(n_729)
);

OAI22xp33_ASAP7_75t_L g730 ( 
.A1(n_474),
.A2(n_214),
.B1(n_165),
.B2(n_303),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_452),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_539),
.B(n_404),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_565),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_539),
.B(n_445),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_445),
.B(n_406),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_571),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_494),
.B(n_230),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_577),
.B(n_532),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_571),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_569),
.B(n_241),
.Y(n_740)
);

INVxp33_ASAP7_75t_L g741 ( 
.A(n_522),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_554),
.B(n_406),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_491),
.A2(n_417),
.B(n_391),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_507),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_445),
.B(n_406),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_507),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_508),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_564),
.B(n_243),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_572),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_472),
.B(n_248),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_472),
.B(n_409),
.Y(n_751)
);

NAND2xp33_ASAP7_75t_L g752 ( 
.A(n_562),
.B(n_253),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_516),
.A2(n_165),
.B1(n_303),
.B2(n_298),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_508),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_574),
.B(n_254),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_583),
.B(n_174),
.Y(n_756)
);

INVx8_ASAP7_75t_L g757 ( 
.A(n_548),
.Y(n_757)
);

NAND2xp33_ASAP7_75t_SL g758 ( 
.A(n_548),
.B(n_189),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_562),
.A2(n_444),
.B1(n_409),
.B2(n_412),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_517),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_517),
.Y(n_761)
);

OAI221xp5_ASAP7_75t_L g762 ( 
.A1(n_574),
.A2(n_189),
.B1(n_214),
.B2(n_235),
.C(n_250),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_572),
.Y(n_763)
);

OAI221xp5_ASAP7_75t_L g764 ( 
.A1(n_518),
.A2(n_260),
.B1(n_265),
.B2(n_269),
.C(n_272),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_672),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_712),
.A2(n_562),
.B1(n_536),
.B2(n_586),
.Y(n_766)
);

AOI21x1_ASAP7_75t_L g767 ( 
.A1(n_618),
.A2(n_521),
.B(n_530),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_597),
.A2(n_491),
.B(n_509),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_600),
.Y(n_769)
);

OAI21xp5_ASAP7_75t_L g770 ( 
.A1(n_610),
.A2(n_521),
.B(n_530),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_611),
.B(n_484),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_688),
.B(n_478),
.Y(n_772)
);

NAND2x1p5_ASAP7_75t_L g773 ( 
.A(n_710),
.B(n_451),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_621),
.A2(n_680),
.B(n_710),
.Y(n_774)
);

AO21x1_ASAP7_75t_L g775 ( 
.A1(n_680),
.A2(n_550),
.B(n_518),
.Y(n_775)
);

INVx8_ASAP7_75t_L g776 ( 
.A(n_721),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_619),
.B(n_484),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_599),
.B(n_475),
.Y(n_778)
);

O2A1O1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_612),
.A2(n_524),
.B(n_541),
.C(n_586),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_621),
.A2(n_483),
.B(n_509),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_710),
.A2(n_483),
.B(n_509),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_623),
.Y(n_782)
);

A2O1A1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_605),
.A2(n_712),
.B(n_634),
.C(n_619),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_634),
.B(n_484),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_633),
.A2(n_475),
.B(n_483),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_593),
.A2(n_562),
.B1(n_524),
.B2(n_541),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_615),
.B(n_514),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_600),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_731),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_616),
.A2(n_661),
.B(n_622),
.C(n_624),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_627),
.A2(n_668),
.B(n_729),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_603),
.B(n_514),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_688),
.B(n_261),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_627),
.A2(n_475),
.B(n_451),
.Y(n_794)
);

INVxp67_ASAP7_75t_L g795 ( 
.A(n_623),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_601),
.A2(n_595),
.B1(n_651),
.B2(n_647),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_673),
.B(n_264),
.Y(n_797)
);

BUFx4f_ASAP7_75t_L g798 ( 
.A(n_721),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_701),
.A2(n_538),
.B(n_546),
.Y(n_799)
);

OR2x2_ASAP7_75t_SL g800 ( 
.A(n_756),
.B(n_265),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_620),
.A2(n_538),
.B(n_546),
.Y(n_801)
);

AO21x1_ASAP7_75t_L g802 ( 
.A1(n_668),
.A2(n_580),
.B(n_559),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_705),
.B(n_266),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_672),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_603),
.B(n_514),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_729),
.A2(n_454),
.B(n_451),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_695),
.A2(n_454),
.B(n_451),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_695),
.A2(n_709),
.B(n_649),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_602),
.B(n_617),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_661),
.B(n_550),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_595),
.A2(n_580),
.B1(n_559),
.B2(n_581),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_695),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_626),
.B(n_581),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_695),
.A2(n_451),
.B(n_454),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_630),
.B(n_589),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_695),
.A2(n_481),
.B(n_489),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_594),
.A2(n_298),
.B(n_284),
.C(n_272),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_709),
.B(n_454),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_594),
.A2(n_284),
.B(n_269),
.C(n_591),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_669),
.B(n_589),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_628),
.A2(n_591),
.B(n_480),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_709),
.A2(n_481),
.B(n_489),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_683),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_709),
.A2(n_481),
.B(n_489),
.Y(n_824)
);

NAND2x1p5_ASAP7_75t_L g825 ( 
.A(n_709),
.B(n_454),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_617),
.B(n_515),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_677),
.A2(n_470),
.B(n_481),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_622),
.A2(n_480),
.B(n_448),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_690),
.A2(n_488),
.B(n_453),
.C(n_460),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_595),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_705),
.B(n_271),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_693),
.B(n_470),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_635),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_679),
.A2(n_470),
.B(n_481),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_681),
.A2(n_489),
.B(n_470),
.Y(n_835)
);

O2A1O1Ixp5_ASAP7_75t_L g836 ( 
.A1(n_708),
.A2(n_448),
.B(n_453),
.C(n_460),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_690),
.A2(n_468),
.B(n_469),
.C(n_477),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_693),
.B(n_470),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_742),
.B(n_275),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_734),
.A2(n_489),
.B(n_479),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_624),
.B(n_515),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_635),
.B(n_515),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_686),
.A2(n_479),
.B(n_512),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_685),
.Y(n_844)
);

O2A1O1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_653),
.A2(n_654),
.B(n_646),
.C(n_606),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_700),
.Y(n_846)
);

NOR3xp33_ASAP7_75t_L g847 ( 
.A(n_738),
.B(n_280),
.C(n_279),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_702),
.A2(n_479),
.B(n_512),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_742),
.B(n_282),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_733),
.B(n_479),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_637),
.B(n_515),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_598),
.B(n_515),
.Y(n_852)
);

AOI21xp33_ASAP7_75t_L g853 ( 
.A1(n_593),
.A2(n_304),
.B(n_300),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_637),
.B(n_528),
.Y(n_854)
);

AOI21x1_ASAP7_75t_L g855 ( 
.A1(n_743),
.A2(n_469),
.B(n_468),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_644),
.B(n_528),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_644),
.A2(n_477),
.B(n_488),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_645),
.A2(n_502),
.B(n_493),
.Y(n_858)
);

AOI222xp33_ASAP7_75t_L g859 ( 
.A1(n_717),
.A2(n_283),
.B1(n_289),
.B2(n_293),
.C1(n_297),
.C2(n_562),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_706),
.A2(n_671),
.B(n_719),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_642),
.A2(n_479),
.B(n_512),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_593),
.A2(n_640),
.B1(n_641),
.B2(n_650),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_642),
.A2(n_512),
.B(n_528),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_733),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_751),
.B(n_493),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_751),
.B(n_528),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_613),
.B(n_694),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_645),
.B(n_528),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_652),
.B(n_502),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_652),
.B(n_562),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_696),
.B(n_4),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_659),
.B(n_409),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_659),
.B(n_412),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_647),
.A2(n_431),
.B1(n_412),
.B2(n_414),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_648),
.B(n_4),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_704),
.B(n_62),
.Y(n_876)
);

INVx5_ASAP7_75t_L g877 ( 
.A(n_721),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_728),
.B(n_431),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_728),
.B(n_431),
.Y(n_879)
);

NOR3xp33_ASAP7_75t_L g880 ( 
.A(n_685),
.B(n_444),
.C(n_414),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_651),
.B(n_414),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_643),
.B(n_512),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_656),
.A2(n_552),
.B(n_527),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_SL g884 ( 
.A1(n_607),
.A2(n_444),
.B(n_415),
.C(n_419),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_700),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_656),
.A2(n_552),
.B(n_527),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_657),
.B(n_415),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_657),
.A2(n_435),
.B(n_419),
.C(n_415),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_643),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_714),
.B(n_670),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_662),
.B(n_419),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_636),
.A2(n_512),
.B(n_552),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_690),
.A2(n_435),
.B(n_433),
.C(n_438),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_678),
.A2(n_435),
.B1(n_438),
.B2(n_433),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_674),
.B(n_438),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_683),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_674),
.B(n_438),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_638),
.A2(n_552),
.B(n_527),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_664),
.A2(n_552),
.B(n_527),
.Y(n_899)
);

AOI21xp33_ASAP7_75t_L g900 ( 
.A1(n_593),
.A2(n_6),
.B(n_10),
.Y(n_900)
);

BUFx8_ASAP7_75t_SL g901 ( 
.A(n_704),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_692),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_735),
.A2(n_552),
.B(n_527),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_684),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_670),
.B(n_433),
.Y(n_905)
);

A2O1A1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_753),
.A2(n_438),
.B(n_433),
.C(n_442),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_675),
.B(n_433),
.Y(n_907)
);

AOI21xp33_ASAP7_75t_L g908 ( 
.A1(n_667),
.A2(n_6),
.B(n_10),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_721),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_711),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_675),
.A2(n_527),
.B(n_433),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_745),
.A2(n_380),
.B(n_391),
.Y(n_912)
);

NAND2x1p5_ASAP7_75t_L g913 ( 
.A(n_676),
.B(n_438),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_676),
.A2(n_438),
.B(n_433),
.Y(n_914)
);

OR2x2_ASAP7_75t_SL g915 ( 
.A(n_756),
.B(n_11),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_655),
.B(n_440),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_762),
.A2(n_442),
.B(n_417),
.C(n_411),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_711),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_692),
.B(n_11),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_718),
.A2(n_417),
.B(n_411),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_744),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_726),
.A2(n_417),
.B(n_411),
.Y(n_922)
);

OAI21xp33_ASAP7_75t_L g923 ( 
.A1(n_596),
.A2(n_442),
.B(n_417),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_704),
.A2(n_442),
.B(n_417),
.C(n_411),
.Y(n_924)
);

NOR2xp67_ASAP7_75t_L g925 ( 
.A(n_625),
.B(n_114),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_658),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_684),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_655),
.B(n_440),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_655),
.B(n_442),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_732),
.A2(n_417),
.B(n_411),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_604),
.A2(n_411),
.B(n_391),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_687),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_608),
.A2(n_411),
.B(n_391),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_609),
.A2(n_391),
.B(n_380),
.Y(n_934)
);

BUFx2_ASAP7_75t_SL g935 ( 
.A(n_687),
.Y(n_935)
);

INVx4_ASAP7_75t_L g936 ( 
.A(n_757),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_744),
.B(n_440),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_689),
.Y(n_938)
);

AO21x1_ASAP7_75t_L g939 ( 
.A1(n_666),
.A2(n_15),
.B(n_16),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_632),
.A2(n_440),
.B1(n_425),
.B2(n_391),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_725),
.A2(n_391),
.B(n_380),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_746),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_678),
.A2(n_440),
.B1(n_425),
.B2(n_380),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_663),
.B(n_380),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_639),
.B(n_746),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_747),
.B(n_754),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_725),
.A2(n_380),
.B(n_440),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_748),
.A2(n_380),
.B(n_440),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_689),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_758),
.A2(n_440),
.B(n_425),
.C(n_18),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_747),
.B(n_440),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_678),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_740),
.A2(n_440),
.B(n_425),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_909),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_SL g955 ( 
.A(n_789),
.B(n_741),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_846),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_809),
.B(n_795),
.Y(n_957)
);

CKINVDCx8_ASAP7_75t_R g958 ( 
.A(n_909),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_774),
.A2(n_703),
.B(n_682),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_860),
.A2(n_665),
.B(n_761),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_783),
.A2(n_754),
.B(n_761),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_809),
.B(n_614),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_783),
.A2(n_760),
.B(n_763),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_865),
.B(n_755),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_778),
.A2(n_629),
.B1(n_691),
.B2(n_698),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_R g966 ( 
.A(n_798),
.B(n_758),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_808),
.A2(n_760),
.B(n_763),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_780),
.A2(n_757),
.B(n_752),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_778),
.A2(n_660),
.B1(n_757),
.B2(n_724),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_839),
.B(n_631),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_771),
.A2(n_757),
.B(n_752),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_SL g972 ( 
.A1(n_871),
.A2(n_764),
.B(n_722),
.C(n_720),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_768),
.A2(n_720),
.B(n_697),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_867),
.B(n_750),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_867),
.A2(n_871),
.B1(n_875),
.B2(n_890),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_885),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_801),
.A2(n_727),
.B(n_749),
.Y(n_977)
);

OAI21xp33_ASAP7_75t_L g978 ( 
.A1(n_849),
.A2(n_631),
.B(n_730),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_876),
.B(n_737),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_910),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_918),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_853),
.A2(n_716),
.B(n_697),
.C(n_699),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_844),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_866),
.B(n_793),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_921),
.Y(n_985)
);

OR2x6_ASAP7_75t_L g986 ( 
.A(n_776),
.B(n_909),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_813),
.A2(n_722),
.B(n_749),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_SL g988 ( 
.A1(n_915),
.A2(n_926),
.B1(n_800),
.B2(n_875),
.Y(n_988)
);

OAI22xp33_ASAP7_75t_L g989 ( 
.A1(n_952),
.A2(n_759),
.B1(n_739),
.B2(n_736),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_845),
.A2(n_852),
.B(n_866),
.C(n_862),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_782),
.B(n_739),
.Y(n_991)
);

AO21x1_ASAP7_75t_L g992 ( 
.A1(n_900),
.A2(n_736),
.B(n_727),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_782),
.B(n_723),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_890),
.B(n_723),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_876),
.B(n_715),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_852),
.A2(n_715),
.B(n_713),
.C(n_707),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_908),
.A2(n_713),
.B(n_707),
.C(n_699),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_847),
.A2(n_678),
.B1(n_425),
.B2(n_147),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_803),
.B(n_425),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_945),
.A2(n_425),
.B1(n_142),
.B2(n_141),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_815),
.A2(n_425),
.B(n_138),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_831),
.B(n_425),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_770),
.A2(n_425),
.B(n_126),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_772),
.B(n_16),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_796),
.A2(n_105),
.B(n_93),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_925),
.A2(n_111),
.B1(n_91),
.B2(n_87),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_864),
.Y(n_1007)
);

BUFx8_ASAP7_75t_L g1008 ( 
.A(n_902),
.Y(n_1008)
);

AOI33xp33_ASAP7_75t_L g1009 ( 
.A1(n_833),
.A2(n_17),
.A3(n_20),
.B1(n_21),
.B2(n_22),
.B3(n_23),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_909),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_949),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_817),
.A2(n_21),
.B(n_22),
.C(n_24),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_911),
.A2(n_68),
.B(n_28),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_864),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_797),
.B(n_25),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_766),
.A2(n_29),
.B(n_31),
.C(n_34),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_817),
.A2(n_29),
.B(n_35),
.C(n_39),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_769),
.B(n_39),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_936),
.B(n_40),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_901),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_788),
.B(n_889),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_776),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_798),
.B(n_42),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_777),
.B(n_45),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_784),
.B(n_891),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_936),
.B(n_47),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_950),
.A2(n_790),
.B(n_880),
.C(n_819),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_790),
.A2(n_48),
.B(n_49),
.C(n_51),
.Y(n_1028)
);

AOI21x1_ASAP7_75t_L g1029 ( 
.A1(n_946),
.A2(n_767),
.B(n_791),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_799),
.A2(n_49),
.B(n_52),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_889),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_786),
.A2(n_842),
.B(n_826),
.C(n_878),
.Y(n_1032)
);

OAI21xp33_ASAP7_75t_SL g1033 ( 
.A1(n_946),
.A2(n_58),
.B(n_914),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_919),
.B(n_830),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_787),
.B(n_879),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_942),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_826),
.A2(n_842),
.B(n_923),
.C(n_779),
.Y(n_1037)
);

NAND2xp33_ASAP7_75t_SL g1038 ( 
.A(n_812),
.B(n_895),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_830),
.A2(n_812),
.B1(n_913),
.B2(n_820),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_810),
.B(n_897),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_765),
.B(n_804),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_939),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_823),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_949),
.Y(n_1044)
);

BUFx10_ASAP7_75t_L g1045 ( 
.A(n_812),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_877),
.B(n_812),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_913),
.A2(n_773),
.B1(n_935),
.B2(n_825),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_776),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_877),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_819),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_896),
.B(n_904),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_877),
.B(n_924),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_927),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_932),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_773),
.A2(n_785),
.B(n_825),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_859),
.A2(n_916),
.B1(n_928),
.B2(n_929),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_807),
.A2(n_824),
.B(n_822),
.Y(n_1057)
);

AOI21xp33_ASAP7_75t_L g1058 ( 
.A1(n_916),
.A2(n_928),
.B(n_870),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_814),
.A2(n_816),
.B(n_781),
.Y(n_1059)
);

NOR3xp33_ASAP7_75t_SL g1060 ( 
.A(n_893),
.B(n_906),
.C(n_832),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_R g1061 ( 
.A(n_877),
.B(n_855),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_938),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_792),
.B(n_805),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_832),
.B(n_838),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_881),
.Y(n_1065)
);

NAND2x1p5_ASAP7_75t_L g1066 ( 
.A(n_838),
.B(n_850),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_894),
.B(n_943),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_850),
.B(n_837),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_894),
.B(n_943),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_841),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_905),
.B(n_907),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_869),
.B(n_872),
.Y(n_1072)
);

NOR3xp33_ASAP7_75t_SL g1073 ( 
.A(n_906),
.B(n_888),
.C(n_818),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_873),
.B(n_887),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_882),
.A2(n_802),
.B1(n_944),
.B2(n_818),
.Y(n_1075)
);

AO21x1_ASAP7_75t_L g1076 ( 
.A1(n_882),
.A2(n_883),
.B(n_886),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_937),
.B(n_888),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_851),
.B(n_856),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_854),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_868),
.A2(n_829),
.B1(n_827),
.B2(n_834),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_948),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_821),
.B(n_835),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_868),
.B(n_951),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_937),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_840),
.A2(n_920),
.B(n_848),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_843),
.B(n_858),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_775),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_SL g1088 ( 
.A1(n_917),
.A2(n_806),
.B(n_794),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_874),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_SL g1090 ( 
.A(n_953),
.B(n_931),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_933),
.B(n_934),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_912),
.A2(n_922),
.B(n_930),
.C(n_836),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_828),
.B(n_857),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_811),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_884),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_884),
.B(n_892),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_941),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_898),
.A2(n_899),
.B(n_861),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_947),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_863),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_903),
.B(n_940),
.Y(n_1101)
);

INVx5_ASAP7_75t_L g1102 ( 
.A(n_986),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1065),
.B(n_984),
.Y(n_1103)
);

BUFx10_ASAP7_75t_L g1104 ( 
.A(n_1020),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_976),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1025),
.B(n_1067),
.Y(n_1106)
);

AOI221x1_ASAP7_75t_L g1107 ( 
.A1(n_1030),
.A2(n_1005),
.B1(n_1013),
.B2(n_990),
.C(n_1003),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_SL g1108 ( 
.A1(n_1032),
.A2(n_1037),
.B(n_969),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_962),
.A2(n_975),
.B(n_974),
.C(n_978),
.Y(n_1109)
);

OR2x2_ASAP7_75t_L g1110 ( 
.A(n_983),
.B(n_970),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_980),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_981),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1082),
.A2(n_968),
.B(n_960),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_967),
.A2(n_1059),
.B(n_1057),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_967),
.A2(n_973),
.B(n_1098),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_985),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_961),
.A2(n_963),
.B(n_1003),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_961),
.A2(n_963),
.B(n_1033),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1069),
.B(n_1035),
.Y(n_1119)
);

CKINVDCx11_ASAP7_75t_R g1120 ( 
.A(n_958),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_1008),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_986),
.Y(n_1122)
);

CKINVDCx16_ASAP7_75t_R g1123 ( 
.A(n_955),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1036),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1048),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_957),
.B(n_1062),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_SL g1127 ( 
.A1(n_1016),
.A2(n_979),
.B(n_972),
.C(n_1095),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_1008),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_960),
.A2(n_1086),
.B(n_1074),
.Y(n_1129)
);

AO21x2_ASAP7_75t_L g1130 ( 
.A1(n_1085),
.A2(n_1098),
.B(n_992),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1085),
.A2(n_1093),
.B(n_1055),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_988),
.B(n_1015),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1030),
.A2(n_1004),
.B(n_1023),
.C(n_965),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1019),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_1013),
.A2(n_1027),
.B(n_1005),
.C(n_998),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1029),
.A2(n_987),
.B(n_977),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_991),
.B(n_993),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_964),
.B(n_1021),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_987),
.A2(n_977),
.B(n_1080),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1040),
.B(n_1079),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1088),
.A2(n_959),
.B(n_1091),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_986),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1101),
.A2(n_996),
.B(n_1096),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1072),
.B(n_1089),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_959),
.A2(n_971),
.B(n_1039),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_SL g1146 ( 
.A(n_1022),
.B(n_1019),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1078),
.A2(n_1047),
.B(n_982),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_SL g1148 ( 
.A(n_1026),
.B(n_1028),
.Y(n_1148)
);

CKINVDCx8_ASAP7_75t_R g1149 ( 
.A(n_1048),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1048),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1071),
.A2(n_1063),
.B(n_1097),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1075),
.A2(n_1073),
.B(n_1060),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_999),
.A2(n_1002),
.B(n_1090),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_954),
.Y(n_1154)
);

OA21x2_ASAP7_75t_L g1155 ( 
.A1(n_1087),
.A2(n_1001),
.B(n_1092),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_1076),
.A2(n_1042),
.A3(n_1001),
.B(n_1000),
.Y(n_1156)
);

INVx2_ASAP7_75t_SL g1157 ( 
.A(n_1026),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1038),
.A2(n_995),
.B(n_1083),
.Y(n_1158)
);

O2A1O1Ixp5_ASAP7_75t_SL g1159 ( 
.A1(n_1031),
.A2(n_1024),
.B(n_1018),
.C(n_1043),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1034),
.B(n_1056),
.Y(n_1160)
);

AOI221xp5_ASAP7_75t_L g1161 ( 
.A1(n_1012),
.A2(n_1017),
.B1(n_1050),
.B2(n_989),
.C(n_994),
.Y(n_1161)
);

INVxp67_ASAP7_75t_L g1162 ( 
.A(n_1053),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_1054),
.B(n_1011),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1066),
.A2(n_997),
.B(n_1051),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1081),
.A2(n_1064),
.B1(n_1006),
.B2(n_1068),
.Y(n_1165)
);

INVx5_ASAP7_75t_L g1166 ( 
.A(n_954),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1094),
.B(n_1070),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1041),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1077),
.A2(n_1068),
.B(n_1058),
.Y(n_1169)
);

NAND3xp33_ASAP7_75t_L g1170 ( 
.A(n_1009),
.B(n_1084),
.C(n_1100),
.Y(n_1170)
);

INVxp67_ASAP7_75t_L g1171 ( 
.A(n_1044),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1007),
.B(n_1014),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1066),
.A2(n_1046),
.B(n_1007),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_SL g1174 ( 
.A(n_1049),
.B(n_1010),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1014),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_954),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1099),
.A2(n_1100),
.B(n_1052),
.Y(n_1177)
);

O2A1O1Ixp5_ASAP7_75t_L g1178 ( 
.A1(n_1052),
.A2(n_1061),
.B(n_1099),
.C(n_966),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1099),
.A2(n_774),
.B(n_710),
.Y(n_1179)
);

OA21x2_ASAP7_75t_L g1180 ( 
.A1(n_1045),
.A2(n_990),
.B(n_1003),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1045),
.A2(n_975),
.B1(n_1069),
.B2(n_1067),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_974),
.B(n_310),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1082),
.A2(n_774),
.B(n_710),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_956),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_SL g1185 ( 
.A(n_958),
.B(n_516),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_1008),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_992),
.A2(n_990),
.A3(n_1076),
.B(n_775),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_974),
.B(n_310),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_962),
.A2(n_871),
.B(n_605),
.C(n_497),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_967),
.A2(n_1059),
.B(n_1057),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1082),
.A2(n_774),
.B(n_710),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1065),
.B(n_984),
.Y(n_1192)
);

AO21x1_ASAP7_75t_L g1193 ( 
.A1(n_1030),
.A2(n_1013),
.B(n_1005),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_992),
.A2(n_990),
.A3(n_1076),
.B(n_775),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1048),
.B(n_986),
.Y(n_1195)
);

AO31x2_ASAP7_75t_L g1196 ( 
.A1(n_992),
.A2(n_990),
.A3(n_1076),
.B(n_775),
.Y(n_1196)
);

CKINVDCx6p67_ASAP7_75t_R g1197 ( 
.A(n_1010),
.Y(n_1197)
);

AO31x2_ASAP7_75t_L g1198 ( 
.A1(n_992),
.A2(n_990),
.A3(n_1076),
.B(n_775),
.Y(n_1198)
);

BUFx12f_ASAP7_75t_L g1199 ( 
.A(n_983),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1082),
.A2(n_774),
.B(n_710),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1082),
.A2(n_774),
.B(n_710),
.Y(n_1201)
);

AO21x2_ASAP7_75t_L g1202 ( 
.A1(n_990),
.A2(n_1003),
.B(n_1085),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_962),
.A2(n_975),
.B(n_974),
.C(n_867),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1082),
.A2(n_774),
.B(n_710),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_975),
.B(n_962),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_974),
.B(n_310),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1082),
.A2(n_774),
.B(n_710),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1082),
.A2(n_774),
.B(n_710),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_974),
.B(n_310),
.Y(n_1209)
);

AO21x1_ASAP7_75t_L g1210 ( 
.A1(n_1030),
.A2(n_1013),
.B(n_1005),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_983),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1082),
.A2(n_774),
.B(n_710),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1065),
.B(n_984),
.Y(n_1213)
);

AOI21xp33_ASAP7_75t_L g1214 ( 
.A1(n_975),
.A2(n_871),
.B(n_605),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1065),
.B(n_984),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_967),
.A2(n_1059),
.B(n_1057),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_983),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1082),
.A2(n_774),
.B(n_710),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_962),
.B(n_809),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_983),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1008),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_970),
.B(n_839),
.Y(n_1222)
);

INVx2_ASAP7_75t_SL g1223 ( 
.A(n_983),
.Y(n_1223)
);

AOI21xp33_ASAP7_75t_L g1224 ( 
.A1(n_975),
.A2(n_871),
.B(n_605),
.Y(n_1224)
);

INVxp67_ASAP7_75t_SL g1225 ( 
.A(n_991),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_967),
.A2(n_1059),
.B(n_1057),
.Y(n_1226)
);

AO31x2_ASAP7_75t_L g1227 ( 
.A1(n_992),
.A2(n_990),
.A3(n_1076),
.B(n_775),
.Y(n_1227)
);

AO31x2_ASAP7_75t_L g1228 ( 
.A1(n_992),
.A2(n_990),
.A3(n_1076),
.B(n_775),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_983),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1082),
.A2(n_774),
.B(n_710),
.Y(n_1230)
);

NAND2x1p5_ASAP7_75t_L g1231 ( 
.A(n_1049),
.B(n_877),
.Y(n_1231)
);

AOI31xp67_ASAP7_75t_L g1232 ( 
.A1(n_1096),
.A2(n_1082),
.A3(n_1093),
.B(n_975),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1065),
.B(n_984),
.Y(n_1233)
);

CKINVDCx11_ASAP7_75t_R g1234 ( 
.A(n_958),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1065),
.B(n_984),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_967),
.A2(n_1059),
.B(n_1057),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_956),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_974),
.A2(n_516),
.B1(n_871),
.B2(n_605),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1082),
.A2(n_774),
.B(n_710),
.Y(n_1239)
);

AO21x1_ASAP7_75t_L g1240 ( 
.A1(n_1030),
.A2(n_1013),
.B(n_1005),
.Y(n_1240)
);

BUFx5_ASAP7_75t_L g1241 ( 
.A(n_1095),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1082),
.A2(n_774),
.B(n_710),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_975),
.B(n_731),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_967),
.A2(n_1059),
.B(n_1057),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1008),
.Y(n_1245)
);

NAND2x1p5_ASAP7_75t_L g1246 ( 
.A(n_1049),
.B(n_877),
.Y(n_1246)
);

BUFx8_ASAP7_75t_L g1247 ( 
.A(n_1121),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_1217),
.Y(n_1248)
);

CKINVDCx11_ASAP7_75t_R g1249 ( 
.A(n_1104),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1134),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1124),
.Y(n_1251)
);

CKINVDCx11_ASAP7_75t_R g1252 ( 
.A(n_1104),
.Y(n_1252)
);

CKINVDCx6p67_ASAP7_75t_R g1253 ( 
.A(n_1120),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1238),
.A2(n_1203),
.B1(n_1219),
.B2(n_1189),
.Y(n_1254)
);

INVx6_ASAP7_75t_L g1255 ( 
.A(n_1166),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1149),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1182),
.A2(n_1206),
.B1(n_1188),
.B2(n_1209),
.Y(n_1257)
);

INVx4_ASAP7_75t_L g1258 ( 
.A(n_1166),
.Y(n_1258)
);

BUFx12f_ASAP7_75t_L g1259 ( 
.A(n_1234),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1205),
.A2(n_1214),
.B1(n_1224),
.B2(n_1132),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1137),
.B(n_1103),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1148),
.A2(n_1152),
.B1(n_1123),
.B2(n_1146),
.Y(n_1262)
);

CKINVDCx11_ASAP7_75t_R g1263 ( 
.A(n_1199),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1214),
.A2(n_1224),
.B1(n_1152),
.B2(n_1160),
.Y(n_1264)
);

CKINVDCx11_ASAP7_75t_R g1265 ( 
.A(n_1186),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1160),
.A2(n_1161),
.B1(n_1210),
.B2(n_1240),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1163),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1223),
.Y(n_1268)
);

INVx4_ASAP7_75t_L g1269 ( 
.A(n_1166),
.Y(n_1269)
);

OAI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1148),
.A2(n_1243),
.B1(n_1146),
.B2(n_1165),
.Y(n_1270)
);

INVx6_ASAP7_75t_L g1271 ( 
.A(n_1166),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1193),
.A2(n_1138),
.B1(n_1170),
.B2(n_1213),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_1211),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_SL g1274 ( 
.A1(n_1185),
.A2(n_1126),
.B1(n_1225),
.B2(n_1222),
.Y(n_1274)
);

BUFx2_ASAP7_75t_SL g1275 ( 
.A(n_1220),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1170),
.A2(n_1235),
.B1(n_1103),
.B2(n_1233),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1192),
.A2(n_1235),
.B1(n_1213),
.B2(n_1233),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1105),
.Y(n_1278)
);

INVx1_ASAP7_75t_SL g1279 ( 
.A(n_1110),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1192),
.A2(n_1215),
.B1(n_1202),
.B2(n_1106),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1111),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1116),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1215),
.A2(n_1202),
.B1(n_1106),
.B2(n_1119),
.Y(n_1283)
);

INVx8_ASAP7_75t_L g1284 ( 
.A(n_1102),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1184),
.Y(n_1285)
);

INVx6_ASAP7_75t_L g1286 ( 
.A(n_1102),
.Y(n_1286)
);

OAI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1167),
.A2(n_1119),
.B1(n_1185),
.B2(n_1144),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1117),
.A2(n_1181),
.B1(n_1169),
.B2(n_1118),
.Y(n_1288)
);

INVx4_ASAP7_75t_L g1289 ( 
.A(n_1102),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1109),
.A2(n_1135),
.B1(n_1108),
.B2(n_1167),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1133),
.A2(n_1140),
.B1(n_1157),
.B2(n_1169),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1168),
.B(n_1144),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_SL g1293 ( 
.A1(n_1117),
.A2(n_1174),
.B1(n_1118),
.B2(n_1181),
.Y(n_1293)
);

CKINVDCx11_ASAP7_75t_R g1294 ( 
.A(n_1221),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1151),
.A2(n_1143),
.B1(n_1237),
.B2(n_1180),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1195),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1174),
.A2(n_1229),
.B1(n_1142),
.B2(n_1102),
.Y(n_1297)
);

INVx6_ASAP7_75t_L g1298 ( 
.A(n_1142),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1175),
.Y(n_1299)
);

BUFx2_ASAP7_75t_SL g1300 ( 
.A(n_1125),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_SL g1301 ( 
.A1(n_1107),
.A2(n_1128),
.B(n_1177),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_1245),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1162),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1142),
.A2(n_1171),
.B1(n_1122),
.B2(n_1158),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_SL g1305 ( 
.A(n_1195),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1142),
.A2(n_1122),
.B1(n_1197),
.B2(n_1180),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1154),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1176),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1143),
.A2(n_1155),
.B1(n_1130),
.B2(n_1129),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1154),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1155),
.A2(n_1130),
.B1(n_1131),
.B2(n_1172),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1127),
.B(n_1159),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1173),
.Y(n_1313)
);

BUFx12f_ASAP7_75t_L g1314 ( 
.A(n_1125),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1154),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1179),
.A2(n_1246),
.B1(n_1231),
.B2(n_1200),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1232),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_SL g1318 ( 
.A1(n_1241),
.A2(n_1147),
.B1(n_1145),
.B2(n_1150),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1153),
.A2(n_1139),
.B1(n_1242),
.B2(n_1208),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1231),
.A2(n_1246),
.B1(n_1239),
.B2(n_1230),
.Y(n_1320)
);

BUFx8_ASAP7_75t_L g1321 ( 
.A(n_1150),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1183),
.A2(n_1218),
.B1(n_1191),
.B2(n_1204),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1241),
.Y(n_1323)
);

CKINVDCx11_ASAP7_75t_R g1324 ( 
.A(n_1150),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1201),
.A2(n_1207),
.B1(n_1212),
.B2(n_1164),
.Y(n_1325)
);

CKINVDCx11_ASAP7_75t_R g1326 ( 
.A(n_1241),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1187),
.B(n_1196),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1187),
.B(n_1196),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1136),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1178),
.A2(n_1141),
.B1(n_1113),
.B2(n_1115),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1114),
.A2(n_1216),
.B1(n_1190),
.B2(n_1236),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1194),
.B(n_1196),
.Y(n_1332)
);

BUFx8_ASAP7_75t_L g1333 ( 
.A(n_1194),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1198),
.Y(n_1334)
);

BUFx8_ASAP7_75t_L g1335 ( 
.A(n_1198),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1198),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1227),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1227),
.Y(n_1338)
);

BUFx12f_ASAP7_75t_L g1339 ( 
.A(n_1227),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1226),
.A2(n_1244),
.B1(n_1156),
.B2(n_1228),
.Y(n_1340)
);

BUFx12f_ASAP7_75t_L g1341 ( 
.A(n_1228),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1228),
.B(n_1156),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1156),
.Y(n_1343)
);

CKINVDCx11_ASAP7_75t_R g1344 ( 
.A(n_1104),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1134),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1112),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1112),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1180),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1217),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1243),
.B(n_1140),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1238),
.A2(n_1203),
.B1(n_1219),
.B2(n_975),
.Y(n_1351)
);

NAND2x1p5_ASAP7_75t_L g1352 ( 
.A(n_1102),
.B(n_1142),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1189),
.A2(n_1224),
.B(n_1214),
.Y(n_1353)
);

CKINVDCx11_ASAP7_75t_R g1354 ( 
.A(n_1104),
.Y(n_1354)
);

NAND2x1p5_ASAP7_75t_L g1355 ( 
.A(n_1102),
.B(n_1142),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1217),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1182),
.A2(n_516),
.B1(n_1206),
.B2(n_1188),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1102),
.Y(n_1358)
);

BUFx10_ASAP7_75t_L g1359 ( 
.A(n_1126),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1219),
.B(n_1137),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1217),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1112),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1222),
.B(n_793),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1120),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1205),
.A2(n_1238),
.B1(n_1224),
.B2(n_1214),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1205),
.A2(n_1238),
.B1(n_1224),
.B2(n_1214),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1238),
.A2(n_1203),
.B1(n_1219),
.B2(n_975),
.Y(n_1367)
);

INVx3_ASAP7_75t_SL g1368 ( 
.A(n_1123),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1238),
.A2(n_1203),
.B1(n_1219),
.B2(n_975),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1112),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1112),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1205),
.A2(n_1238),
.B1(n_1224),
.B2(n_1214),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1189),
.A2(n_1224),
.B(n_1214),
.Y(n_1373)
);

BUFx10_ASAP7_75t_L g1374 ( 
.A(n_1126),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1205),
.A2(n_1238),
.B1(n_1224),
.B2(n_1214),
.Y(n_1375)
);

AND2x4_ASAP7_75t_SL g1376 ( 
.A(n_1211),
.B(n_1220),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1336),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1337),
.Y(n_1378)
);

AO21x2_ASAP7_75t_L g1379 ( 
.A1(n_1353),
.A2(n_1373),
.B(n_1312),
.Y(n_1379)
);

OAI222xp33_ASAP7_75t_L g1380 ( 
.A1(n_1262),
.A2(n_1254),
.B1(n_1369),
.B2(n_1351),
.C1(n_1367),
.C2(n_1290),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1333),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1325),
.A2(n_1331),
.B(n_1322),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1257),
.B(n_1279),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1365),
.A2(n_1372),
.B(n_1366),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1293),
.A2(n_1288),
.B(n_1309),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1261),
.B(n_1277),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1317),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1313),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1327),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1328),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1332),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1323),
.B(n_1358),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1348),
.Y(n_1393)
);

AO21x2_ASAP7_75t_L g1394 ( 
.A1(n_1343),
.A2(n_1329),
.B(n_1301),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1357),
.B(n_1248),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1326),
.Y(n_1396)
);

OAI211xp5_ASAP7_75t_L g1397 ( 
.A1(n_1260),
.A2(n_1366),
.B(n_1365),
.C(n_1372),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1288),
.B(n_1283),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1325),
.A2(n_1331),
.B(n_1322),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1333),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1348),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1334),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1334),
.Y(n_1403)
);

AO21x1_ASAP7_75t_SL g1404 ( 
.A1(n_1266),
.A2(n_1342),
.B(n_1295),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1283),
.B(n_1280),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1284),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1335),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1338),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1270),
.A2(n_1375),
.B1(n_1260),
.B2(n_1264),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1277),
.B(n_1360),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1335),
.Y(n_1411)
);

INVx8_ASAP7_75t_L g1412 ( 
.A(n_1284),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1292),
.B(n_1350),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1280),
.B(n_1266),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1270),
.A2(n_1375),
.B1(n_1264),
.B2(n_1274),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1281),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1339),
.Y(n_1417)
);

OR2x6_ASAP7_75t_L g1418 ( 
.A(n_1306),
.B(n_1352),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1368),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1319),
.A2(n_1309),
.B(n_1320),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1341),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1319),
.A2(n_1295),
.B(n_1311),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1278),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1282),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1311),
.A2(n_1272),
.B(n_1291),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1363),
.A2(n_1287),
.B1(n_1368),
.B2(n_1272),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1285),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1304),
.A2(n_1316),
.B(n_1299),
.Y(n_1428)
);

INVx4_ASAP7_75t_L g1429 ( 
.A(n_1286),
.Y(n_1429)
);

NAND2x1_ASAP7_75t_L g1430 ( 
.A(n_1298),
.B(n_1289),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1276),
.A2(n_1362),
.B(n_1346),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1267),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1251),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1347),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1370),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1371),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1352),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1340),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1318),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1273),
.B(n_1374),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1355),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1330),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1276),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1358),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1250),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1355),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1298),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1297),
.A2(n_1269),
.B(n_1258),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1275),
.A2(n_1345),
.B1(n_1356),
.B2(n_1361),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1303),
.B(n_1361),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1349),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1315),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1255),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1349),
.B(n_1356),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1376),
.B(n_1296),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1296),
.B(n_1310),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1271),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1296),
.B(n_1268),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1307),
.Y(n_1459)
);

OAI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1308),
.A2(n_1256),
.B(n_1302),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1305),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1305),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1376),
.B(n_1374),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1321),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1391),
.B(n_1359),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1384),
.A2(n_1359),
.B1(n_1249),
.B2(n_1252),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1413),
.B(n_1256),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1432),
.B(n_1456),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1423),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1417),
.B(n_1364),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1424),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1380),
.B(n_1344),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1408),
.B(n_1253),
.Y(n_1473)
);

AOI221xp5_ASAP7_75t_L g1474 ( 
.A1(n_1397),
.A2(n_1300),
.B1(n_1247),
.B2(n_1354),
.C(n_1265),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1408),
.B(n_1247),
.Y(n_1475)
);

BUFx12f_ASAP7_75t_SL g1476 ( 
.A(n_1463),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1391),
.B(n_1294),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1456),
.B(n_1324),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1451),
.B(n_1314),
.Y(n_1479)
);

AND2x2_ASAP7_75t_SL g1480 ( 
.A(n_1425),
.B(n_1422),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1386),
.B(n_1321),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1451),
.B(n_1259),
.Y(n_1482)
);

AOI221xp5_ASAP7_75t_L g1483 ( 
.A1(n_1409),
.A2(n_1263),
.B1(n_1415),
.B2(n_1385),
.C(n_1443),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1410),
.B(n_1434),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1449),
.A2(n_1426),
.B1(n_1395),
.B2(n_1383),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1414),
.A2(n_1398),
.B(n_1443),
.C(n_1420),
.Y(n_1486)
);

AOI221xp5_ASAP7_75t_L g1487 ( 
.A1(n_1398),
.A2(n_1379),
.B1(n_1405),
.B2(n_1442),
.C(n_1438),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1417),
.B(n_1421),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1421),
.B(n_1392),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1382),
.A2(n_1399),
.B(n_1442),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1392),
.B(n_1446),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1396),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1454),
.B(n_1450),
.Y(n_1494)
);

A2O1A1Ixp33_ASAP7_75t_L g1495 ( 
.A1(n_1414),
.A2(n_1420),
.B(n_1405),
.C(n_1399),
.Y(n_1495)
);

AOI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1379),
.A2(n_1438),
.B1(n_1445),
.B2(n_1439),
.C(n_1419),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_SL g1497 ( 
.A(n_1396),
.Y(n_1497)
);

NAND3xp33_ASAP7_75t_L g1498 ( 
.A(n_1425),
.B(n_1439),
.C(n_1448),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1423),
.B(n_1379),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1450),
.B(n_1411),
.Y(n_1500)
);

O2A1O1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1461),
.A2(n_1462),
.B(n_1440),
.C(n_1411),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1392),
.Y(n_1502)
);

AO32x1_ASAP7_75t_L g1503 ( 
.A1(n_1377),
.A2(n_1378),
.A3(n_1390),
.B1(n_1389),
.B2(n_1403),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1431),
.Y(n_1504)
);

O2A1O1Ixp33_ASAP7_75t_L g1505 ( 
.A1(n_1461),
.A2(n_1462),
.B(n_1425),
.C(n_1464),
.Y(n_1505)
);

OA21x2_ASAP7_75t_L g1506 ( 
.A1(n_1387),
.A2(n_1378),
.B(n_1402),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1431),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1452),
.Y(n_1508)
);

OR2x6_ASAP7_75t_L g1509 ( 
.A(n_1418),
.B(n_1412),
.Y(n_1509)
);

AOI221xp5_ASAP7_75t_L g1510 ( 
.A1(n_1436),
.A2(n_1427),
.B1(n_1452),
.B2(n_1390),
.C(n_1389),
.Y(n_1510)
);

OR2x6_ASAP7_75t_L g1511 ( 
.A(n_1418),
.B(n_1412),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1433),
.B(n_1435),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1460),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1444),
.B(n_1396),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1381),
.B(n_1400),
.Y(n_1515)
);

OAI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1425),
.A2(n_1447),
.B(n_1430),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1416),
.B(n_1435),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1444),
.B(n_1459),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1464),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1422),
.A2(n_1428),
.B(n_1418),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1446),
.B(n_1418),
.Y(n_1521)
);

O2A1O1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1464),
.A2(n_1447),
.B(n_1455),
.C(n_1457),
.Y(n_1522)
);

A2O1A1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1381),
.A2(n_1400),
.B(n_1407),
.C(n_1404),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1431),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1407),
.B(n_1429),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1506),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1484),
.B(n_1393),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1506),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1496),
.B(n_1437),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1469),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1480),
.B(n_1422),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1469),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1502),
.B(n_1388),
.Y(n_1533)
);

INVx2_ASAP7_75t_SL g1534 ( 
.A(n_1502),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1480),
.B(n_1422),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1499),
.B(n_1394),
.Y(n_1536)
);

OAI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1483),
.A2(n_1430),
.B1(n_1441),
.B2(n_1457),
.C(n_1453),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1504),
.B(n_1393),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1499),
.B(n_1394),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1471),
.Y(n_1540)
);

NAND2x1p5_ASAP7_75t_L g1541 ( 
.A(n_1520),
.B(n_1431),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1490),
.B(n_1394),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1521),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1485),
.A2(n_1404),
.B1(n_1458),
.B2(n_1428),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1507),
.B(n_1401),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1495),
.B(n_1403),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1517),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1495),
.B(n_1402),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1524),
.B(n_1401),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1503),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1472),
.A2(n_1458),
.B1(n_1428),
.B2(n_1436),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1500),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1512),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1552),
.B(n_1494),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1538),
.Y(n_1555)
);

AOI221xp5_ASAP7_75t_L g1556 ( 
.A1(n_1529),
.A2(n_1487),
.B1(n_1498),
.B2(n_1472),
.C(n_1466),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1538),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1540),
.B(n_1486),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1543),
.Y(n_1559)
);

INVx4_ASAP7_75t_L g1560 ( 
.A(n_1533),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1538),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1545),
.Y(n_1562)
);

NAND3xp33_ASAP7_75t_L g1563 ( 
.A(n_1529),
.B(n_1466),
.C(n_1544),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1531),
.B(n_1535),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1528),
.Y(n_1565)
);

NAND4xp25_ASAP7_75t_L g1566 ( 
.A(n_1551),
.B(n_1474),
.C(n_1501),
.D(n_1505),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1540),
.B(n_1486),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1531),
.B(n_1491),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1531),
.B(n_1493),
.Y(n_1569)
);

OAI33xp33_ASAP7_75t_L g1570 ( 
.A1(n_1527),
.A2(n_1508),
.A3(n_1467),
.B1(n_1481),
.B2(n_1477),
.B3(n_1522),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1534),
.Y(n_1571)
);

INVxp67_ASAP7_75t_L g1572 ( 
.A(n_1527),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1547),
.B(n_1549),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1552),
.B(n_1553),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1535),
.B(n_1521),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_R g1576 ( 
.A(n_1544),
.B(n_1513),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1537),
.B(n_1473),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1528),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1535),
.B(n_1521),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1530),
.Y(n_1580)
);

AOI33xp33_ASAP7_75t_L g1581 ( 
.A1(n_1551),
.A2(n_1465),
.A3(n_1510),
.B1(n_1468),
.B2(n_1514),
.B3(n_1518),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1530),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1530),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1532),
.Y(n_1584)
);

NAND2xp33_ASAP7_75t_SL g1585 ( 
.A(n_1546),
.B(n_1513),
.Y(n_1585)
);

AOI211xp5_ASAP7_75t_L g1586 ( 
.A1(n_1537),
.A2(n_1523),
.B(n_1488),
.C(n_1515),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1580),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1573),
.B(n_1555),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1572),
.B(n_1553),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1564),
.B(n_1536),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1559),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1580),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1582),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1578),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1560),
.B(n_1528),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1582),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1564),
.B(n_1536),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1583),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1583),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1584),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1578),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1584),
.Y(n_1602)
);

NOR3xp33_ASAP7_75t_L g1603 ( 
.A(n_1563),
.B(n_1488),
.C(n_1475),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1560),
.B(n_1536),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1573),
.B(n_1550),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1555),
.B(n_1550),
.Y(n_1606)
);

NOR2xp67_ASAP7_75t_L g1607 ( 
.A(n_1560),
.B(n_1526),
.Y(n_1607)
);

AND2x2_ASAP7_75t_SL g1608 ( 
.A(n_1556),
.B(n_1546),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1560),
.B(n_1539),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1557),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1578),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1557),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1561),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1561),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1565),
.Y(n_1615)
);

INVxp67_ASAP7_75t_SL g1616 ( 
.A(n_1558),
.Y(n_1616)
);

INVx4_ASAP7_75t_L g1617 ( 
.A(n_1559),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1571),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1574),
.B(n_1553),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1565),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1587),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1590),
.B(n_1597),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1616),
.B(n_1558),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1591),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1587),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1608),
.B(n_1577),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1590),
.B(n_1597),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1608),
.B(n_1581),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1592),
.Y(n_1629)
);

OR2x2_ASAP7_75t_SL g1630 ( 
.A(n_1608),
.B(n_1563),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1592),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1593),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1616),
.B(n_1567),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1593),
.Y(n_1634)
);

AOI21xp33_ASAP7_75t_L g1635 ( 
.A1(n_1608),
.A2(n_1567),
.B(n_1586),
.Y(n_1635)
);

AND3x1_ASAP7_75t_L g1636 ( 
.A(n_1603),
.B(n_1586),
.C(n_1515),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1588),
.B(n_1610),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1596),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1596),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1598),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1603),
.B(n_1569),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1598),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1599),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1619),
.B(n_1569),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1591),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1588),
.B(n_1562),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1590),
.B(n_1575),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1619),
.B(n_1554),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1606),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1599),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1600),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1589),
.B(n_1585),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1589),
.B(n_1570),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1597),
.B(n_1575),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1604),
.B(n_1579),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1600),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1606),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1602),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1588),
.B(n_1470),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1604),
.B(n_1579),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1617),
.B(n_1562),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1606),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1623),
.B(n_1605),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1626),
.B(n_1659),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1645),
.Y(n_1665)
);

AOI211xp5_ASAP7_75t_L g1666 ( 
.A1(n_1635),
.A2(n_1566),
.B(n_1576),
.C(n_1523),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1625),
.Y(n_1667)
);

AND2x2_ASAP7_75t_SL g1668 ( 
.A(n_1636),
.B(n_1617),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1647),
.B(n_1617),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1645),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1647),
.B(n_1617),
.Y(n_1671)
);

AND3x2_ASAP7_75t_L g1672 ( 
.A(n_1624),
.B(n_1618),
.C(n_1470),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1653),
.B(n_1610),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1622),
.B(n_1617),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1628),
.A2(n_1470),
.B(n_1618),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1622),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_SL g1677 ( 
.A(n_1652),
.B(n_1641),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1648),
.B(n_1612),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1623),
.B(n_1612),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1627),
.B(n_1604),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1627),
.B(n_1609),
.Y(n_1681)
);

OAI21xp33_ASAP7_75t_SL g1682 ( 
.A1(n_1630),
.A2(n_1607),
.B(n_1609),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1633),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1655),
.B(n_1609),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1633),
.B(n_1613),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1637),
.B(n_1605),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1630),
.Y(n_1687)
);

NAND4xp25_ASAP7_75t_SL g1688 ( 
.A(n_1654),
.B(n_1482),
.C(n_1478),
.D(n_1605),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1637),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1621),
.B(n_1613),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1625),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1642),
.B(n_1614),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1644),
.B(n_1497),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1643),
.B(n_1614),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1661),
.A2(n_1511),
.B1(n_1509),
.B2(n_1489),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1656),
.B(n_1602),
.Y(n_1696)
);

INVx2_ASAP7_75t_SL g1697 ( 
.A(n_1661),
.Y(n_1697)
);

NAND2x1_ASAP7_75t_L g1698 ( 
.A(n_1676),
.B(n_1661),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1665),
.Y(n_1699)
);

OAI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1687),
.A2(n_1542),
.B(n_1607),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1687),
.B(n_1673),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1687),
.B(n_1655),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1677),
.A2(n_1658),
.B(n_1629),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1670),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1670),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1666),
.A2(n_1519),
.B1(n_1541),
.B2(n_1550),
.Y(n_1706)
);

OAI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1666),
.A2(n_1638),
.B1(n_1631),
.B2(n_1632),
.C(n_1651),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_SL g1708 ( 
.A(n_1668),
.B(n_1672),
.Y(n_1708)
);

AOI311xp33_ASAP7_75t_L g1709 ( 
.A1(n_1673),
.A2(n_1629),
.A3(n_1638),
.B(n_1639),
.C(n_1640),
.Y(n_1709)
);

OAI22xp33_ASAP7_75t_SL g1710 ( 
.A1(n_1675),
.A2(n_1646),
.B1(n_1657),
.B2(n_1662),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1668),
.A2(n_1548),
.B1(n_1546),
.B2(n_1660),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1664),
.B(n_1660),
.Y(n_1712)
);

OAI21xp33_ASAP7_75t_L g1713 ( 
.A1(n_1668),
.A2(n_1683),
.B(n_1682),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1670),
.B(n_1631),
.Y(n_1714)
);

INVxp67_ASAP7_75t_SL g1715 ( 
.A(n_1676),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1689),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1667),
.Y(n_1717)
);

OA21x2_ASAP7_75t_L g1718 ( 
.A1(n_1667),
.A2(n_1662),
.B(n_1657),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1697),
.B(n_1649),
.Y(n_1719)
);

OAI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1676),
.A2(n_1492),
.B1(n_1646),
.B2(n_1511),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1676),
.B(n_1568),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1688),
.B(n_1519),
.Y(n_1722)
);

OAI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1708),
.A2(n_1697),
.B1(n_1689),
.B2(n_1663),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1710),
.B(n_1682),
.Y(n_1724)
);

OAI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1711),
.A2(n_1663),
.B1(n_1686),
.B2(n_1685),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1715),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_1698),
.Y(n_1727)
);

AOI322xp5_ASAP7_75t_L g1728 ( 
.A1(n_1713),
.A2(n_1680),
.A3(n_1681),
.B1(n_1684),
.B2(n_1669),
.C1(n_1671),
.C2(n_1674),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1702),
.B(n_1669),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1719),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1704),
.Y(n_1731)
);

O2A1O1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1701),
.A2(n_1679),
.B(n_1685),
.C(n_1678),
.Y(n_1732)
);

NOR3xp33_ASAP7_75t_L g1733 ( 
.A(n_1707),
.B(n_1693),
.C(n_1691),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1716),
.B(n_1671),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1705),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1712),
.B(n_1678),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1699),
.B(n_1674),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1718),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1718),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1714),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1714),
.B(n_1686),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1730),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1734),
.B(n_1703),
.Y(n_1743)
);

AOI21xp33_ASAP7_75t_SL g1744 ( 
.A1(n_1723),
.A2(n_1706),
.B(n_1722),
.Y(n_1744)
);

AOI221xp5_ASAP7_75t_L g1745 ( 
.A1(n_1724),
.A2(n_1706),
.B1(n_1700),
.B2(n_1717),
.C(n_1720),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1725),
.A2(n_1732),
.B(n_1727),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1726),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1727),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1734),
.B(n_1719),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1726),
.Y(n_1750)
);

NAND2x1p5_ASAP7_75t_L g1751 ( 
.A(n_1737),
.B(n_1492),
.Y(n_1751)
);

INVxp67_ASAP7_75t_L g1752 ( 
.A(n_1737),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1733),
.A2(n_1721),
.B1(n_1700),
.B2(n_1695),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1748),
.B(n_1729),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1753),
.A2(n_1739),
.B1(n_1736),
.B2(n_1729),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1742),
.B(n_1728),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_SL g1757 ( 
.A(n_1743),
.B(n_1741),
.Y(n_1757)
);

NAND4xp25_ASAP7_75t_L g1758 ( 
.A(n_1746),
.B(n_1709),
.C(n_1740),
.D(n_1735),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1745),
.A2(n_1739),
.B(n_1738),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1752),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1747),
.Y(n_1761)
);

OAI221xp5_ASAP7_75t_L g1762 ( 
.A1(n_1744),
.A2(n_1741),
.B1(n_1739),
.B2(n_1738),
.C(n_1740),
.Y(n_1762)
);

NAND2xp33_ASAP7_75t_R g1763 ( 
.A(n_1749),
.B(n_1731),
.Y(n_1763)
);

AOI221xp5_ASAP7_75t_SL g1764 ( 
.A1(n_1759),
.A2(n_1744),
.B1(n_1762),
.B2(n_1758),
.C(n_1755),
.Y(n_1764)
);

AOI222xp33_ASAP7_75t_L g1765 ( 
.A1(n_1757),
.A2(n_1750),
.B1(n_1735),
.B2(n_1731),
.C1(n_1691),
.C2(n_1694),
.Y(n_1765)
);

NAND3xp33_ASAP7_75t_L g1766 ( 
.A(n_1763),
.B(n_1756),
.C(n_1754),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1760),
.A2(n_1751),
.B(n_1694),
.Y(n_1767)
);

O2A1O1Ixp33_ASAP7_75t_L g1768 ( 
.A1(n_1761),
.A2(n_1692),
.B(n_1690),
.C(n_1696),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1764),
.A2(n_1681),
.B1(n_1680),
.B2(n_1684),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1766),
.Y(n_1770)
);

AOI222xp33_ASAP7_75t_L g1771 ( 
.A1(n_1765),
.A2(n_1692),
.B1(n_1690),
.B2(n_1696),
.C1(n_1649),
.C2(n_1650),
.Y(n_1771)
);

AOI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1767),
.A2(n_1492),
.B1(n_1650),
.B2(n_1640),
.Y(n_1772)
);

OAI211xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1768),
.A2(n_1651),
.B(n_1639),
.C(n_1634),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1768),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1769),
.B(n_1634),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1770),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1774),
.B(n_1632),
.Y(n_1777)
);

OAI211xp5_ASAP7_75t_SL g1778 ( 
.A1(n_1772),
.A2(n_1500),
.B(n_1525),
.C(n_1516),
.Y(n_1778)
);

NOR2x1p5_ASAP7_75t_L g1779 ( 
.A(n_1773),
.B(n_1492),
.Y(n_1779)
);

OAI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1775),
.A2(n_1771),
.B(n_1595),
.Y(n_1780)
);

NAND4xp25_ASAP7_75t_L g1781 ( 
.A(n_1777),
.B(n_1525),
.C(n_1479),
.D(n_1465),
.Y(n_1781)
);

OAI321xp33_ASAP7_75t_L g1782 ( 
.A1(n_1778),
.A2(n_1541),
.A3(n_1509),
.B1(n_1511),
.B2(n_1453),
.C(n_1548),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1780),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1783),
.A2(n_1776),
.B1(n_1779),
.B2(n_1781),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1784),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1785),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1786),
.Y(n_1787)
);

OA21x2_ASAP7_75t_L g1788 ( 
.A1(n_1787),
.A2(n_1782),
.B(n_1601),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1788),
.A2(n_1611),
.B(n_1594),
.Y(n_1789)
);

AO21x2_ASAP7_75t_L g1790 ( 
.A1(n_1789),
.A2(n_1611),
.B(n_1594),
.Y(n_1790)
);

OAI222xp33_ASAP7_75t_L g1791 ( 
.A1(n_1789),
.A2(n_1611),
.B1(n_1601),
.B2(n_1594),
.C1(n_1615),
.C2(n_1620),
.Y(n_1791)
);

OAI221xp5_ASAP7_75t_R g1792 ( 
.A1(n_1790),
.A2(n_1412),
.B1(n_1601),
.B2(n_1476),
.C(n_1615),
.Y(n_1792)
);

AOI211xp5_ASAP7_75t_L g1793 ( 
.A1(n_1792),
.A2(n_1791),
.B(n_1406),
.C(n_1458),
.Y(n_1793)
);


endmodule