module real_aes_2948_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_741;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_0), .B(n_113), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_1), .A2(n_122), .B(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_2), .B(n_760), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_3), .B(n_113), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_4), .B(n_129), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_5), .B(n_129), .Y(n_498) );
INVx1_ASAP7_75t_L g120 ( .A(n_6), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_7), .B(n_129), .Y(n_469) );
CKINVDCx16_ASAP7_75t_R g760 ( .A(n_8), .Y(n_760) );
NAND2xp33_ASAP7_75t_L g479 ( .A(n_9), .B(n_131), .Y(n_479) );
AND2x2_ASAP7_75t_L g149 ( .A(n_10), .B(n_138), .Y(n_149) );
AND2x2_ASAP7_75t_L g158 ( .A(n_11), .B(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g135 ( .A(n_12), .Y(n_135) );
AOI221x1_ASAP7_75t_L g520 ( .A1(n_13), .A2(n_24), .B1(n_113), .B2(n_122), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_14), .B(n_129), .Y(n_168) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_15), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_16), .B(n_113), .Y(n_475) );
AO21x2_ASAP7_75t_L g473 ( .A1(n_17), .A2(n_138), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_18), .B(n_133), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_19), .B(n_129), .Y(n_458) );
AO21x1_ASAP7_75t_L g493 ( .A1(n_20), .A2(n_113), .B(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_21), .B(n_113), .Y(n_183) );
INVx1_ASAP7_75t_L g444 ( .A(n_22), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_23), .A2(n_89), .B1(n_113), .B2(n_222), .Y(n_221) );
NAND2x1_ASAP7_75t_L g507 ( .A(n_25), .B(n_129), .Y(n_507) );
NAND2x1_ASAP7_75t_L g468 ( .A(n_26), .B(n_131), .Y(n_468) );
OR2x2_ASAP7_75t_L g136 ( .A(n_27), .B(n_86), .Y(n_136) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_27), .A2(n_86), .B(n_135), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_28), .B(n_131), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_29), .B(n_129), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_30), .Y(n_779) );
AO21x2_ASAP7_75t_L g163 ( .A1(n_31), .A2(n_159), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_32), .B(n_131), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_33), .A2(n_122), .B(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_34), .B(n_129), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_35), .A2(n_122), .B(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g119 ( .A(n_36), .B(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g123 ( .A(n_36), .B(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g230 ( .A(n_36), .Y(n_230) );
OR2x6_ASAP7_75t_L g442 ( .A(n_37), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_38), .B(n_113), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_39), .B(n_113), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_40), .B(n_129), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_41), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_42), .B(n_131), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_43), .B(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_44), .A2(n_122), .B(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_45), .A2(n_122), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_46), .B(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_47), .B(n_131), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_48), .B(n_113), .Y(n_165) );
INVx1_ASAP7_75t_L g116 ( .A(n_49), .Y(n_116) );
INVx1_ASAP7_75t_L g126 ( .A(n_49), .Y(n_126) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_50), .A2(n_66), .B1(n_769), .B2(n_770), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_50), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_51), .B(n_129), .Y(n_156) );
AND2x2_ASAP7_75t_L g194 ( .A(n_52), .B(n_133), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_53), .B(n_131), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_54), .B(n_129), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_55), .B(n_131), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_56), .A2(n_122), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_57), .B(n_113), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_58), .B(n_113), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_59), .A2(n_122), .B(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g189 ( .A(n_60), .B(n_134), .Y(n_189) );
AO21x1_ASAP7_75t_L g495 ( .A1(n_61), .A2(n_122), .B(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_62), .B(n_113), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_63), .A2(n_80), .B1(n_742), .B2(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_63), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_64), .B(n_131), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_65), .B(n_113), .Y(n_470) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_66), .A2(n_101), .B1(n_753), .B2(n_764), .C1(n_780), .C2(n_784), .Y(n_100) );
INVx1_ASAP7_75t_L g770 ( .A(n_66), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_67), .B(n_131), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_68), .A2(n_94), .B1(n_122), .B2(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_69), .B(n_129), .Y(n_186) );
AND2x2_ASAP7_75t_L g543 ( .A(n_70), .B(n_134), .Y(n_543) );
INVx1_ASAP7_75t_L g118 ( .A(n_71), .Y(n_118) );
INVx1_ASAP7_75t_L g124 ( .A(n_71), .Y(n_124) );
AND2x2_ASAP7_75t_L g471 ( .A(n_72), .B(n_159), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_73), .B(n_131), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_74), .A2(n_122), .B(n_198), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_75), .A2(n_122), .B(n_127), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_76), .A2(n_122), .B(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g180 ( .A(n_77), .B(n_134), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_78), .B(n_133), .Y(n_219) );
INVx1_ASAP7_75t_L g445 ( .A(n_79), .Y(n_445) );
INVx1_ASAP7_75t_L g743 ( .A(n_80), .Y(n_743) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_81), .B(n_113), .Y(n_460) );
AND2x2_ASAP7_75t_L g481 ( .A(n_82), .B(n_159), .Y(n_481) );
AOI22xp33_ASAP7_75t_SL g744 ( .A1(n_83), .A2(n_741), .B1(n_745), .B2(n_749), .Y(n_744) );
AND2x2_ASAP7_75t_L g137 ( .A(n_84), .B(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g494 ( .A(n_85), .B(n_170), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_87), .B(n_131), .Y(n_459) );
AND2x2_ASAP7_75t_L g510 ( .A(n_88), .B(n_159), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_90), .B(n_129), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_91), .A2(n_122), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_92), .B(n_131), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_93), .A2(n_122), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_95), .B(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_96), .B(n_129), .Y(n_486) );
BUFx2_ASAP7_75t_L g188 ( .A(n_97), .Y(n_188) );
BUFx2_ASAP7_75t_L g761 ( .A(n_98), .Y(n_761) );
BUFx2_ASAP7_75t_SL g790 ( .A(n_98), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_99), .A2(n_122), .B(n_477), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_741), .B(n_744), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_439), .B1(n_446), .B2(n_737), .Y(n_103) );
INVx1_ASAP7_75t_L g746 ( .A(n_104), .Y(n_746) );
OAI22xp5_ASAP7_75t_SL g766 ( .A1(n_104), .A2(n_767), .B1(n_768), .B2(n_771), .Y(n_766) );
INVx5_ASAP7_75t_L g767 ( .A(n_104), .Y(n_767) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_343), .Y(n_104) );
NOR3xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_268), .C(n_304), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_242), .Y(n_106) );
AOI211xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_160), .B(n_190), .C(n_215), .Y(n_107) );
AND2x2_ASAP7_75t_L g333 ( .A(n_108), .B(n_192), .Y(n_333) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_140), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_109), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g366 ( .A(n_109), .B(n_248), .Y(n_366) );
AND2x2_ASAP7_75t_L g382 ( .A(n_109), .B(n_207), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_109), .B(n_392), .Y(n_391) );
NAND2x1p5_ASAP7_75t_L g415 ( .A(n_109), .B(n_416), .Y(n_415) );
INVx4_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x4_ASAP7_75t_SL g202 ( .A(n_110), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g237 ( .A(n_110), .Y(n_237) );
AND2x2_ASAP7_75t_L g284 ( .A(n_110), .B(n_217), .Y(n_284) );
AND2x2_ASAP7_75t_L g303 ( .A(n_110), .B(n_140), .Y(n_303) );
BUFx2_ASAP7_75t_L g308 ( .A(n_110), .Y(n_308) );
AND2x2_ASAP7_75t_L g352 ( .A(n_110), .B(n_150), .Y(n_352) );
AND2x4_ASAP7_75t_L g424 ( .A(n_110), .B(n_425), .Y(n_424) );
NOR2x1_ASAP7_75t_L g436 ( .A(n_110), .B(n_206), .Y(n_436) );
OR2x6_ASAP7_75t_L g110 ( .A(n_111), .B(n_137), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_121), .B(n_133), .Y(n_111) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_119), .Y(n_113) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
AND2x6_ASAP7_75t_L g131 ( .A(n_115), .B(n_124), .Y(n_131) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g129 ( .A(n_117), .B(n_126), .Y(n_129) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx5_ASAP7_75t_L g132 ( .A(n_119), .Y(n_132) );
AND2x2_ASAP7_75t_L g125 ( .A(n_120), .B(n_126), .Y(n_125) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_120), .Y(n_225) );
AND2x6_ASAP7_75t_L g122 ( .A(n_123), .B(n_125), .Y(n_122) );
BUFx3_ASAP7_75t_L g226 ( .A(n_123), .Y(n_226) );
INVx2_ASAP7_75t_L g232 ( .A(n_124), .Y(n_232) );
AND2x4_ASAP7_75t_L g228 ( .A(n_125), .B(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g224 ( .A(n_126), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_130), .B(n_132), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_131), .B(n_188), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_132), .A2(n_146), .B(n_147), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_132), .A2(n_155), .B(n_156), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_132), .A2(n_168), .B(n_169), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_132), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_132), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_132), .A2(n_199), .B(n_200), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_132), .A2(n_458), .B(n_459), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_132), .A2(n_468), .B(n_469), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_132), .A2(n_478), .B(n_479), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_132), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_132), .A2(n_497), .B(n_498), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_132), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_132), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_132), .A2(n_540), .B(n_541), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_133), .Y(n_142) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_133), .A2(n_221), .B(n_227), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_133), .A2(n_483), .B(n_484), .Y(n_482) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_133), .A2(n_520), .B(n_524), .Y(n_519) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_133), .A2(n_520), .B(n_524), .Y(n_531) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_SL g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x4_ASAP7_75t_L g170 ( .A(n_135), .B(n_136), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_138), .A2(n_183), .B(n_184), .Y(n_182) );
BUFx4f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx3_ASAP7_75t_L g151 ( .A(n_139), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_140), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g355 ( .A(n_140), .Y(n_355) );
BUFx2_ASAP7_75t_L g404 ( .A(n_140), .Y(n_404) );
INVx1_ASAP7_75t_L g426 ( .A(n_140), .Y(n_426) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_150), .Y(n_140) );
INVx3_ASAP7_75t_L g203 ( .A(n_141), .Y(n_203) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_141), .Y(n_392) );
AOI21x1_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_149), .Y(n_141) );
AO21x2_ASAP7_75t_L g464 ( .A1(n_142), .A2(n_465), .B(n_471), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
INVx2_ASAP7_75t_L g206 ( .A(n_150), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_150), .B(n_203), .Y(n_207) );
INVx2_ASAP7_75t_L g292 ( .A(n_150), .Y(n_292) );
OR2x2_ASAP7_75t_L g299 ( .A(n_150), .B(n_248), .Y(n_299) );
AO21x2_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_158), .Y(n_150) );
INVx4_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_157), .Y(n_152) );
INVx3_ASAP7_75t_L g173 ( .A(n_159), .Y(n_173) );
AND2x2_ASAP7_75t_L g254 ( .A(n_160), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g288 ( .A(n_160), .B(n_251), .Y(n_288) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_171), .Y(n_160) );
AND2x2_ASAP7_75t_L g324 ( .A(n_161), .B(n_213), .Y(n_324) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g281 ( .A(n_162), .B(n_172), .Y(n_281) );
AND2x2_ASAP7_75t_L g400 ( .A(n_162), .B(n_181), .Y(n_400) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g212 ( .A(n_163), .Y(n_212) );
INVx1_ASAP7_75t_L g240 ( .A(n_163), .Y(n_240) );
AND2x2_ASAP7_75t_L g296 ( .A(n_163), .B(n_172), .Y(n_296) );
AND2x2_ASAP7_75t_L g301 ( .A(n_163), .B(n_193), .Y(n_301) );
OR2x2_ASAP7_75t_L g364 ( .A(n_163), .B(n_181), .Y(n_364) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_163), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_170), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_170), .A2(n_196), .B(n_197), .Y(n_195) );
INVx1_ASAP7_75t_SL g454 ( .A(n_170), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_170), .A2(n_475), .B(n_476), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_170), .B(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g192 ( .A(n_171), .B(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g241 ( .A(n_171), .Y(n_241) );
NOR2x1_ASAP7_75t_SL g171 ( .A(n_172), .B(n_181), .Y(n_171) );
AO21x1_ASAP7_75t_SL g172 ( .A1(n_173), .A2(n_174), .B(n_180), .Y(n_172) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_173), .A2(n_174), .B(n_180), .Y(n_214) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_173), .A2(n_504), .B(n_510), .Y(n_503) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_173), .A2(n_537), .B(n_543), .Y(n_536) );
AO21x2_ASAP7_75t_L g572 ( .A1(n_173), .A2(n_537), .B(n_543), .Y(n_572) );
AO21x2_ASAP7_75t_L g575 ( .A1(n_173), .A2(n_504), .B(n_510), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_179), .Y(n_174) );
AND2x2_ASAP7_75t_L g209 ( .A(n_181), .B(n_210), .Y(n_209) );
INVx2_ASAP7_75t_SL g267 ( .A(n_181), .Y(n_267) );
NAND2x1_ASAP7_75t_L g277 ( .A(n_181), .B(n_193), .Y(n_277) );
OR2x2_ASAP7_75t_L g282 ( .A(n_181), .B(n_210), .Y(n_282) );
BUFx2_ASAP7_75t_L g338 ( .A(n_181), .Y(n_338) );
AND2x2_ASAP7_75t_L g374 ( .A(n_181), .B(n_253), .Y(n_374) );
AND2x2_ASAP7_75t_L g385 ( .A(n_181), .B(n_213), .Y(n_385) );
OR2x6_ASAP7_75t_L g181 ( .A(n_182), .B(n_189), .Y(n_181) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_201), .B1(n_207), .B2(n_208), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_192), .A2(n_382), .B1(n_432), .B2(n_437), .Y(n_431) );
INVx4_ASAP7_75t_L g210 ( .A(n_193), .Y(n_210) );
INVx2_ASAP7_75t_L g251 ( .A(n_193), .Y(n_251) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_193), .Y(n_322) );
OR2x2_ASAP7_75t_L g337 ( .A(n_193), .B(n_213), .Y(n_337) );
OR2x2_ASAP7_75t_SL g363 ( .A(n_193), .B(n_364), .Y(n_363) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_202), .B(n_204), .Y(n_201) );
INVx2_ASAP7_75t_SL g244 ( .A(n_202), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_202), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g312 ( .A(n_202), .B(n_260), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_202), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g234 ( .A(n_203), .Y(n_234) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_203), .Y(n_259) );
AND2x2_ASAP7_75t_L g315 ( .A(n_203), .B(n_292), .Y(n_315) );
INVx1_ASAP7_75t_L g425 ( .A(n_203), .Y(n_425) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_205), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_205), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g233 ( .A(n_206), .B(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_207), .B(n_366), .Y(n_365) );
AOI321xp33_ASAP7_75t_L g387 ( .A1(n_208), .A2(n_289), .A3(n_357), .B1(n_388), .B2(n_389), .C(n_393), .Y(n_387) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_211), .Y(n_208) );
INVxp67_ASAP7_75t_SL g286 ( .A(n_209), .Y(n_286) );
AND2x2_ASAP7_75t_L g311 ( .A(n_209), .B(n_240), .Y(n_311) );
AND2x2_ASAP7_75t_L g386 ( .A(n_209), .B(n_296), .Y(n_386) );
INVx1_ASAP7_75t_L g255 ( .A(n_210), .Y(n_255) );
BUFx2_ASAP7_75t_L g265 ( .A(n_210), .Y(n_265) );
NOR2xp67_ASAP7_75t_L g372 ( .A(n_210), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g310 ( .A(n_211), .Y(n_310) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
BUFx2_ASAP7_75t_L g317 ( .A(n_212), .Y(n_317) );
INVx2_ASAP7_75t_L g253 ( .A(n_213), .Y(n_253) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_213), .Y(n_276) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AOI21xp33_ASAP7_75t_SL g215 ( .A1(n_216), .A2(n_235), .B(n_238), .Y(n_215) );
NOR2xp67_ASAP7_75t_L g369 ( .A(n_216), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_233), .Y(n_217) );
INVx3_ASAP7_75t_L g260 ( .A(n_218), .Y(n_260) );
AND2x2_ASAP7_75t_L g291 ( .A(n_218), .B(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
AND2x4_ASAP7_75t_L g248 ( .A(n_219), .B(n_220), .Y(n_248) );
AND2x4_ASAP7_75t_L g222 ( .A(n_223), .B(n_226), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
NOR2x1p5_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
INVx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g331 ( .A(n_233), .Y(n_331) );
INVx1_ASAP7_75t_SL g416 ( .A(n_234), .Y(n_416) );
INVxp33_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_237), .B(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g342 ( .A(n_237), .B(n_299), .Y(n_342) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_241), .Y(n_238) );
AND2x2_ASAP7_75t_L g346 ( .A(n_239), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_239), .B(n_361), .Y(n_360) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_240), .B(n_277), .Y(n_332) );
NOR4xp25_ASAP7_75t_L g427 ( .A(n_240), .B(n_271), .C(n_428), .D(n_429), .Y(n_427) );
OR2x2_ASAP7_75t_L g395 ( .A(n_241), .B(n_396), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_249), .B1(n_254), .B2(n_256), .C(n_261), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
AND2x2_ASAP7_75t_L g270 ( .A(n_245), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g307 ( .A(n_246), .B(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g327 ( .A(n_247), .Y(n_327) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
BUFx3_ASAP7_75t_L g350 ( .A(n_248), .Y(n_350) );
AND2x2_ASAP7_75t_L g357 ( .A(n_248), .B(n_358), .Y(n_357) );
INVxp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
OR2x2_ASAP7_75t_L g294 ( .A(n_251), .B(n_295), .Y(n_294) );
INVxp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_253), .B(n_267), .Y(n_266) );
INVxp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
INVx2_ASAP7_75t_L g271 ( .A(n_258), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_258), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g263 ( .A(n_260), .Y(n_263) );
OAI321xp33_ASAP7_75t_L g375 ( .A1(n_260), .A2(n_368), .A3(n_376), .B1(n_381), .B2(n_383), .C(n_387), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
OR2x2_ASAP7_75t_L g330 ( .A(n_263), .B(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_L g430 ( .A(n_266), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_267), .B(n_310), .Y(n_309) );
NAND2xp33_ASAP7_75t_SL g410 ( .A(n_267), .B(n_281), .Y(n_410) );
OAI211xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_272), .B(n_283), .C(n_287), .Y(n_268) );
INVxp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NOR2x1_ASAP7_75t_L g272 ( .A(n_273), .B(n_278), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g379 ( .A(n_276), .Y(n_379) );
INVx3_ASAP7_75t_L g318 ( .A(n_277), .Y(n_318) );
OR2x2_ASAP7_75t_L g421 ( .A(n_277), .B(n_295), .Y(n_421) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_279), .A2(n_363), .B1(n_365), .B2(n_367), .Y(n_362) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_SL g361 ( .A(n_282), .Y(n_361) );
OR2x2_ASAP7_75t_L g438 ( .A(n_282), .B(n_295), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AOI21xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_289), .B(n_293), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_291), .B(n_308), .Y(n_407) );
AND2x2_ASAP7_75t_L g413 ( .A(n_291), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g358 ( .A(n_292), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_297), .B1(n_300), .B2(n_302), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_L g339 ( .A1(n_295), .A2(n_338), .B(n_340), .C(n_342), .Y(n_339) );
INVx2_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_298), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_298), .B(n_390), .Y(n_412) );
INVx2_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g384 ( .A(n_301), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g334 ( .A1(n_303), .A2(n_335), .B(n_338), .C(n_339), .Y(n_334) );
NAND3xp33_ASAP7_75t_SL g304 ( .A(n_305), .B(n_319), .C(n_334), .Y(n_304) );
AOI222xp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_309), .B1(n_311), .B2(n_312), .C1(n_313), .C2(n_316), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g368 ( .A(n_308), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_308), .B(n_341), .Y(n_394) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_SL g328 ( .A(n_315), .Y(n_328) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
OR2x2_ASAP7_75t_L g433 ( .A(n_317), .B(n_350), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_318), .A2(n_409), .B1(n_411), .B2(n_413), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_325), .B1(n_329), .B2(n_332), .C(n_333), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI21xp5_ASAP7_75t_SL g393 ( .A1(n_326), .A2(n_394), .B(n_395), .Y(n_393) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx2_ASAP7_75t_L g341 ( .A(n_327), .Y(n_341) );
AND2x2_ASAP7_75t_L g435 ( .A(n_327), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g419 ( .A(n_331), .Y(n_419) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g348 ( .A(n_337), .B(n_338), .Y(n_348) );
INVx1_ASAP7_75t_L g401 ( .A(n_337), .Y(n_401) );
NOR3xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_375), .C(n_397), .Y(n_343) );
OAI211xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_349), .B(n_351), .C(n_356), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI21xp33_ASAP7_75t_L g351 ( .A1(n_346), .A2(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI211xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_359), .B(n_362), .C(n_369), .Y(n_356) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g380 ( .A(n_363), .Y(n_380) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_364), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_366), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g428 ( .A(n_366), .Y(n_428) );
AND2x2_ASAP7_75t_L g418 ( .A(n_368), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g388 ( .A(n_370), .Y(n_388) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx1_ASAP7_75t_L g396 ( .A(n_372), .Y(n_396) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_384), .A2(n_418), .B1(n_420), .B2(n_422), .C(n_427), .Y(n_417) );
OAI21xp33_ASAP7_75t_SL g432 ( .A1(n_389), .A2(n_433), .B(n_434), .Y(n_432) );
INVx2_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND4xp25_ASAP7_75t_L g397 ( .A(n_398), .B(n_408), .C(n_417), .D(n_431), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_402), .B1(n_405), .B2(n_406), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_426), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx3_ASAP7_75t_SL g748 ( .A(n_439), .Y(n_748) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_440), .Y(n_439) );
AND2x6_ASAP7_75t_SL g440 ( .A(n_441), .B(n_442), .Y(n_440) );
OR2x6_ASAP7_75t_SL g739 ( .A(n_441), .B(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g752 ( .A(n_441), .B(n_442), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_441), .B(n_740), .Y(n_763) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_442), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_447), .A2(n_739), .B1(n_746), .B2(n_747), .Y(n_745) );
OR2x6_ASAP7_75t_L g447 ( .A(n_448), .B(n_635), .Y(n_447) );
NAND3xp33_ASAP7_75t_SL g448 ( .A(n_449), .B(n_547), .C(n_602), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_488), .B1(n_511), .B2(n_515), .C(n_525), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_472), .Y(n_450) );
AND2x2_ASAP7_75t_SL g513 ( .A(n_451), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g546 ( .A(n_451), .Y(n_546) );
AND2x2_ASAP7_75t_L g591 ( .A(n_451), .B(n_528), .Y(n_591) );
AND2x4_ASAP7_75t_L g451 ( .A(n_452), .B(n_463), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g579 ( .A(n_453), .Y(n_579) );
INVx1_ASAP7_75t_L g589 ( .A(n_453), .Y(n_589) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_455), .B(n_461), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_454), .B(n_462), .Y(n_461) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_454), .A2(n_455), .B(n_461), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_460), .Y(n_455) );
OR2x2_ASAP7_75t_L g568 ( .A(n_463), .B(n_473), .Y(n_568) );
NAND2x1p5_ASAP7_75t_L g599 ( .A(n_463), .B(n_514), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_463), .B(n_480), .Y(n_612) );
INVx2_ASAP7_75t_L g621 ( .A(n_463), .Y(n_621) );
AND2x2_ASAP7_75t_L g642 ( .A(n_463), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g726 ( .A(n_463), .B(n_545), .Y(n_726) );
INVx4_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g554 ( .A(n_464), .B(n_480), .Y(n_554) );
AND2x2_ASAP7_75t_L g687 ( .A(n_464), .B(n_514), .Y(n_687) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_464), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_470), .Y(n_465) );
AND2x4_ASAP7_75t_L g641 ( .A(n_472), .B(n_642), .Y(n_641) );
AOI321xp33_ASAP7_75t_L g655 ( .A1(n_472), .A2(n_584), .A3(n_585), .B1(n_617), .B2(n_656), .C(n_659), .Y(n_655) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_480), .Y(n_472) );
BUFx3_ASAP7_75t_L g512 ( .A(n_473), .Y(n_512) );
INVx2_ASAP7_75t_L g545 ( .A(n_473), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_473), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g578 ( .A(n_473), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g611 ( .A(n_473), .Y(n_611) );
INVx5_ASAP7_75t_L g514 ( .A(n_480), .Y(n_514) );
NOR2x1_ASAP7_75t_SL g563 ( .A(n_480), .B(n_553), .Y(n_563) );
BUFx2_ASAP7_75t_L g658 ( .A(n_480), .Y(n_658) );
OR2x6_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVxp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_501), .Y(n_489) );
NOR2xp33_ASAP7_75t_SL g556 ( .A(n_490), .B(n_557), .Y(n_556) );
NOR4xp25_ASAP7_75t_L g659 ( .A(n_490), .B(n_653), .C(n_657), .D(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g697 ( .A(n_490), .Y(n_697) );
AND2x2_ASAP7_75t_L g731 ( .A(n_490), .B(n_671), .Y(n_731) );
BUFx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g532 ( .A(n_491), .Y(n_532) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g586 ( .A(n_492), .Y(n_586) );
OAI21x1_ASAP7_75t_SL g492 ( .A1(n_493), .A2(n_495), .B(n_499), .Y(n_492) );
INVx1_ASAP7_75t_L g500 ( .A(n_494), .Y(n_500) );
AOI33xp33_ASAP7_75t_L g727 ( .A1(n_501), .A2(n_529), .A3(n_560), .B1(n_576), .B2(n_682), .B3(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g517 ( .A(n_502), .B(n_518), .Y(n_517) );
AND2x4_ASAP7_75t_L g527 ( .A(n_502), .B(n_528), .Y(n_527) );
BUFx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g534 ( .A(n_503), .Y(n_534) );
INVxp67_ASAP7_75t_L g615 ( .A(n_503), .Y(n_615) );
AND2x2_ASAP7_75t_L g671 ( .A(n_503), .B(n_536), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_509), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_511), .A2(n_693), .B(n_694), .Y(n_692) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
AND2x2_ASAP7_75t_L g680 ( .A(n_512), .B(n_554), .Y(n_680) );
AND3x2_ASAP7_75t_L g682 ( .A(n_512), .B(n_566), .C(n_621), .Y(n_682) );
INVx3_ASAP7_75t_SL g634 ( .A(n_513), .Y(n_634) );
INVx4_ASAP7_75t_L g528 ( .A(n_514), .Y(n_528) );
AND2x2_ASAP7_75t_L g566 ( .A(n_514), .B(n_553), .Y(n_566) );
INVxp67_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g560 ( .A(n_518), .Y(n_560) );
AND2x4_ASAP7_75t_L g585 ( .A(n_518), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g648 ( .A(n_518), .B(n_536), .Y(n_648) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g618 ( .A(n_519), .Y(n_618) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_519), .Y(n_640) );
O2A1O1Ixp33_ASAP7_75t_R g525 ( .A1(n_526), .A2(n_529), .B(n_533), .C(n_544), .Y(n_525) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g577 ( .A(n_528), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_528), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_528), .B(n_545), .Y(n_706) );
INVx1_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g688 ( .A(n_530), .B(n_678), .Y(n_688) );
AND2x2_ASAP7_75t_SL g530 ( .A(n_531), .B(n_532), .Y(n_530) );
AND2x2_ASAP7_75t_L g535 ( .A(n_531), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g557 ( .A(n_531), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g573 ( .A(n_531), .B(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g606 ( .A(n_531), .B(n_586), .Y(n_606) );
AND2x4_ASAP7_75t_L g571 ( .A(n_532), .B(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g595 ( .A(n_532), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g633 ( .A(n_532), .B(n_558), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
AND2x2_ASAP7_75t_L g561 ( .A(n_534), .B(n_558), .Y(n_561) );
AND2x2_ASAP7_75t_L g576 ( .A(n_534), .B(n_536), .Y(n_576) );
BUFx2_ASAP7_75t_L g632 ( .A(n_534), .Y(n_632) );
AND2x2_ASAP7_75t_L g646 ( .A(n_534), .B(n_557), .Y(n_646) );
INVx2_ASAP7_75t_L g558 ( .A(n_536), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_538), .B(n_542), .Y(n_537) );
OAI22xp33_ASAP7_75t_L g594 ( .A1(n_544), .A2(n_595), .B1(n_597), .B2(n_601), .Y(n_594) );
INVx2_ASAP7_75t_SL g625 ( .A(n_544), .Y(n_625) );
OR2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
AND2x2_ASAP7_75t_L g600 ( .A(n_545), .B(n_553), .Y(n_600) );
INVx1_ASAP7_75t_L g707 ( .A(n_546), .Y(n_707) );
NOR3xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_580), .C(n_594), .Y(n_547) );
OAI221xp5_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_555), .B1(n_559), .B2(n_562), .C(n_564), .Y(n_548) );
INVx1_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .Y(n_550) );
INVxp67_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g608 ( .A(n_552), .Y(n_608) );
INVxp67_ASAP7_75t_SL g736 ( .A(n_552), .Y(n_736) );
INVx1_ASAP7_75t_L g699 ( .A(n_554), .Y(n_699) );
AND2x2_ASAP7_75t_SL g709 ( .A(n_554), .B(n_578), .Y(n_709) );
INVxp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_558), .B(n_586), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
OR2x2_ASAP7_75t_L g592 ( .A(n_560), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g670 ( .A(n_560), .Y(n_670) );
AND2x2_ASAP7_75t_L g605 ( .A(n_561), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g651 ( .A(n_563), .B(n_611), .Y(n_651) );
AND2x2_ASAP7_75t_L g728 ( .A(n_563), .B(n_726), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_569), .B1(n_576), .B2(n_577), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g587 ( .A(n_568), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
INVx2_ASAP7_75t_L g593 ( .A(n_571), .Y(n_593) );
AND2x4_ASAP7_75t_L g617 ( .A(n_571), .B(n_618), .Y(n_617) );
OAI21xp33_ASAP7_75t_SL g647 ( .A1(n_571), .A2(n_648), .B(n_649), .Y(n_647) );
AND2x2_ASAP7_75t_L g674 ( .A(n_571), .B(n_632), .Y(n_674) );
INVx2_ASAP7_75t_L g596 ( .A(n_572), .Y(n_596) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_572), .Y(n_629) );
INVx1_ASAP7_75t_SL g653 ( .A(n_573), .Y(n_653) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx2_ASAP7_75t_L g584 ( .A(n_575), .Y(n_584) );
AND2x4_ASAP7_75t_SL g678 ( .A(n_575), .B(n_596), .Y(n_678) );
AND2x2_ASAP7_75t_L g675 ( .A(n_578), .B(n_621), .Y(n_675) );
AND2x2_ASAP7_75t_L g701 ( .A(n_578), .B(n_687), .Y(n_701) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_579), .Y(n_623) );
INVx1_ASAP7_75t_L g643 ( .A(n_579), .Y(n_643) );
OAI22xp33_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_587), .B1(n_590), .B2(n_592), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_585), .B(n_596), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_585), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g724 ( .A(n_585), .Y(n_724) );
INVx2_ASAP7_75t_SL g649 ( .A(n_587), .Y(n_649) );
AND2x2_ASAP7_75t_L g661 ( .A(n_589), .B(n_621), .Y(n_661) );
INVx2_ASAP7_75t_L g667 ( .A(n_589), .Y(n_667) );
INVxp33_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g626 ( .A(n_592), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_595), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g717 ( .A(n_595), .Y(n_717) );
INVx1_ASAP7_75t_L g645 ( .A(n_597), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_598), .B(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g656 ( .A(n_600), .B(n_657), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_600), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_729) );
NOR3xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_624), .C(n_627), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_607), .B1(n_609), .B2(n_613), .C(n_616), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_SL g722 ( .A(n_607), .Y(n_722) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g691 ( .A(n_608), .B(n_657), .Y(n_691) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g622 ( .A(n_611), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g693 ( .A(n_613), .Y(n_693) );
OR2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g690 ( .A(n_614), .Y(n_690) );
INVx1_ASAP7_75t_L g696 ( .A(n_615), .Y(n_696) );
OR2x2_ASAP7_75t_L g719 ( .A(n_615), .B(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
INVx1_ASAP7_75t_SL g628 ( .A(n_618), .Y(n_628) );
AND2x2_ASAP7_75t_L g698 ( .A(n_618), .B(n_678), .Y(n_698) );
AND2x2_ASAP7_75t_SL g730 ( .A(n_618), .B(n_631), .Y(n_730) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
INVx1_ASAP7_75t_L g735 ( .A(n_621), .Y(n_735) );
INVx1_ASAP7_75t_L g685 ( .A(n_623), .Y(n_685) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
O2A1O1Ixp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B(n_630), .C(n_634), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_628), .B(n_678), .Y(n_702) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_631), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
AND2x2_ASAP7_75t_L g639 ( .A(n_633), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g720 ( .A(n_633), .Y(n_720) );
NAND4xp75_ASAP7_75t_L g635 ( .A(n_636), .B(n_692), .C(n_708), .D(n_729), .Y(n_635) );
NOR3x1_ASAP7_75t_L g636 ( .A(n_637), .B(n_654), .C(n_676), .Y(n_636) );
NAND4xp75_ASAP7_75t_L g637 ( .A(n_638), .B(n_644), .C(n_647), .D(n_650), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_639), .B(n_641), .Y(n_638) );
AND2x2_ASAP7_75t_L g689 ( .A(n_640), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g714 ( .A(n_641), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_SL g703 ( .A(n_646), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_662), .Y(n_654) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_658), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_668), .B(n_672), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI322xp33_ASAP7_75t_L g694 ( .A1(n_666), .A2(n_695), .A3(n_699), .B1(n_700), .B2(n_702), .C1(n_703), .C2(n_704), .Y(n_694) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_667), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_670), .B(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_671), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
OAI211xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_679), .B(n_681), .C(n_683), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_688), .B1(n_689), .B2(n_691), .Y(n_683) );
NOR2xp33_ASAP7_75t_SL g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx2_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B(n_698), .Y(n_695) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_701), .B(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_705), .B(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g711 ( .A(n_706), .B(n_712), .Y(n_711) );
O2A1O1Ixp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_710), .B(n_715), .C(n_718), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_711), .B(n_714), .Y(n_710) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OAI221xp5_ASAP7_75t_SL g718 ( .A1(n_719), .A2(n_721), .B1(n_723), .B2(n_725), .C(n_727), .Y(n_718) );
INVxp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
CKINVDCx11_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
CKINVDCx6p67_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_762), .Y(n_755) );
INVxp67_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g757 ( .A(n_758), .B(n_761), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_SL g783 ( .A(n_759), .B(n_761), .Y(n_783) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_759), .A2(n_788), .B(n_791), .Y(n_787) );
BUFx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
BUFx2_ASAP7_75t_L g773 ( .A(n_763), .Y(n_773) );
BUFx3_ASAP7_75t_L g778 ( .A(n_763), .Y(n_778) );
INVxp67_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AOI21xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_772), .B(n_774), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_768), .Y(n_771) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g791 ( .A(n_773), .Y(n_791) );
NOR2xp33_ASAP7_75t_SL g774 ( .A(n_775), .B(n_779), .Y(n_774) );
INVx1_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
BUFx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
CKINVDCx11_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
CKINVDCx8_ASAP7_75t_R g789 ( .A(n_790), .Y(n_789) );
endmodule