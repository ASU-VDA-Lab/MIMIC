module real_jpeg_16787_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_2),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_2),
.B(n_127),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_3),
.Y(n_125)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_4),
.Y(n_109)
);

AND2x4_ASAP7_75t_SL g16 ( 
.A(n_5),
.B(n_17),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_5),
.B(n_49),
.Y(n_48)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_5),
.B(n_57),
.Y(n_56)
);

AND2x4_ASAP7_75t_SL g68 ( 
.A(n_5),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_5),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_6),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_6),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_6),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_7),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_7),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_7),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_7),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_8),
.B(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_9),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_98),
.Y(n_11)
);

AOI21x1_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_64),
.B(n_97),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_53),
.Y(n_13)
);

NOR2xp67_ASAP7_75t_SL g97 ( 
.A(n_14),
.B(n_53),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_32),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_15),
.B(n_33),
.C(n_43),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_20),
.Y(n_15)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_16),
.Y(n_104)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_21),
.B(n_27),
.C(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_25),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_42),
.B2(n_43),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_39),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AO22x1_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_48),
.B(n_51),
.Y(n_121)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_56),
.C(n_60),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_55),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_60),
.B1(n_61),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_82),
.B(n_96),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_78),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_72),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_68),
.B1(n_72),
.B2(n_89),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2x1_ASAP7_75t_L g123 ( 
.A(n_68),
.B(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_90),
.B(n_95),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_88),
.Y(n_95)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_130),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_101),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_120),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.Y(n_105)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_110)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);


endmodule