module fake_netlist_5_2061_n_1812 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1812);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1812;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_783;
wire n_555;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1752;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_43),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_92),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_152),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_95),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_141),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_40),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_9),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_59),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_37),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_91),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_132),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_96),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_36),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_99),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_11),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_86),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_74),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_69),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_76),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_40),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_30),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_33),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_77),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_44),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_123),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_52),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_50),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_68),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_22),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_70),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_130),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_89),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_20),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_82),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_21),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_18),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_80),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_78),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_51),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_97),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_17),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_63),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_1),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_18),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_53),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_33),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_39),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_124),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_62),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_154),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_55),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_66),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_53),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_50),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_21),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_115),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_13),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_85),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_58),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_15),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_136),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_120),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_110),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_71),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_117),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_49),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_101),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_36),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_35),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_72),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_100),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_14),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_23),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_127),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_118),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_138),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_48),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_113),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_145),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_11),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_30),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_0),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_139),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_39),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_73),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_13),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_98),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_153),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_8),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_28),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_109),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_65),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_29),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_105),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_88),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_133),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_94),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_35),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_79),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_14),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_6),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_104),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_160),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_32),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_121),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_149),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_146),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_112),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_60),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_19),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_90),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_84),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_46),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_122),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_42),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_0),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_126),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_34),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_51),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_48),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_61),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_108),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_26),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_87),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_144),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_8),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_157),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_47),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_17),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_107),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_128),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_67),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_57),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_26),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_81),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_27),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_64),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_34),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_9),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_111),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_10),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_150),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_19),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_29),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_22),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_119),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_44),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_140),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_142),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_55),
.Y(n_316)
);

BUFx10_ASAP7_75t_L g317 ( 
.A(n_114),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_32),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_2),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_164),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g321 ( 
.A(n_255),
.B(n_1),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_172),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_284),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_173),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_208),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_R g326 ( 
.A(n_294),
.B(n_159),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_181),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_245),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_162),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_163),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_165),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g332 ( 
.A(n_255),
.B(n_2),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_174),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_284),
.Y(n_334)
);

NAND2xp33_ASAP7_75t_R g335 ( 
.A(n_171),
.B(n_3),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_277),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_287),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_284),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_293),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_284),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_176),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_189),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_208),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_189),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_178),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_192),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_280),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_309),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_192),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_179),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_171),
.B(n_3),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_280),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_168),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_264),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_264),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_307),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_307),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_290),
.B(n_4),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_290),
.B(n_4),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_193),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_187),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_191),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_182),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_258),
.B(n_5),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_182),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_198),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_258),
.B(n_5),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_309),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_202),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_274),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_186),
.Y(n_372)
);

INVxp33_ASAP7_75t_L g373 ( 
.A(n_186),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_205),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_199),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_274),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_201),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_213),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_214),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_240),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_199),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_215),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_196),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_161),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_169),
.B(n_6),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_291),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_212),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_169),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_222),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_224),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_212),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_238),
.B(n_7),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_225),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_227),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_188),
.B(n_7),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_323),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_321),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_371),
.B(n_232),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_323),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_334),
.B(n_180),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_390),
.Y(n_401)
);

CKINVDCx11_ASAP7_75t_R g402 ( 
.A(n_348),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_321),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_334),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_338),
.Y(n_405)
);

OA21x2_ASAP7_75t_L g406 ( 
.A1(n_388),
.A2(n_194),
.B(n_188),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_337),
.Y(n_407)
);

NAND2x1_ASAP7_75t_L g408 ( 
.A(n_337),
.B(n_287),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_337),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_337),
.Y(n_410)
);

AND2x6_ASAP7_75t_L g411 ( 
.A(n_337),
.B(n_287),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_338),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_337),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_339),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_365),
.B(n_228),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_339),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_341),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_341),
.B(n_180),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_358),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_358),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_388),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_364),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_376),
.B(n_232),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_364),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_343),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_376),
.B(n_194),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_376),
.B(n_195),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_343),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_366),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_345),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_366),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_368),
.B(n_230),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_372),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_375),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_375),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_385),
.B(n_233),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_345),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_381),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_332),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_395),
.B(n_236),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_381),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_387),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_377),
.B(n_195),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_387),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_391),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_380),
.B(n_237),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_347),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_335),
.A2(n_247),
.B1(n_319),
.B2(n_204),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_347),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_391),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_350),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_350),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_355),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_377),
.B(n_203),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_355),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_356),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_356),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_357),
.B(n_241),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_357),
.B(n_352),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_392),
.B(n_185),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_377),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_392),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_359),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_329),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_332),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_463),
.B(n_330),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_401),
.Y(n_469)
);

AND2x6_ASAP7_75t_L g470 ( 
.A(n_465),
.B(n_185),
.Y(n_470)
);

BUFx4f_ASAP7_75t_L g471 ( 
.A(n_406),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_406),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_450),
.A2(n_360),
.B1(n_361),
.B2(n_325),
.Y(n_473)
);

OR2x6_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_203),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_466),
.B(n_331),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_333),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_401),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_407),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_422),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_466),
.B(n_342),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_373),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_R g482 ( 
.A(n_398),
.B(n_346),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_406),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_417),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_407),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_417),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_406),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_407),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_417),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_463),
.B(n_351),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_L g492 ( 
.A(n_438),
.B(n_326),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_396),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_396),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_463),
.B(n_362),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_407),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_399),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_399),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_397),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_402),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_404),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_404),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_463),
.B(n_207),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_405),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_416),
.B(n_383),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_405),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_412),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_412),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_424),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_407),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_465),
.B(n_363),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_422),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_407),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_414),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_438),
.B(n_367),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_450),
.A2(n_344),
.B1(n_369),
.B2(n_353),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_465),
.B(n_370),
.Y(n_517)
);

AND3x2_ASAP7_75t_L g518 ( 
.A(n_397),
.B(n_349),
.C(n_262),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_414),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_418),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_427),
.B(n_207),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_424),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_407),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_418),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_416),
.B(n_383),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_442),
.B(n_374),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_462),
.A2(n_266),
.B1(n_238),
.B2(n_243),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_422),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_426),
.Y(n_529)
);

AO22x1_ASAP7_75t_L g530 ( 
.A1(n_462),
.A2(n_250),
.B1(n_266),
.B2(n_259),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_400),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_403),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_403),
.B(n_386),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_467),
.B(n_386),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_422),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_462),
.A2(n_259),
.B1(n_311),
.B2(n_305),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_422),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_441),
.B(n_378),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_427),
.B(n_379),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_415),
.B(n_382),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_442),
.B(n_389),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_415),
.B(n_393),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_409),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_448),
.B(n_394),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_448),
.B(n_354),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_426),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_434),
.B(n_257),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_400),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_427),
.B(n_217),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_422),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_409),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_400),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_441),
.B(n_467),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_400),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_409),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_398),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_428),
.B(n_217),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_426),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_426),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_426),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_462),
.A2(n_243),
.B1(n_318),
.B2(n_289),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_434),
.B(n_340),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_400),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_422),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_419),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_426),
.Y(n_566)
);

AO22x2_ASAP7_75t_L g567 ( 
.A1(n_462),
.A2(n_292),
.B1(n_289),
.B2(n_305),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_445),
.B(n_273),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_424),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_398),
.B(n_201),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_419),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_419),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_409),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_445),
.B(n_242),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_426),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_409),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_419),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_429),
.Y(n_578)
);

BUFx6f_ASAP7_75t_SL g579 ( 
.A(n_464),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_419),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_429),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_429),
.Y(n_582)
);

INVx6_ASAP7_75t_L g583 ( 
.A(n_428),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_423),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_464),
.B(n_201),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_428),
.B(n_445),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_456),
.A2(n_235),
.B1(n_197),
.B2(n_316),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_429),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_456),
.B(n_249),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_429),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_456),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_429),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_423),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_425),
.Y(n_594)
);

INVxp33_ASAP7_75t_L g595 ( 
.A(n_402),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_425),
.Y(n_596)
);

BUFx10_ASAP7_75t_L g597 ( 
.A(n_430),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_429),
.Y(n_598)
);

AND2x6_ASAP7_75t_L g599 ( 
.A(n_461),
.B(n_218),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_439),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_430),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_439),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_409),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_461),
.A2(n_318),
.B1(n_292),
.B2(n_248),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_408),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_432),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_460),
.B(n_320),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_409),
.Y(n_608)
);

INVx5_ASAP7_75t_L g609 ( 
.A(n_411),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_432),
.B(n_229),
.Y(n_610)
);

BUFx6f_ASAP7_75t_SL g611 ( 
.A(n_433),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_439),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_460),
.B(n_433),
.Y(n_613)
);

INVx5_ASAP7_75t_L g614 ( 
.A(n_411),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_435),
.B(n_253),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_435),
.B(n_263),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_436),
.B(n_229),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_408),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_471),
.B(n_287),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_509),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_509),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_556),
.B(n_322),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_515),
.B(n_431),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_493),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_493),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_599),
.A2(n_250),
.B1(n_248),
.B2(n_311),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_482),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_509),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_522),
.B(n_436),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_501),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_526),
.B(n_431),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_501),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_599),
.A2(n_486),
.B1(n_567),
.B2(n_472),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_499),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_556),
.B(n_324),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_504),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_541),
.B(n_431),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_569),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_511),
.B(n_166),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_522),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_547),
.B(n_431),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_471),
.A2(n_410),
.B(n_408),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_517),
.B(n_167),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_499),
.B(n_170),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_597),
.B(n_327),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_471),
.B(n_540),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_534),
.B(n_542),
.Y(n_647)
);

NOR3xp33_ASAP7_75t_L g648 ( 
.A(n_505),
.B(n_256),
.C(n_184),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_591),
.B(n_431),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_522),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_591),
.B(n_449),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_583),
.Y(n_652)
);

O2A1O1Ixp5_ASAP7_75t_L g653 ( 
.A1(n_472),
.A2(n_218),
.B(n_262),
.C(n_260),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_534),
.B(n_175),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_613),
.B(n_449),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_597),
.B(n_328),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_597),
.B(n_336),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_481),
.B(n_437),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_504),
.Y(n_659)
);

OR2x2_ASAP7_75t_SL g660 ( 
.A(n_544),
.B(n_562),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_586),
.B(n_449),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_583),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_492),
.A2(n_299),
.B1(n_265),
.B2(n_268),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_583),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_506),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_586),
.B(n_449),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_553),
.B(n_177),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_481),
.B(n_449),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_583),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_521),
.B(n_437),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_475),
.B(n_439),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_480),
.B(n_439),
.Y(n_672)
);

NOR2xp67_ASAP7_75t_L g673 ( 
.A(n_545),
.B(n_440),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_597),
.B(n_269),
.Y(n_674)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_525),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_584),
.B(n_439),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_584),
.B(n_439),
.Y(n_677)
);

NOR3xp33_ASAP7_75t_L g678 ( 
.A(n_533),
.B(n_246),
.C(n_239),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_607),
.B(n_183),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_539),
.B(n_532),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_521),
.B(n_440),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_593),
.B(n_231),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_506),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_507),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_593),
.B(n_231),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_516),
.B(n_443),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_507),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_594),
.B(n_244),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_594),
.B(n_244),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_520),
.Y(n_690)
);

INVx8_ASAP7_75t_L g691 ( 
.A(n_579),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_596),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_596),
.B(n_251),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_601),
.B(n_251),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_486),
.B(n_287),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_601),
.B(n_254),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_539),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_532),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_606),
.B(n_254),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_486),
.B(n_271),
.Y(n_700)
);

AO221x1_ASAP7_75t_L g701 ( 
.A1(n_567),
.A2(n_260),
.B1(n_261),
.B2(n_272),
.C(n_298),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_520),
.Y(n_702)
);

AND2x2_ASAP7_75t_SL g703 ( 
.A(n_468),
.B(n_476),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_606),
.B(n_261),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_491),
.B(n_272),
.Y(n_705)
);

BUFx8_ASAP7_75t_L g706 ( 
.A(n_579),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_532),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_570),
.B(n_190),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_494),
.Y(n_709)
);

OR2x6_ASAP7_75t_L g710 ( 
.A(n_530),
.B(n_298),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_531),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_531),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_548),
.Y(n_713)
);

INVx5_ASAP7_75t_L g714 ( 
.A(n_470),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_538),
.B(n_200),
.Y(n_715)
);

NOR2xp67_ASAP7_75t_L g716 ( 
.A(n_495),
.B(n_443),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_494),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_532),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_548),
.B(n_275),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_497),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_SL g721 ( 
.A(n_579),
.B(n_201),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_568),
.B(n_283),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_516),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_605),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_518),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_585),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_477),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_497),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_549),
.B(n_301),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_587),
.B(n_288),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_549),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_587),
.B(n_296),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_574),
.B(n_303),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_552),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_483),
.B(n_301),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_605),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_473),
.B(n_444),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_498),
.Y(n_738)
);

NAND2xp33_ASAP7_75t_L g739 ( 
.A(n_599),
.B(n_306),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_473),
.B(n_206),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_552),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_483),
.B(n_308),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_521),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_521),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_488),
.B(n_308),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_488),
.B(n_315),
.Y(n_746)
);

INVxp33_ASAP7_75t_L g747 ( 
.A(n_610),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_554),
.Y(n_748)
);

NOR3xp33_ASAP7_75t_L g749 ( 
.A(n_469),
.B(n_220),
.C(n_209),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_554),
.B(n_315),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_L g751 ( 
.A(n_589),
.B(n_444),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_563),
.B(n_446),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_563),
.B(n_446),
.Y(n_753)
);

NOR2x1p5_ASAP7_75t_L g754 ( 
.A(n_615),
.B(n_210),
.Y(n_754)
);

BUFx5_ASAP7_75t_L g755 ( 
.A(n_605),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_616),
.B(n_211),
.Y(n_756)
);

AND2x6_ASAP7_75t_SL g757 ( 
.A(n_474),
.B(n_223),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_474),
.A2(n_312),
.B1(n_314),
.B2(n_452),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_474),
.B(n_216),
.Y(n_759)
);

NOR2xp67_ASAP7_75t_L g760 ( 
.A(n_565),
.B(n_447),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_565),
.B(n_413),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_571),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_571),
.B(n_447),
.Y(n_763)
);

INVxp67_ASAP7_75t_SL g764 ( 
.A(n_478),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_SL g765 ( 
.A(n_579),
.B(n_611),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_557),
.B(n_452),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_572),
.B(n_410),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_572),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_474),
.B(n_219),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_557),
.B(n_278),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_474),
.B(n_221),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_618),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_498),
.B(n_226),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_577),
.B(n_410),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_577),
.B(n_410),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_502),
.B(n_234),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_502),
.B(n_252),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_557),
.B(n_278),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_557),
.B(n_453),
.Y(n_779)
);

OAI221xp5_ASAP7_75t_L g780 ( 
.A1(n_604),
.A2(n_536),
.B1(n_527),
.B2(n_561),
.C(n_617),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_580),
.B(n_451),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_SL g782 ( 
.A(n_611),
.B(n_500),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_508),
.B(n_267),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_580),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_610),
.B(n_617),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_508),
.B(n_270),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_514),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_503),
.B(n_413),
.Y(n_788)
);

NOR2xp67_ASAP7_75t_L g789 ( 
.A(n_514),
.B(n_453),
.Y(n_789)
);

INVxp67_ASAP7_75t_SL g790 ( 
.A(n_478),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_530),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_785),
.B(n_599),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_644),
.Y(n_793)
);

NOR2x1_ASAP7_75t_L g794 ( 
.A(n_647),
.B(n_618),
.Y(n_794)
);

OAI321xp33_ASAP7_75t_L g795 ( 
.A1(n_740),
.A2(n_519),
.A3(n_524),
.B1(n_455),
.B2(n_459),
.C(n_454),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_724),
.A2(n_611),
.B1(n_618),
.B2(n_503),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_731),
.B(n_599),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_L g798 ( 
.A1(n_695),
.A2(n_503),
.B(n_599),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_658),
.B(n_599),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_671),
.A2(n_550),
.B(n_479),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_713),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_672),
.A2(n_550),
.B(n_479),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_642),
.A2(n_619),
.B(n_668),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_647),
.A2(n_679),
.B1(n_697),
.B2(n_743),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_713),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_619),
.A2(n_550),
.B(n_479),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_772),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_623),
.A2(n_550),
.B(n_479),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_755),
.B(n_609),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_673),
.B(n_519),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_631),
.A2(n_528),
.B(n_564),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_709),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_637),
.A2(n_528),
.B(n_564),
.Y(n_813)
);

BUFx12f_ASAP7_75t_L g814 ( 
.A(n_727),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_695),
.A2(n_503),
.B(n_524),
.Y(n_815)
);

AOI21xp33_ASAP7_75t_L g816 ( 
.A1(n_679),
.A2(n_567),
.B(n_595),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_772),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_724),
.A2(n_611),
.B1(n_567),
.B2(n_537),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_646),
.A2(n_528),
.B(n_564),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_SL g820 ( 
.A(n_765),
.B(n_691),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_634),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_755),
.B(n_609),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_736),
.A2(n_512),
.B1(n_537),
.B2(n_535),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_646),
.A2(n_528),
.B(n_564),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_639),
.B(n_470),
.Y(n_825)
);

AOI21xp33_ASAP7_75t_L g826 ( 
.A1(n_740),
.A2(n_313),
.B(n_281),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_736),
.A2(n_512),
.B1(n_535),
.B2(n_537),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_780),
.A2(n_459),
.B(n_454),
.C(n_455),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_709),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_639),
.B(n_643),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_627),
.B(n_478),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_661),
.A2(n_513),
.B(n_551),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_666),
.A2(n_513),
.B(n_551),
.Y(n_833)
);

AOI221xp5_ASAP7_75t_L g834 ( 
.A1(n_723),
.A2(n_715),
.B1(n_644),
.B2(n_708),
.C(n_654),
.Y(n_834)
);

AO21x1_ASAP7_75t_L g835 ( 
.A1(n_700),
.A2(n_512),
.B(n_535),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_691),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_641),
.A2(n_655),
.B(n_664),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_664),
.A2(n_551),
.B(n_513),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_643),
.B(n_470),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_638),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_788),
.A2(n_551),
.B(n_513),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_629),
.B(n_470),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_747),
.B(n_223),
.Y(n_843)
);

NAND3xp33_ASAP7_75t_L g844 ( 
.A(n_654),
.B(n_302),
.C(n_304),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_717),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_737),
.A2(n_300),
.B(n_310),
.C(n_295),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_686),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_SL g848 ( 
.A(n_691),
.B(n_278),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_788),
.A2(n_513),
.B(n_551),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_755),
.B(n_609),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_717),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_629),
.B(n_470),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_660),
.B(n_478),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_711),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_755),
.B(n_609),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_756),
.B(n_692),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_756),
.B(n_470),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_649),
.A2(n_513),
.B(n_551),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_751),
.B(n_670),
.Y(n_859)
);

INVx4_ASAP7_75t_L g860 ( 
.A(n_772),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_670),
.B(n_470),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_633),
.A2(n_559),
.B1(n_612),
.B2(n_529),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_681),
.B(n_485),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_675),
.B(n_223),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_720),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_651),
.A2(n_576),
.B(n_614),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_720),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_772),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_764),
.A2(n_576),
.B(n_614),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_681),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_766),
.B(n_728),
.Y(n_871)
);

AO21x1_ASAP7_75t_L g872 ( 
.A1(n_700),
.A2(n_612),
.B(n_582),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_790),
.A2(n_576),
.B(n_614),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_755),
.B(n_609),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_766),
.B(n_529),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_728),
.B(n_485),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_738),
.B(n_485),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_653),
.A2(n_742),
.B(n_735),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_620),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_698),
.B(n_223),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_738),
.B(n_485),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_791),
.B(n_489),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_779),
.Y(n_883)
);

OAI21xp33_ASAP7_75t_L g884 ( 
.A1(n_715),
.A2(n_285),
.B(n_279),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_767),
.A2(n_576),
.B(n_614),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_787),
.B(n_489),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_787),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_716),
.B(n_489),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_774),
.A2(n_576),
.B(n_614),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_775),
.A2(n_576),
.B(n_614),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_755),
.B(n_609),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_624),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_781),
.A2(n_546),
.B(n_558),
.Y(n_893)
);

NAND3xp33_ASAP7_75t_L g894 ( 
.A(n_667),
.B(n_276),
.C(n_282),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_779),
.B(n_489),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_712),
.B(n_496),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_701),
.A2(n_278),
.B1(n_297),
.B2(n_317),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_708),
.A2(n_286),
.B(n_420),
.C(n_421),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_621),
.Y(n_899)
);

NOR2x1_ASAP7_75t_R g900 ( 
.A(n_622),
.B(n_297),
.Y(n_900)
);

BUFx12f_ASAP7_75t_L g901 ( 
.A(n_706),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_734),
.B(n_496),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_744),
.A2(n_546),
.B1(n_558),
.B2(n_602),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_741),
.B(n_748),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_762),
.B(n_768),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_745),
.A2(n_559),
.B(n_560),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_784),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_628),
.B(n_496),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_746),
.A2(n_761),
.B(n_703),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_640),
.B(n_496),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_650),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_624),
.Y(n_912)
);

BUFx8_ASAP7_75t_L g913 ( 
.A(n_725),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_703),
.B(n_510),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_705),
.B(n_510),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_761),
.A2(n_560),
.B(n_566),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_625),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_635),
.B(n_510),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_759),
.A2(n_420),
.B(n_421),
.C(n_458),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_759),
.A2(n_769),
.B(n_771),
.C(n_729),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_625),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_760),
.A2(n_566),
.B(n_575),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_710),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_680),
.B(n_510),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_633),
.A2(n_588),
.B1(n_575),
.B2(n_602),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_SL g926 ( 
.A1(n_730),
.A2(n_592),
.B(n_598),
.C(n_600),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_752),
.A2(n_763),
.B(n_753),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_652),
.A2(n_588),
.B(n_578),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_773),
.B(n_608),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_630),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_773),
.B(n_608),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_662),
.A2(n_578),
.B(n_581),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_714),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_669),
.B(n_581),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_726),
.A2(n_582),
.B1(n_590),
.B2(n_600),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_707),
.B(n_297),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_632),
.A2(n_590),
.B(n_592),
.Y(n_937)
);

AOI211xp5_ASAP7_75t_L g938 ( 
.A1(n_667),
.A2(n_732),
.B(n_648),
.C(n_678),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_776),
.B(n_608),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_632),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_776),
.B(n_608),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_777),
.B(n_783),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_719),
.A2(n_676),
.B(n_677),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_636),
.Y(n_944)
);

O2A1O1Ixp5_ASAP7_75t_L g945 ( 
.A1(n_719),
.A2(n_600),
.B(n_598),
.C(n_592),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_777),
.B(n_603),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_636),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_659),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_718),
.B(n_297),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_783),
.B(n_603),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_786),
.B(n_317),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_659),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_710),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_665),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_665),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_750),
.A2(n_598),
.B(n_603),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_786),
.B(n_603),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_789),
.B(n_683),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_683),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_684),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_714),
.A2(n_573),
.B(n_555),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_684),
.A2(n_573),
.B(n_555),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_687),
.A2(n_573),
.B(n_555),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_714),
.B(n_573),
.Y(n_964)
);

AO21x1_ASAP7_75t_L g965 ( 
.A1(n_769),
.A2(n_484),
.B(n_487),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_687),
.B(n_555),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_682),
.A2(n_484),
.B(n_487),
.C(n_490),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_690),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_690),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_754),
.B(n_749),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_702),
.B(n_543),
.Y(n_971)
);

AOI21x1_ASAP7_75t_L g972 ( 
.A1(n_733),
.A2(n_702),
.B(n_688),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_685),
.Y(n_973)
);

INVx11_ASAP7_75t_L g974 ( 
.A(n_706),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_689),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_771),
.A2(n_543),
.B1(n_523),
.B2(n_490),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_693),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_714),
.B(n_543),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_739),
.A2(n_523),
.B(n_543),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_645),
.B(n_317),
.Y(n_980)
);

NOR2xp67_ASAP7_75t_L g981 ( 
.A(n_663),
.B(n_523),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_694),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_696),
.Y(n_983)
);

NOR2xp67_ASAP7_75t_L g984 ( 
.A(n_814),
.B(n_656),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_803),
.A2(n_778),
.B(n_770),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_836),
.B(n_657),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_821),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_812),
.Y(n_988)
);

AOI21xp33_ASAP7_75t_L g989 ( 
.A1(n_830),
.A2(n_721),
.B(n_626),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_812),
.Y(n_990)
);

OAI22x1_ASAP7_75t_L g991 ( 
.A1(n_793),
.A2(n_847),
.B1(n_804),
.B2(n_923),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_942),
.A2(n_722),
.B(n_674),
.C(n_699),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_837),
.A2(n_626),
.B(n_413),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_817),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_834),
.A2(n_710),
.B1(n_704),
.B2(n_758),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_829),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_829),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_856),
.B(n_782),
.Y(n_998)
);

OAI21xp33_ASAP7_75t_L g999 ( 
.A1(n_826),
.A2(n_757),
.B(n_458),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_927),
.A2(n_413),
.B(n_523),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_983),
.B(n_458),
.Y(n_1001)
);

OAI21xp33_ASAP7_75t_SL g1002 ( 
.A1(n_815),
.A2(n_798),
.B(n_973),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_SL g1003 ( 
.A1(n_853),
.A2(n_457),
.B(n_451),
.C(n_317),
.Y(n_1003)
);

AOI21x1_ASAP7_75t_L g1004 ( 
.A1(n_914),
.A2(n_457),
.B(n_451),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_843),
.B(n_457),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_865),
.Y(n_1006)
);

NAND2xp33_ASAP7_75t_L g1007 ( 
.A(n_920),
.B(n_411),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_800),
.A2(n_802),
.B(n_878),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_920),
.A2(n_457),
.B(n_451),
.C(n_413),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_R g1010 ( 
.A(n_820),
.B(n_158),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_951),
.A2(n_411),
.B1(n_413),
.B2(n_148),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_865),
.Y(n_1012)
);

BUFx2_ASAP7_75t_SL g1013 ( 
.A(n_836),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_864),
.B(n_10),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_867),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_977),
.B(n_411),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_853),
.A2(n_938),
.B1(n_859),
.B2(n_918),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_913),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_982),
.B(n_411),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_867),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_840),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_SL g1022 ( 
.A1(n_898),
.A2(n_147),
.B(n_143),
.C(n_137),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_904),
.A2(n_413),
.B1(n_15),
.B2(n_16),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_817),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_905),
.A2(n_12),
.B1(n_16),
.B2(n_20),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_817),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_868),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_840),
.B(n_816),
.Y(n_1028)
);

NOR2x1_ASAP7_75t_SL g1029 ( 
.A(n_868),
.B(n_103),
.Y(n_1029)
);

CKINVDCx11_ASAP7_75t_R g1030 ( 
.A(n_901),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_975),
.B(n_411),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_806),
.A2(n_411),
.B(n_135),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_808),
.A2(n_411),
.B(n_134),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_884),
.B(n_12),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_887),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_SL g1036 ( 
.A1(n_898),
.A2(n_131),
.B(n_129),
.C(n_102),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_868),
.Y(n_1037)
);

INVx4_ASAP7_75t_L g1038 ( 
.A(n_868),
.Y(n_1038)
);

CKINVDCx16_ASAP7_75t_R g1039 ( 
.A(n_848),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_882),
.B(n_411),
.Y(n_1040)
);

OAI21xp33_ASAP7_75t_L g1041 ( 
.A1(n_980),
.A2(n_23),
.B(n_24),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_811),
.A2(n_93),
.B(n_83),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_882),
.B(n_75),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_R g1044 ( 
.A(n_807),
.B(n_56),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_923),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_909),
.A2(n_24),
.B(n_25),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_R g1047 ( 
.A(n_807),
.B(n_25),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_813),
.A2(n_56),
.B(n_28),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_953),
.B(n_27),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_857),
.A2(n_31),
.B(n_37),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_918),
.A2(n_31),
.B(n_38),
.C(n_41),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_953),
.B(n_38),
.Y(n_1052)
);

BUFx12f_ASAP7_75t_L g1053 ( 
.A(n_913),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_854),
.B(n_41),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_907),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_794),
.B(n_45),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_879),
.B(n_46),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_870),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_879),
.B(n_47),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_871),
.A2(n_846),
.B1(n_828),
.B2(n_883),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_825),
.A2(n_49),
.B(n_52),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_899),
.B(n_54),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_899),
.B(n_54),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_839),
.A2(n_838),
.B(n_891),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_801),
.B(n_805),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_809),
.A2(n_891),
.B(n_855),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_809),
.A2(n_850),
.B(n_855),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_822),
.A2(n_850),
.B(n_874),
.Y(n_1068)
);

INVx4_ASAP7_75t_L g1069 ( 
.A(n_870),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_870),
.B(n_844),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_846),
.A2(n_810),
.B(n_828),
.C(n_919),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_970),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_SL g1073 ( 
.A1(n_924),
.A2(n_831),
.B(n_795),
.C(n_897),
.Y(n_1073)
);

O2A1O1Ixp5_ASAP7_75t_L g1074 ( 
.A1(n_965),
.A2(n_872),
.B(n_835),
.C(n_919),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_970),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_894),
.B(n_936),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_845),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_822),
.A2(n_874),
.B(n_824),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_831),
.B(n_911),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_880),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_949),
.B(n_900),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_851),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_875),
.B(n_892),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_912),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_875),
.B(n_860),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_892),
.B(n_921),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_819),
.A2(n_929),
.B(n_931),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_799),
.A2(n_818),
.B1(n_792),
.B2(n_939),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_924),
.A2(n_943),
.B(n_797),
.C(n_950),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_863),
.B(n_895),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_941),
.B(n_946),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_957),
.A2(n_833),
.B(n_832),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_921),
.B(n_940),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_860),
.B(n_796),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_932),
.A2(n_915),
.B(n_963),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_935),
.A2(n_926),
.B(n_925),
.C(n_862),
.Y(n_1096)
);

O2A1O1Ixp5_ASAP7_75t_L g1097 ( 
.A1(n_945),
.A2(n_972),
.B(n_979),
.C(n_906),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_933),
.Y(n_1098)
);

BUFx12f_ASAP7_75t_L g1099 ( 
.A(n_974),
.Y(n_1099)
);

BUFx12f_ASAP7_75t_L g1100 ( 
.A(n_933),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_933),
.Y(n_1101)
);

INVxp67_ASAP7_75t_SL g1102 ( 
.A(n_955),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_926),
.A2(n_958),
.B(n_861),
.C(n_842),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_917),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_852),
.A2(n_897),
.B1(n_940),
.B2(n_948),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_962),
.A2(n_858),
.B(n_873),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_981),
.A2(n_976),
.B(n_893),
.C(n_967),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_869),
.A2(n_841),
.B(n_849),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_948),
.B(n_952),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_896),
.A2(n_902),
.B(n_947),
.C(n_968),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_866),
.A2(n_888),
.B(n_964),
.Y(n_1111)
);

INVx4_ASAP7_75t_L g1112 ( 
.A(n_952),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_934),
.A2(n_930),
.B1(n_944),
.B2(n_960),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_954),
.A2(n_969),
.B1(n_959),
.B2(n_903),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_954),
.B(n_959),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_934),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_969),
.A2(n_910),
.B1(n_908),
.B2(n_876),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_877),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_881),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_964),
.A2(n_978),
.B(n_886),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_966),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_971),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_978),
.B(n_823),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_937),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_827),
.B(n_956),
.Y(n_1125)
);

O2A1O1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_916),
.A2(n_928),
.B(n_922),
.C(n_890),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_885),
.A2(n_889),
.B(n_961),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_803),
.A2(n_471),
.B(n_837),
.Y(n_1128)
);

INVx3_ASAP7_75t_SL g1129 ( 
.A(n_970),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_R g1130 ( 
.A(n_814),
.B(n_727),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_834),
.B(n_942),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_803),
.A2(n_471),
.B(n_837),
.Y(n_1132)
);

INVx5_ASAP7_75t_L g1133 ( 
.A(n_933),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1131),
.A2(n_998),
.B(n_989),
.C(n_995),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1087),
.A2(n_1008),
.B(n_1128),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1132),
.A2(n_1091),
.B(n_1106),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1092),
.A2(n_1095),
.B(n_1089),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1021),
.B(n_987),
.Y(n_1138)
);

INVx6_ASAP7_75t_SL g1139 ( 
.A(n_986),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1078),
.A2(n_1108),
.B(n_1127),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_1080),
.B(n_1028),
.Y(n_1141)
);

AO31x2_ASAP7_75t_L g1142 ( 
.A1(n_1009),
.A2(n_1107),
.A3(n_1088),
.B(n_1125),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_SL g1143 ( 
.A1(n_1073),
.A2(n_989),
.B(n_992),
.C(n_1046),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1127),
.A2(n_1111),
.B(n_1064),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1017),
.B(n_1090),
.Y(n_1145)
);

BUFx12f_ASAP7_75t_L g1146 ( 
.A(n_1030),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_995),
.A2(n_1046),
.B(n_1034),
.C(n_1051),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_988),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1014),
.B(n_1072),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_985),
.A2(n_1002),
.B(n_993),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1081),
.A2(n_1076),
.B1(n_999),
.B2(n_1075),
.Y(n_1151)
);

NOR2xp67_ASAP7_75t_L g1152 ( 
.A(n_991),
.B(n_1099),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1097),
.A2(n_1126),
.B(n_1066),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1096),
.A2(n_1088),
.B(n_1094),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_1060),
.A2(n_1105),
.A3(n_1114),
.B(n_1124),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1041),
.A2(n_1023),
.B(n_1025),
.C(n_1062),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_1045),
.B(n_1129),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1060),
.A2(n_1105),
.A3(n_1114),
.B(n_1117),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_SL g1159 ( 
.A1(n_1029),
.A2(n_1071),
.B(n_1079),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1116),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1084),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1039),
.B(n_1057),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1104),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1067),
.A2(n_1068),
.B(n_1000),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1023),
.A2(n_1025),
.B(n_1063),
.C(n_1054),
.Y(n_1165)
);

AOI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1004),
.A2(n_1043),
.B(n_1070),
.Y(n_1166)
);

OAI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_984),
.A2(n_1056),
.B1(n_1043),
.B2(n_1059),
.Y(n_1167)
);

OR2x6_ASAP7_75t_L g1168 ( 
.A(n_1013),
.B(n_1100),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1005),
.B(n_1118),
.Y(n_1169)
);

NOR2xp67_ASAP7_75t_L g1170 ( 
.A(n_986),
.B(n_1069),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1121),
.B(n_1122),
.Y(n_1171)
);

AO21x2_ASAP7_75t_L g1172 ( 
.A1(n_1003),
.A2(n_1007),
.B(n_1033),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1103),
.A2(n_1110),
.B(n_1117),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1120),
.A2(n_1042),
.B(n_1123),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1074),
.A2(n_1048),
.B(n_1061),
.Y(n_1175)
);

AO31x2_ASAP7_75t_L g1176 ( 
.A1(n_1050),
.A2(n_1032),
.A3(n_1112),
.B(n_1040),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1065),
.B(n_1049),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1052),
.B(n_1001),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1011),
.A2(n_1113),
.B(n_1109),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_1133),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_SL g1181 ( 
.A1(n_1053),
.A2(n_1018),
.B1(n_1055),
.B2(n_1069),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1119),
.B(n_1077),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_1024),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1109),
.A2(n_1086),
.B(n_1093),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1082),
.B(n_1044),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_L g1186 ( 
.A(n_1055),
.B(n_1022),
.C(n_1036),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1058),
.B(n_1010),
.Y(n_1187)
);

NAND2xp33_ASAP7_75t_SL g1188 ( 
.A(n_1130),
.B(n_1058),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1115),
.A2(n_1006),
.B(n_1035),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1083),
.B(n_990),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1016),
.A2(n_1019),
.B(n_1015),
.C(n_1012),
.Y(n_1191)
);

BUFx12f_ASAP7_75t_L g1192 ( 
.A(n_1024),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1047),
.B(n_996),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_997),
.A2(n_1031),
.B(n_1020),
.C(n_1085),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1112),
.A2(n_994),
.A3(n_1038),
.B(n_1102),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1133),
.A2(n_994),
.B(n_1038),
.Y(n_1196)
);

OA21x2_ASAP7_75t_L g1197 ( 
.A1(n_1027),
.A2(n_1026),
.B(n_1037),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1026),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1026),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1133),
.A2(n_1101),
.B(n_1037),
.Y(n_1200)
);

CKINVDCx16_ASAP7_75t_R g1201 ( 
.A(n_1037),
.Y(n_1201)
);

O2A1O1Ixp5_ASAP7_75t_L g1202 ( 
.A1(n_1098),
.A2(n_830),
.B(n_942),
.C(n_1131),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_SL g1203 ( 
.A(n_1018),
.Y(n_1203)
);

O2A1O1Ixp33_ASAP7_75t_SL g1204 ( 
.A1(n_1131),
.A2(n_830),
.B(n_942),
.C(n_920),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1131),
.A2(n_942),
.B1(n_830),
.B2(n_834),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1131),
.A2(n_834),
.B(n_830),
.C(n_942),
.Y(n_1206)
);

NOR4xp25_ASAP7_75t_L g1207 ( 
.A(n_1131),
.B(n_942),
.C(n_830),
.D(n_1051),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_987),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1078),
.A2(n_1108),
.B(n_1127),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1078),
.A2(n_1108),
.B(n_1127),
.Y(n_1210)
);

NAND3xp33_ASAP7_75t_SL g1211 ( 
.A(n_1131),
.B(n_834),
.C(n_830),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1084),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_987),
.Y(n_1213)
);

NOR2x1_ASAP7_75t_R g1214 ( 
.A(n_1099),
.B(n_727),
.Y(n_1214)
);

CKINVDCx11_ASAP7_75t_R g1215 ( 
.A(n_1030),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_987),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1078),
.A2(n_1108),
.B(n_1127),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1131),
.B(n_793),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1100),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_SL g1220 ( 
.A1(n_1131),
.A2(n_834),
.B(n_740),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1080),
.B(n_847),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1131),
.A2(n_830),
.B(n_942),
.C(n_834),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1131),
.A2(n_834),
.B(n_830),
.C(n_942),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1080),
.B(n_834),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1084),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1131),
.B(n_830),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1087),
.A2(n_830),
.B(n_1008),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1080),
.B(n_847),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1100),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1084),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1087),
.A2(n_830),
.B(n_1008),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1131),
.A2(n_830),
.B(n_1009),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_SL g1233 ( 
.A1(n_1039),
.A2(n_660),
.B1(n_723),
.B2(n_740),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1084),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1131),
.B(n_830),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1087),
.A2(n_830),
.B(n_1008),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_SL g1237 ( 
.A1(n_1131),
.A2(n_830),
.B(n_942),
.C(n_920),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1131),
.A2(n_830),
.B(n_942),
.C(n_834),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1009),
.A2(n_965),
.A3(n_872),
.B(n_835),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1100),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1078),
.A2(n_1108),
.B(n_1127),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1131),
.B(n_830),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1078),
.A2(n_1108),
.B(n_1127),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1131),
.B(n_847),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_SL g1245 ( 
.A1(n_1131),
.A2(n_830),
.B(n_942),
.C(n_920),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_SL g1246 ( 
.A1(n_1131),
.A2(n_830),
.B(n_942),
.C(n_920),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1008),
.A2(n_830),
.B(n_1087),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1008),
.A2(n_830),
.B(n_1087),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_SL g1249 ( 
.A(n_1039),
.B(n_765),
.Y(n_1249)
);

AO21x1_ASAP7_75t_L g1250 ( 
.A1(n_1131),
.A2(n_830),
.B(n_942),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1084),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1100),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1131),
.B(n_830),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1131),
.B(n_830),
.Y(n_1254)
);

AO21x1_ASAP7_75t_L g1255 ( 
.A1(n_1131),
.A2(n_830),
.B(n_942),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1087),
.A2(n_830),
.B(n_1008),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1131),
.A2(n_830),
.B(n_1009),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1078),
.A2(n_1108),
.B(n_1127),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_SL g1259 ( 
.A1(n_1029),
.A2(n_1046),
.B(n_1071),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1131),
.B(n_830),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_987),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1087),
.A2(n_830),
.B(n_1008),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1098),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1100),
.Y(n_1264)
);

NAND3xp33_ASAP7_75t_L g1265 ( 
.A(n_1131),
.B(n_834),
.C(n_830),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1130),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1131),
.B(n_830),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1084),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1009),
.A2(n_965),
.A3(n_872),
.B(n_835),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1131),
.A2(n_830),
.B(n_1009),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1078),
.A2(n_1108),
.B(n_1127),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1131),
.A2(n_834),
.B(n_830),
.C(n_942),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1078),
.A2(n_1108),
.B(n_1127),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1078),
.A2(n_1108),
.B(n_1127),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1131),
.A2(n_830),
.B(n_1009),
.Y(n_1275)
);

INVx5_ASAP7_75t_L g1276 ( 
.A(n_1100),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1211),
.A2(n_1265),
.B1(n_1205),
.B2(n_1145),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1261),
.Y(n_1278)
);

INVx6_ASAP7_75t_L g1279 ( 
.A(n_1276),
.Y(n_1279)
);

INVx4_ASAP7_75t_L g1280 ( 
.A(n_1276),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_1215),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1265),
.A2(n_1205),
.B1(n_1145),
.B2(n_1177),
.Y(n_1282)
);

INVx4_ASAP7_75t_L g1283 ( 
.A(n_1276),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1163),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1220),
.B(n_1226),
.Y(n_1285)
);

AOI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1220),
.A2(n_1233),
.B1(n_1162),
.B2(n_1218),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1212),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1250),
.A2(n_1255),
.B1(n_1226),
.B2(n_1267),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1216),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1206),
.A2(n_1223),
.B1(n_1272),
.B2(n_1141),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1235),
.A2(n_1267),
.B1(n_1254),
.B2(n_1242),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1146),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1235),
.A2(n_1253),
.B1(n_1254),
.B2(n_1242),
.Y(n_1293)
);

CKINVDCx11_ASAP7_75t_R g1294 ( 
.A(n_1219),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1225),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1253),
.A2(n_1260),
.B1(n_1224),
.B2(n_1167),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_1266),
.Y(n_1297)
);

OAI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1244),
.A2(n_1249),
.B1(n_1260),
.B2(n_1171),
.Y(n_1298)
);

INVx3_ASAP7_75t_SL g1299 ( 
.A(n_1219),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1249),
.A2(n_1151),
.B1(n_1178),
.B2(n_1149),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1171),
.A2(n_1147),
.B1(n_1222),
.B2(n_1238),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1221),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1230),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1234),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_1188),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1203),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1251),
.Y(n_1307)
);

INVx6_ASAP7_75t_L g1308 ( 
.A(n_1192),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_1201),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1219),
.Y(n_1310)
);

INVx8_ASAP7_75t_L g1311 ( 
.A(n_1168),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1183),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1259),
.A2(n_1154),
.B1(n_1275),
.B2(n_1232),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1268),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_1160),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1185),
.A2(n_1193),
.B1(n_1169),
.B2(n_1170),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1232),
.A2(n_1275),
.B1(n_1270),
.B2(n_1257),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1190),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1189),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1208),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1139),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1182),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1186),
.A2(n_1257),
.B1(n_1270),
.B2(n_1181),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_1213),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1228),
.B(n_1138),
.Y(n_1325)
);

INVx6_ASAP7_75t_L g1326 ( 
.A(n_1168),
.Y(n_1326)
);

BUFx10_ASAP7_75t_L g1327 ( 
.A(n_1229),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1184),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_1157),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1169),
.A2(n_1139),
.B1(n_1187),
.B2(n_1134),
.Y(n_1330)
);

OAI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1186),
.A2(n_1152),
.B1(n_1173),
.B2(n_1175),
.Y(n_1331)
);

BUFx12f_ASAP7_75t_L g1332 ( 
.A(n_1229),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1198),
.Y(n_1333)
);

CKINVDCx11_ASAP7_75t_R g1334 ( 
.A(n_1229),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1199),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1155),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1180),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1175),
.A2(n_1159),
.B1(n_1179),
.B2(n_1174),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1197),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1197),
.Y(n_1340)
);

CKINVDCx11_ASAP7_75t_R g1341 ( 
.A(n_1240),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1156),
.A2(n_1165),
.B1(n_1194),
.B2(n_1179),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_SL g1343 ( 
.A1(n_1203),
.A2(n_1204),
.B1(n_1237),
.B2(n_1245),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1191),
.A2(n_1136),
.B1(n_1264),
.B2(n_1252),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1240),
.Y(n_1345)
);

OAI22x1_ASAP7_75t_L g1346 ( 
.A1(n_1166),
.A2(n_1207),
.B1(n_1143),
.B2(n_1246),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_1240),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1150),
.A2(n_1247),
.B1(n_1248),
.B2(n_1262),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1247),
.A2(n_1248),
.B1(n_1256),
.B2(n_1236),
.Y(n_1349)
);

INVx8_ASAP7_75t_L g1350 ( 
.A(n_1252),
.Y(n_1350)
);

OAI22xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1207),
.A2(n_1227),
.B1(n_1231),
.B2(n_1202),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1155),
.B(n_1142),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1252),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1263),
.Y(n_1354)
);

INVx6_ASAP7_75t_L g1355 ( 
.A(n_1264),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1195),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1137),
.A2(n_1172),
.B1(n_1135),
.B2(n_1144),
.Y(n_1357)
);

INVx6_ASAP7_75t_L g1358 ( 
.A(n_1214),
.Y(n_1358)
);

OAI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1200),
.A2(n_1196),
.B1(n_1142),
.B2(n_1155),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1142),
.A2(n_1158),
.B1(n_1195),
.B2(n_1176),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1172),
.A2(n_1140),
.B1(n_1273),
.B2(n_1271),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1209),
.A2(n_1274),
.B1(n_1258),
.B2(n_1243),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1210),
.A2(n_1217),
.B1(n_1241),
.B2(n_1158),
.Y(n_1363)
);

BUFx12f_ASAP7_75t_L g1364 ( 
.A(n_1176),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_SL g1365 ( 
.A1(n_1158),
.A2(n_1153),
.B1(n_1164),
.B2(n_1239),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1176),
.A2(n_1211),
.B1(n_1131),
.B2(n_1265),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1239),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1239),
.A2(n_1211),
.B1(n_1131),
.B2(n_1265),
.Y(n_1368)
);

OAI21xp33_ASAP7_75t_L g1369 ( 
.A1(n_1269),
.A2(n_834),
.B(n_1220),
.Y(n_1369)
);

BUFx10_ASAP7_75t_L g1370 ( 
.A(n_1269),
.Y(n_1370)
);

OAI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1269),
.A2(n_1220),
.B1(n_942),
.B2(n_830),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1211),
.A2(n_1131),
.B1(n_1265),
.B2(n_1205),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1177),
.A2(n_830),
.B1(n_942),
.B2(n_1220),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1205),
.B(n_1222),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1205),
.A2(n_1131),
.B1(n_830),
.B2(n_942),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1211),
.A2(n_1131),
.B1(n_1265),
.B2(n_1205),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1220),
.A2(n_834),
.B1(n_401),
.B2(n_830),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1211),
.A2(n_1131),
.B1(n_1265),
.B2(n_1205),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1149),
.B(n_1182),
.Y(n_1379)
);

BUFx12f_ASAP7_75t_L g1380 ( 
.A(n_1215),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1220),
.B(n_1177),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1148),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1216),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1215),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1220),
.A2(n_834),
.B1(n_401),
.B2(n_830),
.Y(n_1385)
);

BUFx8_ASAP7_75t_SL g1386 ( 
.A(n_1146),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1211),
.A2(n_1131),
.B1(n_1265),
.B2(n_1205),
.Y(n_1387)
);

INVx3_ASAP7_75t_SL g1388 ( 
.A(n_1266),
.Y(n_1388)
);

INVx4_ASAP7_75t_L g1389 ( 
.A(n_1276),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1261),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1177),
.A2(n_830),
.B1(n_942),
.B2(n_1220),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1220),
.A2(n_834),
.B1(n_401),
.B2(n_830),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1177),
.A2(n_740),
.B1(n_1205),
.B2(n_942),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1211),
.A2(n_1131),
.B1(n_1265),
.B2(n_1205),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1161),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1328),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1319),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1356),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1285),
.B(n_1277),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1318),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1311),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1349),
.A2(n_1348),
.B(n_1338),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1336),
.Y(n_1403)
);

AO21x2_ASAP7_75t_L g1404 ( 
.A1(n_1331),
.A2(n_1371),
.B(n_1374),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1336),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1357),
.A2(n_1348),
.B(n_1349),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1352),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1322),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1360),
.B(n_1367),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1339),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1340),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1357),
.A2(n_1338),
.B(n_1362),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1331),
.A2(n_1371),
.B(n_1374),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1370),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1370),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1291),
.B(n_1293),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1364),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1346),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1277),
.B(n_1366),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1366),
.B(n_1368),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1326),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1284),
.Y(n_1422)
);

AOI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1342),
.A2(n_1301),
.B(n_1290),
.Y(n_1423)
);

OAI21xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1317),
.A2(n_1313),
.B(n_1394),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1287),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1381),
.B(n_1368),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1295),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1303),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1304),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1326),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1393),
.A2(n_1282),
.B1(n_1373),
.B2(n_1391),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1307),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1317),
.A2(n_1313),
.B(n_1369),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1314),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1395),
.Y(n_1435)
);

CKINVDCx16_ASAP7_75t_R g1436 ( 
.A(n_1347),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1365),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1365),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1359),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1302),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1359),
.Y(n_1441)
);

AO21x1_ASAP7_75t_SL g1442 ( 
.A1(n_1372),
.A2(n_1394),
.B(n_1376),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1386),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1291),
.B(n_1293),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1351),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1282),
.B(n_1372),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1363),
.Y(n_1447)
);

AOI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1344),
.A2(n_1330),
.B(n_1316),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_1311),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1376),
.B(n_1378),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1333),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1362),
.A2(n_1288),
.B(n_1387),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1393),
.A2(n_1387),
.B1(n_1378),
.B2(n_1377),
.Y(n_1453)
);

AOI21xp33_ASAP7_75t_SL g1454 ( 
.A1(n_1385),
.A2(n_1392),
.B(n_1286),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1363),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1288),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1323),
.B(n_1296),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1298),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1298),
.B(n_1296),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1300),
.B(n_1379),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1335),
.Y(n_1461)
);

OR2x6_ASAP7_75t_L g1462 ( 
.A(n_1279),
.B(n_1280),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1323),
.B(n_1382),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1361),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1361),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1354),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1343),
.B(n_1325),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1343),
.B(n_1289),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1375),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1383),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1329),
.A2(n_1315),
.B1(n_1305),
.B2(n_1358),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1283),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1380),
.Y(n_1473)
);

OR2x6_ASAP7_75t_L g1474 ( 
.A(n_1283),
.B(n_1389),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1389),
.B(n_1337),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1320),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1436),
.B(n_1324),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1437),
.B(n_1312),
.Y(n_1478)
);

A2O1A1Ixp33_ASAP7_75t_L g1479 ( 
.A1(n_1454),
.A2(n_1320),
.B(n_1350),
.C(n_1353),
.Y(n_1479)
);

A2O1A1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1454),
.A2(n_1350),
.B(n_1310),
.C(n_1321),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1439),
.B(n_1441),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1415),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1400),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1453),
.A2(n_1309),
.B1(n_1358),
.B2(n_1308),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1438),
.B(n_1447),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1424),
.A2(n_1350),
.B(n_1390),
.C(n_1278),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1399),
.B(n_1390),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1415),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1410),
.Y(n_1489)
);

OR2x6_ASAP7_75t_L g1490 ( 
.A(n_1402),
.B(n_1358),
.Y(n_1490)
);

CKINVDCx8_ASAP7_75t_R g1491 ( 
.A(n_1436),
.Y(n_1491)
);

AOI211xp5_ASAP7_75t_L g1492 ( 
.A1(n_1457),
.A2(n_1299),
.B(n_1388),
.C(n_1306),
.Y(n_1492)
);

BUFx4f_ASAP7_75t_SL g1493 ( 
.A(n_1440),
.Y(n_1493)
);

BUFx4f_ASAP7_75t_SL g1494 ( 
.A(n_1440),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1399),
.B(n_1299),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1418),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1447),
.B(n_1355),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1431),
.A2(n_1308),
.B1(n_1345),
.B2(n_1355),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_SL g1499 ( 
.A1(n_1423),
.A2(n_1355),
.B(n_1327),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1455),
.B(n_1327),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1411),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1455),
.B(n_1388),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1460),
.B(n_1297),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1446),
.A2(n_1281),
.B(n_1292),
.Y(n_1504)
);

AO21x2_ASAP7_75t_L g1505 ( 
.A1(n_1402),
.A2(n_1332),
.B(n_1294),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1446),
.A2(n_1384),
.B(n_1334),
.Y(n_1506)
);

AO21x2_ASAP7_75t_L g1507 ( 
.A1(n_1445),
.A2(n_1341),
.B(n_1406),
.Y(n_1507)
);

AOI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1457),
.A2(n_1450),
.B1(n_1424),
.B2(n_1458),
.C(n_1419),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1439),
.B(n_1441),
.Y(n_1509)
);

INVx3_ASAP7_75t_L g1510 ( 
.A(n_1422),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1464),
.B(n_1465),
.Y(n_1511)
);

OR2x6_ASAP7_75t_L g1512 ( 
.A(n_1452),
.B(n_1412),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1459),
.A2(n_1450),
.B(n_1448),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1464),
.B(n_1465),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1408),
.B(n_1426),
.Y(n_1515)
);

BUFx12f_ASAP7_75t_L g1516 ( 
.A(n_1443),
.Y(n_1516)
);

AO21x2_ASAP7_75t_L g1517 ( 
.A1(n_1445),
.A2(n_1412),
.B(n_1404),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1459),
.A2(n_1448),
.B(n_1469),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1425),
.B(n_1427),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1404),
.A2(n_1413),
.B(n_1433),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1469),
.A2(n_1419),
.B(n_1458),
.Y(n_1521)
);

CKINVDCx6p67_ASAP7_75t_R g1522 ( 
.A(n_1476),
.Y(n_1522)
);

OAI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1452),
.A2(n_1426),
.B(n_1444),
.Y(n_1523)
);

OAI211xp5_ASAP7_75t_SL g1524 ( 
.A1(n_1468),
.A2(n_1476),
.B(n_1460),
.C(n_1466),
.Y(n_1524)
);

BUFx12f_ASAP7_75t_L g1525 ( 
.A(n_1473),
.Y(n_1525)
);

A2O1A1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1452),
.A2(n_1420),
.B(n_1468),
.C(n_1416),
.Y(n_1526)
);

OA21x2_ASAP7_75t_L g1527 ( 
.A1(n_1412),
.A2(n_1418),
.B(n_1398),
.Y(n_1527)
);

INVx4_ASAP7_75t_L g1528 ( 
.A(n_1474),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1404),
.A2(n_1413),
.B(n_1433),
.Y(n_1529)
);

O2A1O1Ixp33_ASAP7_75t_SL g1530 ( 
.A1(n_1417),
.A2(n_1466),
.B(n_1421),
.C(n_1470),
.Y(n_1530)
);

INVx4_ASAP7_75t_L g1531 ( 
.A(n_1474),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1515),
.B(n_1409),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1511),
.B(n_1407),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1517),
.B(n_1523),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1511),
.B(n_1407),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1514),
.B(n_1404),
.Y(n_1536)
);

AND2x4_ASAP7_75t_SL g1537 ( 
.A(n_1528),
.B(n_1462),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1514),
.B(n_1420),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1512),
.B(n_1413),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1503),
.B(n_1430),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1484),
.A2(n_1433),
.B1(n_1444),
.B2(n_1416),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1512),
.B(n_1413),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1512),
.B(n_1414),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1489),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1517),
.B(n_1409),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1526),
.B(n_1456),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1489),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1512),
.B(n_1433),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1531),
.B(n_1397),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1501),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1501),
.Y(n_1551)
);

NOR2xp67_ASAP7_75t_L g1552 ( 
.A(n_1520),
.B(n_1421),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1485),
.B(n_1456),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1484),
.A2(n_1508),
.B1(n_1491),
.B2(n_1490),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1517),
.B(n_1403),
.Y(n_1555)
);

OAI211xp5_ASAP7_75t_SL g1556 ( 
.A1(n_1518),
.A2(n_1471),
.B(n_1451),
.C(n_1435),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1490),
.A2(n_1442),
.B1(n_1467),
.B2(n_1463),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1527),
.B(n_1403),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1527),
.B(n_1405),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1527),
.B(n_1397),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1519),
.B(n_1397),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1519),
.B(n_1396),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1544),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1544),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1554),
.A2(n_1442),
.B1(n_1490),
.B2(n_1513),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1532),
.B(n_1496),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1547),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1547),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1543),
.B(n_1531),
.Y(n_1569)
);

INVxp67_ASAP7_75t_SL g1570 ( 
.A(n_1558),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1550),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1539),
.B(n_1485),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1560),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1551),
.Y(n_1574)
);

AOI222xp33_ASAP7_75t_L g1575 ( 
.A1(n_1554),
.A2(n_1521),
.B1(n_1504),
.B2(n_1506),
.C1(n_1524),
.C2(n_1463),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1543),
.B(n_1531),
.Y(n_1576)
);

AOI221xp5_ASAP7_75t_L g1577 ( 
.A1(n_1541),
.A2(n_1529),
.B1(n_1480),
.B2(n_1486),
.C(n_1479),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1542),
.B(n_1548),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1536),
.B(n_1483),
.Y(n_1579)
);

NAND4xp25_ASAP7_75t_L g1580 ( 
.A(n_1546),
.B(n_1492),
.C(n_1498),
.D(n_1495),
.Y(n_1580)
);

INVx1_ASAP7_75t_SL g1581 ( 
.A(n_1532),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1551),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1556),
.A2(n_1505),
.B1(n_1502),
.B2(n_1507),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1556),
.A2(n_1530),
.B(n_1505),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1558),
.Y(n_1585)
);

OAI33xp33_ASAP7_75t_L g1586 ( 
.A1(n_1541),
.A2(n_1487),
.A3(n_1509),
.B1(n_1481),
.B2(n_1434),
.B3(n_1428),
.Y(n_1586)
);

INVx4_ASAP7_75t_L g1587 ( 
.A(n_1537),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1557),
.A2(n_1491),
.B1(n_1494),
.B2(n_1493),
.Y(n_1588)
);

AO21x2_ASAP7_75t_L g1589 ( 
.A1(n_1552),
.A2(n_1507),
.B(n_1499),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1542),
.B(n_1502),
.Y(n_1590)
);

AOI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1546),
.A2(n_1467),
.B1(n_1461),
.B2(n_1429),
.C(n_1432),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1536),
.B(n_1510),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1543),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1548),
.B(n_1482),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1543),
.B(n_1549),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1560),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1548),
.B(n_1482),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1538),
.B(n_1488),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1545),
.A2(n_1522),
.B1(n_1509),
.B2(n_1481),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1538),
.B(n_1543),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1563),
.Y(n_1601)
);

NOR2xp67_ASAP7_75t_L g1602 ( 
.A(n_1593),
.B(n_1534),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1563),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1564),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1581),
.B(n_1553),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1581),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1600),
.B(n_1507),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1592),
.B(n_1545),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1579),
.B(n_1558),
.Y(n_1609)
);

NAND2x1_ASAP7_75t_SL g1610 ( 
.A(n_1569),
.B(n_1576),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1573),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1600),
.B(n_1561),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1592),
.B(n_1534),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1579),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1564),
.B(n_1559),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1591),
.B(n_1598),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1567),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1567),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1573),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1573),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1578),
.B(n_1561),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1568),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1591),
.B(n_1553),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1598),
.B(n_1533),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1568),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1571),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1578),
.B(n_1561),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1572),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1566),
.B(n_1533),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1572),
.B(n_1535),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1590),
.B(n_1594),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1566),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1590),
.B(n_1535),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1594),
.B(n_1562),
.Y(n_1634)
);

AOI321xp33_ASAP7_75t_L g1635 ( 
.A1(n_1565),
.A2(n_1477),
.A3(n_1540),
.B1(n_1500),
.B2(n_1497),
.C(n_1478),
.Y(n_1635)
);

AOI32xp33_ASAP7_75t_SL g1636 ( 
.A1(n_1616),
.A2(n_1570),
.A3(n_1575),
.B1(n_1582),
.B2(n_1574),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1610),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1623),
.A2(n_1583),
.B1(n_1577),
.B2(n_1584),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1606),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1601),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1601),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1606),
.B(n_1570),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1631),
.B(n_1595),
.Y(n_1643)
);

NOR2x1_ASAP7_75t_L g1644 ( 
.A(n_1602),
.B(n_1584),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1602),
.B(n_1569),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1603),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1611),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1603),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1604),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1604),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1617),
.Y(n_1651)
);

NOR2xp67_ASAP7_75t_L g1652 ( 
.A(n_1632),
.B(n_1587),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1613),
.B(n_1596),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1613),
.B(n_1596),
.Y(n_1654)
);

NAND4xp25_ASAP7_75t_L g1655 ( 
.A(n_1635),
.B(n_1575),
.C(n_1577),
.D(n_1580),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1608),
.B(n_1596),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1611),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1610),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1617),
.Y(n_1659)
);

O2A1O1Ixp33_ASAP7_75t_SL g1660 ( 
.A1(n_1635),
.A2(n_1588),
.B(n_1585),
.C(n_1599),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1618),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1614),
.B(n_1633),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1618),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1622),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1622),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1605),
.B(n_1630),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1631),
.B(n_1595),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1628),
.B(n_1595),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1625),
.Y(n_1669)
);

INVx2_ASAP7_75t_SL g1670 ( 
.A(n_1625),
.Y(n_1670)
);

OR2x2_ASAP7_75t_SL g1671 ( 
.A(n_1608),
.B(n_1585),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1626),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1611),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1607),
.B(n_1595),
.Y(n_1674)
);

OAI32xp33_ASAP7_75t_L g1675 ( 
.A1(n_1609),
.A2(n_1580),
.A3(n_1599),
.B1(n_1588),
.B2(n_1555),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1607),
.B(n_1597),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1624),
.B(n_1597),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1629),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1663),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1665),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1672),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1646),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1637),
.B(n_1626),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1655),
.B(n_1612),
.Y(n_1684)
);

A2O1A1Ixp33_ASAP7_75t_L g1685 ( 
.A1(n_1638),
.A2(n_1609),
.B(n_1552),
.C(n_1569),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1639),
.B(n_1612),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1671),
.B(n_1615),
.Y(n_1687)
);

BUFx2_ASAP7_75t_L g1688 ( 
.A(n_1658),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1646),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1658),
.B(n_1621),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1648),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1637),
.B(n_1621),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1678),
.B(n_1627),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1662),
.B(n_1627),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1671),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1670),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1660),
.B(n_1634),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1644),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1648),
.Y(n_1699)
);

CKINVDCx16_ASAP7_75t_R g1700 ( 
.A(n_1636),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1652),
.B(n_1634),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1670),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1642),
.Y(n_1703)
);

OR2x6_ASAP7_75t_L g1704 ( 
.A(n_1636),
.B(n_1462),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1649),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1666),
.B(n_1629),
.Y(n_1706)
);

NOR2x1_ASAP7_75t_L g1707 ( 
.A(n_1642),
.B(n_1649),
.Y(n_1707)
);

INVx1_ASAP7_75t_SL g1708 ( 
.A(n_1650),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1643),
.B(n_1593),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1645),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1677),
.B(n_1615),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1643),
.B(n_1593),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1667),
.B(n_1593),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1667),
.B(n_1619),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1690),
.B(n_1668),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1688),
.Y(n_1716)
);

A2O1A1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1698),
.A2(n_1675),
.B(n_1645),
.C(n_1668),
.Y(n_1717)
);

OAI211xp5_ASAP7_75t_L g1718 ( 
.A1(n_1695),
.A2(n_1675),
.B(n_1661),
.C(n_1651),
.Y(n_1718)
);

INVxp67_ASAP7_75t_SL g1719 ( 
.A(n_1707),
.Y(n_1719)
);

OAI21xp33_ASAP7_75t_L g1720 ( 
.A1(n_1704),
.A2(n_1645),
.B(n_1641),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1700),
.A2(n_1586),
.B1(n_1640),
.B2(n_1659),
.C(n_1669),
.Y(n_1721)
);

AOI21x1_ASAP7_75t_L g1722 ( 
.A1(n_1688),
.A2(n_1651),
.B(n_1650),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1682),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1700),
.B(n_1695),
.Y(n_1724)
);

INVxp67_ASAP7_75t_SL g1725 ( 
.A(n_1707),
.Y(n_1725)
);

OAI211xp5_ASAP7_75t_SL g1726 ( 
.A1(n_1684),
.A2(n_1661),
.B(n_1664),
.C(n_1669),
.Y(n_1726)
);

A2O1A1Ixp33_ASAP7_75t_SL g1727 ( 
.A1(n_1695),
.A2(n_1657),
.B(n_1647),
.C(n_1673),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1682),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1690),
.Y(n_1729)
);

OAI21xp33_ASAP7_75t_SL g1730 ( 
.A1(n_1704),
.A2(n_1674),
.B(n_1676),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1692),
.B(n_1674),
.Y(n_1731)
);

OAI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1704),
.A2(n_1664),
.B1(n_1653),
.B2(n_1654),
.C(n_1656),
.Y(n_1732)
);

AOI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1704),
.A2(n_1586),
.B1(n_1505),
.B2(n_1576),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1683),
.Y(n_1734)
);

NAND3xp33_ASAP7_75t_SL g1735 ( 
.A(n_1697),
.B(n_1710),
.C(n_1685),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1689),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1689),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1691),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1692),
.B(n_1676),
.Y(n_1739)
);

NOR2x1_ASAP7_75t_SL g1740 ( 
.A(n_1704),
.B(n_1589),
.Y(n_1740)
);

XNOR2x1_ASAP7_75t_L g1741 ( 
.A(n_1716),
.B(n_1687),
.Y(n_1741)
);

NAND3xp33_ASAP7_75t_L g1742 ( 
.A(n_1724),
.B(n_1717),
.C(n_1718),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1729),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1719),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1725),
.B(n_1702),
.Y(n_1745)
);

INVxp33_ASAP7_75t_L g1746 ( 
.A(n_1729),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1734),
.B(n_1702),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1715),
.B(n_1703),
.Y(n_1748)
);

AOI211xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1720),
.A2(n_1679),
.B(n_1680),
.C(n_1681),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1735),
.A2(n_1686),
.B1(n_1701),
.B2(n_1703),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1722),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1715),
.B(n_1701),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1722),
.Y(n_1753)
);

INVx2_ASAP7_75t_SL g1754 ( 
.A(n_1734),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1730),
.B(n_1703),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1739),
.B(n_1679),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1740),
.Y(n_1757)
);

INVxp67_ASAP7_75t_SL g1758 ( 
.A(n_1740),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1723),
.Y(n_1759)
);

AOI21xp33_ASAP7_75t_L g1760 ( 
.A1(n_1742),
.A2(n_1727),
.B(n_1732),
.Y(n_1760)
);

INVx1_ASAP7_75t_SL g1761 ( 
.A(n_1741),
.Y(n_1761)
);

OAI211xp5_ASAP7_75t_L g1762 ( 
.A1(n_1750),
.A2(n_1726),
.B(n_1733),
.C(n_1721),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1752),
.B(n_1731),
.Y(n_1763)
);

INVxp67_ASAP7_75t_SL g1764 ( 
.A(n_1741),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1744),
.A2(n_1731),
.B1(n_1739),
.B2(n_1681),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1749),
.B(n_1756),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1754),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1743),
.B(n_1680),
.Y(n_1768)
);

AOI21xp33_ASAP7_75t_L g1769 ( 
.A1(n_1746),
.A2(n_1696),
.B(n_1708),
.Y(n_1769)
);

OA21x2_ASAP7_75t_L g1770 ( 
.A1(n_1751),
.A2(n_1728),
.B(n_1723),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1748),
.B(n_1693),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1763),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1765),
.B(n_1746),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1761),
.B(n_1745),
.Y(n_1774)
);

NOR3xp33_ASAP7_75t_L g1775 ( 
.A(n_1764),
.B(n_1755),
.C(n_1753),
.Y(n_1775)
);

NOR3x1_ASAP7_75t_L g1776 ( 
.A(n_1766),
.B(n_1754),
.C(n_1755),
.Y(n_1776)
);

AND3x1_ASAP7_75t_L g1777 ( 
.A(n_1767),
.B(n_1768),
.C(n_1753),
.Y(n_1777)
);

AOI211x1_ASAP7_75t_L g1778 ( 
.A1(n_1762),
.A2(n_1759),
.B(n_1728),
.C(n_1736),
.Y(n_1778)
);

NAND3xp33_ASAP7_75t_L g1779 ( 
.A(n_1760),
.B(n_1751),
.C(n_1753),
.Y(n_1779)
);

NAND3xp33_ASAP7_75t_SL g1780 ( 
.A(n_1761),
.B(n_1757),
.C(n_1687),
.Y(n_1780)
);

AOI211x1_ASAP7_75t_SL g1781 ( 
.A1(n_1780),
.A2(n_1769),
.B(n_1757),
.C(n_1702),
.Y(n_1781)
);

O2A1O1Ixp33_ASAP7_75t_L g1782 ( 
.A1(n_1775),
.A2(n_1774),
.B(n_1779),
.C(n_1773),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_R g1783 ( 
.A(n_1772),
.B(n_1525),
.Y(n_1783)
);

A2O1A1Ixp33_ASAP7_75t_L g1784 ( 
.A1(n_1777),
.A2(n_1745),
.B(n_1758),
.C(n_1771),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1776),
.B(n_1516),
.Y(n_1785)
);

AOI221xp5_ASAP7_75t_L g1786 ( 
.A1(n_1782),
.A2(n_1778),
.B1(n_1745),
.B2(n_1747),
.C(n_1736),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1785),
.A2(n_1747),
.B1(n_1770),
.B2(n_1708),
.Y(n_1787)
);

O2A1O1Ixp5_ASAP7_75t_L g1788 ( 
.A1(n_1784),
.A2(n_1747),
.B(n_1737),
.C(n_1738),
.Y(n_1788)
);

AOI221xp5_ASAP7_75t_L g1789 ( 
.A1(n_1783),
.A2(n_1738),
.B1(n_1737),
.B2(n_1699),
.C(n_1691),
.Y(n_1789)
);

AOI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1781),
.A2(n_1699),
.B1(n_1705),
.B2(n_1683),
.C(n_1770),
.Y(n_1790)
);

OAI322xp33_ASAP7_75t_L g1791 ( 
.A1(n_1782),
.A2(n_1705),
.A3(n_1711),
.B1(n_1694),
.B2(n_1706),
.C1(n_1657),
.C2(n_1673),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1788),
.Y(n_1792)
);

NOR2x1_ASAP7_75t_L g1793 ( 
.A(n_1791),
.B(n_1683),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1787),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1786),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1789),
.Y(n_1796)
);

NOR3xp33_ASAP7_75t_L g1797 ( 
.A(n_1794),
.B(n_1790),
.C(n_1525),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1792),
.B(n_1683),
.Y(n_1798)
);

AND2x4_ASAP7_75t_L g1799 ( 
.A(n_1793),
.B(n_1714),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1798),
.A2(n_1795),
.B(n_1796),
.Y(n_1800)
);

AOI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1800),
.A2(n_1799),
.B1(n_1797),
.B2(n_1516),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1801),
.B(n_1711),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1801),
.B(n_1714),
.Y(n_1803)
);

AOI22x1_ASAP7_75t_L g1804 ( 
.A1(n_1802),
.A2(n_1647),
.B1(n_1712),
.B2(n_1709),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1803),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1805),
.Y(n_1806)
);

OAI21x1_ASAP7_75t_L g1807 ( 
.A1(n_1804),
.A2(n_1713),
.B(n_1712),
.Y(n_1807)
);

OAI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1806),
.A2(n_1713),
.B1(n_1709),
.B2(n_1654),
.Y(n_1808)
);

OA21x2_ASAP7_75t_L g1809 ( 
.A1(n_1808),
.A2(n_1807),
.B(n_1653),
.Y(n_1809)
);

XNOR2xp5_ASAP7_75t_L g1810 ( 
.A(n_1809),
.B(n_1401),
.Y(n_1810)
);

OAI221xp5_ASAP7_75t_R g1811 ( 
.A1(n_1810),
.A2(n_1656),
.B1(n_1522),
.B2(n_1620),
.C(n_1619),
.Y(n_1811)
);

AOI211xp5_ASAP7_75t_L g1812 ( 
.A1(n_1811),
.A2(n_1475),
.B(n_1449),
.C(n_1472),
.Y(n_1812)
);


endmodule