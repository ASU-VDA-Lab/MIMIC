module fake_jpeg_31634_n_72 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_72);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_72;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVxp67_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_25),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_0),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_13),
.B1(n_23),
.B2(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_10),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_3),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_37),
.C(n_25),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_27),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_35),
.B1(n_28),
.B2(n_26),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_47),
.A2(n_17),
.B1(n_21),
.B2(n_20),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_24),
.B1(n_19),
.B2(n_18),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_9),
.B1(n_5),
.B2(n_6),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_8),
.Y(n_64)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_42),
.B(n_6),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_59),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_4),
.C(n_7),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_61),
.C(n_63),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_4),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_8),
.C(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_62),
.Y(n_68)
);

A2O1A1O1Ixp25_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_69),
.B(n_59),
.C(n_67),
.D(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVxp33_ASAP7_75t_SL g71 ( 
.A(n_70),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_71),
.B(n_66),
.Y(n_72)
);


endmodule