module real_aes_8601_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_725;
wire n_119;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g177 ( .A1(n_0), .A2(n_178), .B(n_181), .C(n_185), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_1), .B(n_169), .Y(n_188) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_3), .B(n_179), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_4), .A2(n_138), .B(n_500), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_5), .A2(n_143), .B(n_146), .C(n_527), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_6), .A2(n_138), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_7), .B(n_169), .Y(n_506) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_8), .A2(n_171), .B(n_246), .Y(n_245) );
AND2x6_ASAP7_75t_L g143 ( .A(n_9), .B(n_144), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_10), .A2(n_143), .B(n_146), .C(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g540 ( .A(n_11), .Y(n_540) );
INVx1_ASAP7_75t_L g109 ( .A(n_12), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_12), .B(n_42), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_13), .B(n_184), .Y(n_529) );
INVx1_ASAP7_75t_L g164 ( .A(n_14), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_15), .B(n_179), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_16), .A2(n_180), .B(n_560), .C(n_562), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_17), .B(n_169), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_18), .B(n_158), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g145 ( .A1(n_19), .A2(n_146), .B(n_149), .C(n_157), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g547 ( .A1(n_20), .A2(n_183), .B(n_239), .C(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_21), .B(n_184), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_22), .A2(n_40), .B1(n_729), .B2(n_730), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_22), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_23), .B(n_184), .Y(n_514) );
CKINVDCx16_ASAP7_75t_R g474 ( .A(n_24), .Y(n_474) );
INVx1_ASAP7_75t_L g513 ( .A(n_25), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_26), .A2(n_146), .B(n_157), .C(n_249), .Y(n_248) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_27), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_28), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_29), .A2(n_79), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_29), .Y(n_127) );
INVx1_ASAP7_75t_L g491 ( .A(n_30), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_31), .A2(n_138), .B(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g141 ( .A(n_32), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_33), .A2(n_197), .B(n_198), .C(n_202), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_34), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_35), .A2(n_183), .B(n_503), .C(n_505), .Y(n_502) );
INVxp67_ASAP7_75t_L g492 ( .A(n_36), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_37), .B(n_251), .Y(n_250) );
CKINVDCx14_ASAP7_75t_R g501 ( .A(n_38), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_39), .A2(n_146), .B(n_157), .C(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_40), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_41), .A2(n_104), .B1(n_115), .B2(n_739), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_42), .B(n_109), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_43), .A2(n_185), .B(n_538), .C(n_539), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_44), .B(n_137), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_45), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_46), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_47), .B(n_179), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_48), .B(n_138), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_49), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_50), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_51), .A2(n_197), .B(n_202), .C(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g182 ( .A(n_52), .Y(n_182) );
INVx1_ASAP7_75t_L g225 ( .A(n_53), .Y(n_225) );
INVx1_ASAP7_75t_L g546 ( .A(n_54), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_55), .B(n_138), .Y(n_222) );
AOI222xp33_ASAP7_75t_L g456 ( .A1(n_56), .A2(n_457), .B1(n_724), .B2(n_725), .C1(n_731), .C2(n_736), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_57), .Y(n_166) );
CKINVDCx14_ASAP7_75t_R g536 ( .A(n_58), .Y(n_536) );
INVx1_ASAP7_75t_L g144 ( .A(n_59), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_60), .B(n_138), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_61), .B(n_169), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_62), .A2(n_156), .B(n_212), .C(n_214), .Y(n_211) );
INVx1_ASAP7_75t_L g163 ( .A(n_63), .Y(n_163) );
INVx1_ASAP7_75t_SL g504 ( .A(n_64), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_65), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_66), .B(n_179), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_67), .B(n_169), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_68), .B(n_180), .Y(n_236) );
INVx1_ASAP7_75t_L g477 ( .A(n_69), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_70), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_71), .B(n_151), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_72), .A2(n_146), .B(n_202), .C(n_265), .Y(n_264) );
CKINVDCx16_ASAP7_75t_R g210 ( .A(n_73), .Y(n_210) );
INVx1_ASAP7_75t_L g114 ( .A(n_74), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_75), .A2(n_138), .B(n_535), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_76), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_77), .A2(n_138), .B(n_557), .Y(n_556) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_78), .A2(n_124), .B1(n_125), .B2(n_128), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_78), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_79), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_80), .A2(n_137), .B(n_487), .Y(n_486) );
CKINVDCx16_ASAP7_75t_R g510 ( .A(n_81), .Y(n_510) );
INVx1_ASAP7_75t_L g558 ( .A(n_82), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_83), .B(n_154), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_84), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_84), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_85), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_86), .A2(n_138), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g561 ( .A(n_87), .Y(n_561) );
INVx2_ASAP7_75t_L g161 ( .A(n_88), .Y(n_161) );
INVx1_ASAP7_75t_L g528 ( .A(n_89), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_90), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_91), .B(n_184), .Y(n_237) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_92), .B(n_111), .C(n_112), .Y(n_110) );
OR2x2_ASAP7_75t_L g447 ( .A(n_92), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g460 ( .A(n_92), .B(n_449), .Y(n_460) );
INVx2_ASAP7_75t_L g462 ( .A(n_92), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_93), .A2(n_146), .B(n_202), .C(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_94), .B(n_138), .Y(n_195) );
INVx1_ASAP7_75t_L g199 ( .A(n_95), .Y(n_199) );
INVxp67_ASAP7_75t_L g215 ( .A(n_96), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_97), .B(n_171), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_98), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g232 ( .A(n_99), .Y(n_232) );
INVx1_ASAP7_75t_L g266 ( .A(n_100), .Y(n_266) );
INVx2_ASAP7_75t_L g549 ( .A(n_101), .Y(n_549) );
AND2x2_ASAP7_75t_L g227 ( .A(n_102), .B(n_160), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx5_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx9p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g739 ( .A(n_107), .Y(n_739) );
OR2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g449 ( .A(n_111), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_455), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_117), .B(n_451), .C(n_456), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_444), .B(n_451), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_129), .B1(n_442), .B2(n_443), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_123), .Y(n_442) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g443 ( .A(n_129), .Y(n_443) );
OAI22xp5_ASAP7_75t_SL g731 ( .A1(n_129), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
AND2x2_ASAP7_75t_SL g129 ( .A(n_130), .B(n_378), .Y(n_129) );
NOR5xp2_ASAP7_75t_L g130 ( .A(n_131), .B(n_309), .C(n_338), .D(n_358), .E(n_365), .Y(n_130) );
OAI211xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_189), .B(n_253), .C(n_296), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_133), .A2(n_381), .B1(n_383), .B2(n_384), .Y(n_380) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_168), .Y(n_133) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_134), .Y(n_256) );
AND2x4_ASAP7_75t_L g289 ( .A(n_134), .B(n_290), .Y(n_289) );
INVx5_ASAP7_75t_L g307 ( .A(n_134), .Y(n_307) );
AND2x2_ASAP7_75t_L g316 ( .A(n_134), .B(n_308), .Y(n_316) );
AND2x2_ASAP7_75t_L g328 ( .A(n_134), .B(n_193), .Y(n_328) );
AND2x2_ASAP7_75t_L g424 ( .A(n_134), .B(n_292), .Y(n_424) );
OR2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_165), .Y(n_134) );
AOI21xp5_ASAP7_75t_SL g135 ( .A1(n_136), .A2(n_145), .B(n_158), .Y(n_135) );
BUFx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
NAND2x1p5_ASAP7_75t_L g233 ( .A(n_139), .B(n_143), .Y(n_233) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g156 ( .A(n_140), .Y(n_156) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
INVx1_ASAP7_75t_L g240 ( .A(n_141), .Y(n_240) );
INVx1_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_142), .Y(n_152) );
INVx3_ASAP7_75t_L g180 ( .A(n_142), .Y(n_180) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_142), .Y(n_184) );
INVx1_ASAP7_75t_L g251 ( .A(n_142), .Y(n_251) );
BUFx3_ASAP7_75t_L g157 ( .A(n_143), .Y(n_157) );
INVx4_ASAP7_75t_SL g187 ( .A(n_143), .Y(n_187) );
INVx5_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx3_ASAP7_75t_L g186 ( .A(n_147), .Y(n_186) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_147), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_153), .B(n_155), .Y(n_149) );
INVx2_ASAP7_75t_L g154 ( .A(n_151), .Y(n_154) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx4_ASAP7_75t_L g213 ( .A(n_152), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_154), .A2(n_199), .B(n_200), .C(n_201), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_154), .A2(n_201), .B(n_225), .C(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_154), .A2(n_477), .B(n_478), .C(n_479), .Y(n_476) );
O2A1O1Ixp5_ASAP7_75t_L g527 ( .A1(n_154), .A2(n_479), .B(n_528), .C(n_529), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_155), .A2(n_179), .B(n_513), .C(n_514), .Y(n_512) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_156), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_159), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g167 ( .A(n_160), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_160), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_160), .A2(n_222), .B(n_223), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_160), .A2(n_233), .B(n_510), .C(n_511), .Y(n_509) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_160), .A2(n_534), .B(n_541), .Y(n_533) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AND2x2_ASAP7_75t_L g172 ( .A(n_161), .B(n_162), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_167), .A2(n_524), .B(n_530), .Y(n_523) );
INVx2_ASAP7_75t_L g290 ( .A(n_168), .Y(n_290) );
AND2x2_ASAP7_75t_L g308 ( .A(n_168), .B(n_262), .Y(n_308) );
AND2x2_ASAP7_75t_L g327 ( .A(n_168), .B(n_261), .Y(n_327) );
AND2x2_ASAP7_75t_L g367 ( .A(n_168), .B(n_307), .Y(n_367) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_173), .B(n_188), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_170), .B(n_204), .Y(n_203) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_170), .A2(n_231), .B(n_241), .Y(n_230) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_170), .A2(n_263), .B(n_271), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_170), .B(n_272), .Y(n_271) );
AO21x2_ASAP7_75t_L g472 ( .A1(n_170), .A2(n_473), .B(n_480), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_170), .B(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_170), .B(n_531), .Y(n_530) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_171), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_171), .A2(n_247), .B(n_248), .Y(n_246) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g243 ( .A(n_172), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_187), .Y(n_174) );
INVx2_ASAP7_75t_L g197 ( .A(n_176), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_176), .A2(n_187), .B(n_210), .C(n_211), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_SL g487 ( .A1(n_176), .A2(n_187), .B(n_488), .C(n_489), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g500 ( .A1(n_176), .A2(n_187), .B(n_501), .C(n_502), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_SL g535 ( .A1(n_176), .A2(n_187), .B(n_536), .C(n_537), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_SL g545 ( .A1(n_176), .A2(n_187), .B(n_546), .C(n_547), .Y(n_545) );
O2A1O1Ixp33_ASAP7_75t_SL g557 ( .A1(n_176), .A2(n_187), .B(n_558), .C(n_559), .Y(n_557) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_179), .B(n_215), .Y(n_214) );
OAI22xp33_ASAP7_75t_L g490 ( .A1(n_179), .A2(n_213), .B1(n_491), .B2(n_492), .Y(n_490) );
INVx5_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_180), .B(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_183), .B(n_504), .Y(n_503) );
INVx4_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g538 ( .A(n_184), .Y(n_538) );
INVx2_ASAP7_75t_L g479 ( .A(n_185), .Y(n_479) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_186), .Y(n_201) );
INVx1_ASAP7_75t_L g562 ( .A(n_186), .Y(n_562) );
INVx1_ASAP7_75t_L g202 ( .A(n_187), .Y(n_202) );
INVxp67_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_217), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AOI322xp5_ASAP7_75t_L g426 ( .A1(n_192), .A2(n_228), .A3(n_281), .B1(n_289), .B2(n_343), .C1(n_427), .C2(n_430), .Y(n_426) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_205), .Y(n_192) );
INVx5_ASAP7_75t_L g258 ( .A(n_193), .Y(n_258) );
AND2x2_ASAP7_75t_L g275 ( .A(n_193), .B(n_260), .Y(n_275) );
BUFx2_ASAP7_75t_L g353 ( .A(n_193), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_193), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g430 ( .A(n_193), .B(n_337), .Y(n_430) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_203), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_205), .B(n_219), .Y(n_284) );
INVx1_ASAP7_75t_L g311 ( .A(n_205), .Y(n_311) );
AND2x2_ASAP7_75t_L g324 ( .A(n_205), .B(n_244), .Y(n_324) );
AND2x2_ASAP7_75t_L g425 ( .A(n_205), .B(n_343), .Y(n_425) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g279 ( .A(n_206), .B(n_219), .Y(n_279) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_206), .Y(n_287) );
OR2x2_ASAP7_75t_L g294 ( .A(n_206), .B(n_244), .Y(n_294) );
AND2x2_ASAP7_75t_L g304 ( .A(n_206), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_206), .B(n_230), .Y(n_333) );
INVxp67_ASAP7_75t_L g357 ( .A(n_206), .Y(n_357) );
AND2x2_ASAP7_75t_L g364 ( .A(n_206), .B(n_228), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_206), .B(n_244), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_206), .B(n_229), .Y(n_390) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_216), .Y(n_206) );
OA21x2_ASAP7_75t_L g498 ( .A1(n_207), .A2(n_499), .B(n_506), .Y(n_498) );
OA21x2_ASAP7_75t_L g543 ( .A1(n_207), .A2(n_544), .B(n_550), .Y(n_543) );
OA21x2_ASAP7_75t_L g555 ( .A1(n_207), .A2(n_556), .B(n_563), .Y(n_555) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_212), .A2(n_266), .B(n_267), .C(n_268), .Y(n_265) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_213), .B(n_549), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_213), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_228), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_219), .B(n_245), .Y(n_334) );
OR2x2_ASAP7_75t_L g356 ( .A(n_219), .B(n_229), .Y(n_356) );
AND2x2_ASAP7_75t_L g369 ( .A(n_219), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_219), .B(n_324), .Y(n_375) );
OAI211xp5_ASAP7_75t_SL g379 ( .A1(n_219), .A2(n_380), .B(n_385), .C(n_394), .Y(n_379) );
AND2x2_ASAP7_75t_L g440 ( .A(n_219), .B(n_244), .Y(n_440) );
INVx5_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
OR2x2_ASAP7_75t_L g293 ( .A(n_220), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_220), .B(n_299), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_220), .B(n_288), .Y(n_300) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_220), .Y(n_302) );
OR2x2_ASAP7_75t_L g313 ( .A(n_220), .B(n_229), .Y(n_313) );
AND2x2_ASAP7_75t_SL g318 ( .A(n_220), .B(n_304), .Y(n_318) );
AND2x2_ASAP7_75t_L g343 ( .A(n_220), .B(n_229), .Y(n_343) );
AND2x2_ASAP7_75t_L g363 ( .A(n_220), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g401 ( .A(n_220), .B(n_228), .Y(n_401) );
OR2x2_ASAP7_75t_L g404 ( .A(n_220), .B(n_390), .Y(n_404) );
OR2x6_ASAP7_75t_L g220 ( .A(n_221), .B(n_227), .Y(n_220) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_244), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g347 ( .A1(n_229), .A2(n_348), .B(n_351), .C(n_357), .Y(n_347) );
INVx5_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_230), .B(n_244), .Y(n_278) );
AND2x2_ASAP7_75t_L g282 ( .A(n_230), .B(n_245), .Y(n_282) );
OR2x2_ASAP7_75t_L g288 ( .A(n_230), .B(n_244), .Y(n_288) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_234), .Y(n_231) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_233), .A2(n_474), .B(n_475), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_233), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_238), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_238), .A2(n_250), .B(n_252), .Y(n_249) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx2_ASAP7_75t_L g484 ( .A(n_243), .Y(n_484) );
INVx1_ASAP7_75t_SL g305 ( .A(n_244), .Y(n_305) );
OR2x2_ASAP7_75t_L g433 ( .A(n_244), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_273), .B(n_276), .C(n_285), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AOI31xp33_ASAP7_75t_L g358 ( .A1(n_255), .A2(n_359), .A3(n_361), .B(n_362), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_256), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_257), .B(n_289), .Y(n_295) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_258), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g315 ( .A(n_258), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g320 ( .A(n_258), .B(n_290), .Y(n_320) );
AND2x2_ASAP7_75t_L g330 ( .A(n_258), .B(n_289), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_258), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g350 ( .A(n_258), .B(n_307), .Y(n_350) );
AND2x2_ASAP7_75t_L g355 ( .A(n_258), .B(n_327), .Y(n_355) );
OR2x2_ASAP7_75t_L g374 ( .A(n_258), .B(n_260), .Y(n_374) );
OR2x2_ASAP7_75t_L g376 ( .A(n_258), .B(n_377), .Y(n_376) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_258), .Y(n_423) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g323 ( .A(n_260), .B(n_290), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_260), .B(n_307), .Y(n_346) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
BUFx2_ASAP7_75t_L g292 ( .A(n_262), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_270), .Y(n_263) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx3_ASAP7_75t_L g505 ( .A(n_269), .Y(n_505) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g383 ( .A(n_275), .B(n_307), .Y(n_383) );
AOI322xp5_ASAP7_75t_L g385 ( .A1(n_275), .A2(n_289), .A3(n_327), .B1(n_386), .B2(n_387), .C1(n_388), .C2(n_391), .Y(n_385) );
INVx1_ASAP7_75t_L g393 ( .A(n_275), .Y(n_393) );
NAND2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
INVx1_ASAP7_75t_SL g387 ( .A(n_277), .Y(n_387) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
OR2x2_ASAP7_75t_L g339 ( .A(n_278), .B(n_284), .Y(n_339) );
INVx1_ASAP7_75t_L g370 ( .A(n_278), .Y(n_370) );
INVx2_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OAI32xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_289), .A3(n_291), .B1(n_293), .B2(n_295), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AOI21xp33_ASAP7_75t_SL g325 ( .A1(n_288), .A2(n_303), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g340 ( .A(n_289), .Y(n_340) );
AND2x4_ASAP7_75t_L g337 ( .A(n_290), .B(n_307), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_290), .B(n_373), .Y(n_372) );
AOI322xp5_ASAP7_75t_L g402 ( .A1(n_291), .A2(n_318), .A3(n_337), .B1(n_370), .B2(n_403), .C1(n_405), .C2(n_406), .Y(n_402) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_291), .A2(n_368), .B1(n_432), .B2(n_433), .C(n_435), .Y(n_431) );
AND2x2_ASAP7_75t_L g319 ( .A(n_292), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g299 ( .A(n_294), .Y(n_299) );
OR2x2_ASAP7_75t_L g371 ( .A(n_294), .B(n_356), .Y(n_371) );
OAI31xp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_300), .A3(n_301), .B(n_306), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_297), .A2(n_330), .B1(n_331), .B2(n_335), .Y(n_329) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g342 ( .A(n_299), .B(n_343), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_301), .A2(n_342), .B1(n_395), .B2(n_398), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g384 ( .A(n_304), .B(n_353), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_304), .B(n_343), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_305), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g418 ( .A(n_305), .B(n_356), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_306), .A2(n_401), .B1(n_414), .B2(n_417), .Y(n_413) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx2_ASAP7_75t_L g322 ( .A(n_307), .Y(n_322) );
AND2x2_ASAP7_75t_L g405 ( .A(n_307), .B(n_327), .Y(n_405) );
OR2x2_ASAP7_75t_L g407 ( .A(n_307), .B(n_374), .Y(n_407) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_307), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_308), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_308), .B(n_353), .Y(n_361) );
OAI211xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_314), .B(n_317), .C(n_329), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B1(n_321), .B2(n_324), .C(n_325), .Y(n_317) );
INVxp67_ASAP7_75t_L g429 ( .A(n_320), .Y(n_429) );
INVx1_ASAP7_75t_L g396 ( .A(n_321), .Y(n_396) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x2_ASAP7_75t_L g360 ( .A(n_322), .B(n_327), .Y(n_360) );
INVx1_ASAP7_75t_L g377 ( .A(n_323), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_323), .B(n_350), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx1_ASAP7_75t_L g392 ( .A(n_327), .Y(n_392) );
AND2x2_ASAP7_75t_L g398 ( .A(n_327), .B(n_353), .Y(n_398) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_SL g386 ( .A(n_334), .Y(n_386) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_337), .B(n_373), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_341), .B2(n_344), .C(n_347), .Y(n_338) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g434 ( .A(n_343), .Y(n_434) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g352 ( .A(n_346), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_350), .B(n_409), .Y(n_408) );
AOI21xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B(n_356), .Y(n_351) );
OAI211xp5_ASAP7_75t_SL g399 ( .A1(n_354), .A2(n_400), .B(n_402), .C(n_408), .Y(n_399) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g411 ( .A(n_356), .Y(n_411) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI222xp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_368), .B1(n_371), .B2(n_372), .C1(n_375), .C2(n_376), .Y(n_365) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g441 ( .A(n_372), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_373), .B(n_416), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_373), .A2(n_420), .B1(n_422), .B2(n_425), .Y(n_419) );
INVx2_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
NOR4xp25_ASAP7_75t_L g378 ( .A(n_379), .B(n_399), .C(n_412), .D(n_431), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_381), .B(n_411), .Y(n_421) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g388 ( .A(n_386), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_389), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_419), .C(n_426), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx2_ASAP7_75t_L g428 ( .A(n_424), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
OAI21xp5_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_438), .B(n_441), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_443), .A2(n_458), .B1(n_461), .B2(n_463), .Y(n_457) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g454 ( .A(n_447), .Y(n_454) );
NOR2x2_ASAP7_75t_L g738 ( .A(n_448), .B(n_462), .Y(n_738) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g461 ( .A(n_449), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g732 ( .A(n_459), .Y(n_732) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g735 ( .A(n_461), .Y(n_735) );
INVx2_ASAP7_75t_L g733 ( .A(n_463), .Y(n_733) );
OR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_658), .Y(n_463) );
NAND5xp2_ASAP7_75t_L g464 ( .A(n_465), .B(n_587), .C(n_617), .D(n_638), .E(n_644), .Y(n_464) );
AOI221xp5_ASAP7_75t_SL g465 ( .A1(n_466), .A2(n_520), .B1(n_551), .B2(n_553), .C(n_564), .Y(n_465) );
INVxp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_517), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_495), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_SL g638 ( .A1(n_470), .A2(n_507), .B(n_639), .C(n_642), .Y(n_638) );
AND2x2_ASAP7_75t_L g708 ( .A(n_470), .B(n_508), .Y(n_708) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_482), .Y(n_470) );
AND2x2_ASAP7_75t_L g566 ( .A(n_471), .B(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g570 ( .A(n_471), .B(n_567), .Y(n_570) );
OR2x2_ASAP7_75t_L g596 ( .A(n_471), .B(n_508), .Y(n_596) );
AND2x2_ASAP7_75t_L g598 ( .A(n_471), .B(n_498), .Y(n_598) );
AND2x2_ASAP7_75t_L g616 ( .A(n_471), .B(n_497), .Y(n_616) );
INVx1_ASAP7_75t_L g649 ( .A(n_471), .Y(n_649) );
INVx2_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_L g519 ( .A(n_472), .Y(n_519) );
AND2x2_ASAP7_75t_L g552 ( .A(n_472), .B(n_498), .Y(n_552) );
AND2x2_ASAP7_75t_L g705 ( .A(n_472), .B(n_508), .Y(n_705) );
AND2x2_ASAP7_75t_L g586 ( .A(n_482), .B(n_496), .Y(n_586) );
OR2x2_ASAP7_75t_L g590 ( .A(n_482), .B(n_508), .Y(n_590) );
AND2x2_ASAP7_75t_L g615 ( .A(n_482), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g662 ( .A(n_482), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_482), .B(n_624), .Y(n_710) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_485), .B(n_493), .Y(n_482) );
INVx1_ASAP7_75t_L g568 ( .A(n_483), .Y(n_568) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OA21x2_ASAP7_75t_L g567 ( .A1(n_486), .A2(n_494), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OAI322xp33_ASAP7_75t_L g711 ( .A1(n_495), .A2(n_647), .A3(n_670), .B1(n_691), .B2(n_712), .C1(n_714), .C2(n_715), .Y(n_711) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_496), .B(n_567), .Y(n_714) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_507), .Y(n_496) );
AND2x2_ASAP7_75t_L g518 ( .A(n_497), .B(n_519), .Y(n_518) );
AND2x4_ASAP7_75t_L g583 ( .A(n_497), .B(n_508), .Y(n_583) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g624 ( .A(n_498), .B(n_508), .Y(n_624) );
AND2x2_ASAP7_75t_L g668 ( .A(n_498), .B(n_507), .Y(n_668) );
AND2x2_ASAP7_75t_L g551 ( .A(n_507), .B(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g569 ( .A(n_507), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_507), .B(n_598), .Y(n_722) );
INVx3_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g517 ( .A(n_508), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_508), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g636 ( .A(n_508), .B(n_567), .Y(n_636) );
AND2x2_ASAP7_75t_L g663 ( .A(n_508), .B(n_598), .Y(n_663) );
OR2x2_ASAP7_75t_L g719 ( .A(n_508), .B(n_570), .Y(n_719) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_515), .Y(n_508) );
INVx1_ASAP7_75t_SL g605 ( .A(n_517), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_518), .B(n_636), .Y(n_637) );
AND2x2_ASAP7_75t_L g671 ( .A(n_518), .B(n_661), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_518), .B(n_594), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_518), .B(n_716), .Y(n_715) );
OAI31xp33_ASAP7_75t_L g689 ( .A1(n_520), .A2(n_551), .A3(n_690), .B(n_692), .Y(n_689) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_532), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_521), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g672 ( .A(n_521), .B(n_607), .Y(n_672) );
OR2x2_ASAP7_75t_L g679 ( .A(n_521), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g691 ( .A(n_521), .B(n_580), .Y(n_691) );
CKINVDCx16_ASAP7_75t_R g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g625 ( .A(n_522), .B(n_626), .Y(n_625) );
BUFx3_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g553 ( .A(n_523), .B(n_554), .Y(n_553) );
INVx4_ASAP7_75t_L g574 ( .A(n_523), .Y(n_574) );
AND2x2_ASAP7_75t_L g611 ( .A(n_523), .B(n_555), .Y(n_611) );
AND2x2_ASAP7_75t_L g610 ( .A(n_532), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_SL g680 ( .A(n_532), .Y(n_680) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_542), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_533), .B(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g580 ( .A(n_533), .B(n_543), .Y(n_580) );
INVx2_ASAP7_75t_L g600 ( .A(n_533), .Y(n_600) );
AND2x2_ASAP7_75t_L g614 ( .A(n_533), .B(n_543), .Y(n_614) );
AND2x2_ASAP7_75t_L g621 ( .A(n_533), .B(n_577), .Y(n_621) );
BUFx3_ASAP7_75t_L g631 ( .A(n_533), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_533), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g576 ( .A(n_542), .Y(n_576) );
AND2x2_ASAP7_75t_L g584 ( .A(n_542), .B(n_574), .Y(n_584) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g554 ( .A(n_543), .B(n_555), .Y(n_554) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_543), .Y(n_608) );
INVx2_ASAP7_75t_SL g591 ( .A(n_552), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_552), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_552), .B(n_661), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_553), .B(n_631), .Y(n_684) );
INVx1_ASAP7_75t_SL g718 ( .A(n_553), .Y(n_718) );
INVx1_ASAP7_75t_SL g626 ( .A(n_554), .Y(n_626) );
INVx1_ASAP7_75t_SL g577 ( .A(n_555), .Y(n_577) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_555), .Y(n_588) );
OR2x2_ASAP7_75t_L g599 ( .A(n_555), .B(n_574), .Y(n_599) );
AND2x2_ASAP7_75t_L g613 ( .A(n_555), .B(n_574), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_555), .B(n_603), .Y(n_665) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_569), .B(n_571), .C(n_582), .Y(n_564) );
AOI31xp33_ASAP7_75t_L g681 ( .A1(n_565), .A2(n_682), .A3(n_683), .B(n_684), .Y(n_681) );
AND2x2_ASAP7_75t_L g654 ( .A(n_566), .B(n_583), .Y(n_654) );
BUFx3_ASAP7_75t_L g594 ( .A(n_567), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_567), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g630 ( .A(n_567), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_567), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g585 ( .A(n_570), .Y(n_585) );
OAI222xp33_ASAP7_75t_L g694 ( .A1(n_570), .A2(n_695), .B1(n_698), .B2(n_699), .C1(n_700), .C2(n_701), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_578), .Y(n_571) );
INVx1_ASAP7_75t_L g700 ( .A(n_572), .Y(n_700) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_574), .B(n_577), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_574), .B(n_600), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_574), .B(n_575), .Y(n_670) );
INVx1_ASAP7_75t_L g721 ( .A(n_574), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_575), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g723 ( .A(n_575), .Y(n_723) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx2_ASAP7_75t_L g603 ( .A(n_576), .Y(n_603) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_577), .Y(n_646) );
AOI32xp33_ASAP7_75t_L g582 ( .A1(n_578), .A2(n_583), .A3(n_584), .B1(n_585), .B2(n_586), .Y(n_582) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_580), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g657 ( .A(n_580), .Y(n_657) );
OR2x2_ASAP7_75t_L g698 ( .A(n_580), .B(n_599), .Y(n_698) );
INVx1_ASAP7_75t_L g634 ( .A(n_581), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_583), .B(n_594), .Y(n_619) );
INVx3_ASAP7_75t_L g628 ( .A(n_583), .Y(n_628) );
AOI322xp5_ASAP7_75t_L g644 ( .A1(n_583), .A2(n_628), .A3(n_645), .B1(n_647), .B2(n_650), .C1(n_654), .C2(n_655), .Y(n_644) );
AND2x2_ASAP7_75t_L g620 ( .A(n_584), .B(n_621), .Y(n_620) );
INVxp67_ASAP7_75t_L g697 ( .A(n_584), .Y(n_697) );
A2O1A1O1Ixp25_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B(n_592), .C(n_600), .D(n_601), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_588), .B(n_631), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
OAI221xp5_ASAP7_75t_L g601 ( .A1(n_590), .A2(n_602), .B1(n_605), .B2(n_606), .C(n_609), .Y(n_601) );
INVx1_ASAP7_75t_SL g716 ( .A(n_590), .Y(n_716) );
AOI21xp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_597), .B(n_599), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_594), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OAI221xp5_ASAP7_75t_SL g686 ( .A1(n_596), .A2(n_680), .B1(n_687), .B2(n_688), .C(n_689), .Y(n_686) );
OAI222xp33_ASAP7_75t_L g717 ( .A1(n_597), .A2(n_718), .B1(n_719), .B2(n_720), .C1(n_722), .C2(n_723), .Y(n_717) );
AND2x2_ASAP7_75t_L g675 ( .A(n_598), .B(n_661), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_598), .A2(n_613), .B(n_660), .Y(n_687) );
INVx1_ASAP7_75t_L g701 ( .A(n_598), .Y(n_701) );
INVx2_ASAP7_75t_SL g604 ( .A(n_599), .Y(n_604) );
AND2x2_ASAP7_75t_L g607 ( .A(n_600), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_SL g641 ( .A(n_603), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_603), .B(n_613), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_604), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_604), .B(n_614), .Y(n_643) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI21xp5_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_612), .B(n_615), .Y(n_609) );
INVx1_ASAP7_75t_SL g627 ( .A(n_611), .Y(n_627) );
AND2x2_ASAP7_75t_L g674 ( .A(n_611), .B(n_657), .Y(n_674) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g713 ( .A(n_613), .B(n_631), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_614), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g699 ( .A(n_615), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_620), .B1(n_622), .B2(n_629), .C(n_632), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_625), .B1(n_627), .B2(n_628), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_626), .A2(n_633), .B1(n_635), .B2(n_637), .Y(n_632) );
OR2x2_ASAP7_75t_L g703 ( .A(n_627), .B(n_631), .Y(n_703) );
OR2x2_ASAP7_75t_L g706 ( .A(n_627), .B(n_641), .Y(n_706) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g702 ( .A1(n_648), .A2(n_703), .B1(n_704), .B2(n_706), .C(n_707), .Y(n_702) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND3xp33_ASAP7_75t_SL g658 ( .A(n_659), .B(n_673), .C(n_685), .Y(n_658) );
AOI222xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_664), .B1(n_666), .B2(n_669), .C1(n_671), .C2(n_672), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_661), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g683 ( .A(n_663), .Y(n_683) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B1(n_676), .B2(n_678), .C(n_681), .Y(n_673) );
INVx1_ASAP7_75t_L g688 ( .A(n_674), .Y(n_688) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI21xp33_ASAP7_75t_L g707 ( .A1(n_678), .A2(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
NOR5xp2_ASAP7_75t_L g685 ( .A(n_686), .B(n_694), .C(n_702), .D(n_711), .E(n_717), .Y(n_685) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVxp67_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx3_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
endmodule