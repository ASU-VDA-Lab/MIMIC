module fake_jpeg_14299_n_100 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_100);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx4f_ASAP7_75t_SL g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_13),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_23),
.A2(n_24),
.B1(n_11),
.B2(n_17),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_13),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_0),
.C(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_5),
.Y(n_37)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_41),
.Y(n_54)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_18),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_24),
.B1(n_23),
.B2(n_30),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_37),
.B1(n_42),
.B2(n_16),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_50),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_49),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_17),
.B(n_16),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx24_ASAP7_75t_SL g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_52),
.B(n_14),
.Y(n_61)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_31),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_47),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_58),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_33),
.B1(n_37),
.B2(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_64),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_65),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_15),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_70),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_73),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_45),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_55),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_58),
.C(n_63),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_78),
.C(n_80),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_57),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_81),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_37),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_53),
.Y(n_82)
);

AOI221xp5_ASAP7_75t_L g85 ( 
.A1(n_82),
.A2(n_71),
.B1(n_53),
.B2(n_11),
.C(n_5),
.Y(n_85)
);

NOR2xp67_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_82),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_34),
.C(n_39),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_78),
.C(n_80),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_34),
.B1(n_39),
.B2(n_32),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_88),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_32),
.B1(n_11),
.B2(n_6),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_92),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_8),
.B(n_9),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_32),
.C(n_11),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_86),
.B1(n_83),
.B2(n_84),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g96 ( 
.A(n_93),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_97),
.A2(n_6),
.B(n_94),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_94),
.B(n_10),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_99),
.Y(n_100)
);


endmodule