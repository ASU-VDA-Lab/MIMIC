module fake_jpeg_8540_n_301 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_181;
wire n_38;
wire n_26;
wire n_28;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_17),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_30),
.B1(n_33),
.B2(n_20),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_27),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_18),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_18),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_59),
.Y(n_64)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_33),
.B1(n_21),
.B2(n_17),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_62),
.B(n_17),
.Y(n_77)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_55),
.Y(n_66)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_57),
.B(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_30),
.B1(n_20),
.B2(n_23),
.Y(n_76)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_21),
.B1(n_17),
.B2(n_18),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_22),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_86),
.Y(n_96)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_16),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_82),
.B1(n_19),
.B2(n_23),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_79),
.B1(n_46),
.B2(n_54),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_43),
.B(n_18),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_43),
.B1(n_19),
.B2(n_27),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_21),
.B1(n_20),
.B2(n_18),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_88),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_60),
.A2(n_21),
.B1(n_40),
.B2(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_48),
.B(n_24),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_68),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_32),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_34),
.C(n_40),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_105),
.Y(n_136)
);

AO21x1_ASAP7_75t_L g142 ( 
.A1(n_92),
.A2(n_24),
.B(n_25),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_67),
.A2(n_46),
.B1(n_54),
.B2(n_51),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_111),
.B1(n_85),
.B2(n_68),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_75),
.B(n_87),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_16),
.B1(n_25),
.B2(n_26),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_44),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_108),
.Y(n_139)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_110),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_67),
.A2(n_55),
.B1(n_40),
.B2(n_16),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_49),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_113),
.B(n_84),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_115),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_117),
.A2(n_123),
.B1(n_129),
.B2(n_137),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_87),
.B1(n_77),
.B2(n_66),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_64),
.B1(n_73),
.B2(n_78),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_119),
.A2(n_144),
.B1(n_26),
.B2(n_29),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_88),
.B1(n_73),
.B2(n_80),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_120),
.A2(n_134),
.B1(n_141),
.B2(n_115),
.Y(n_166)
);

XNOR2x2_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_80),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_121),
.A2(n_135),
.B(n_29),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_128),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_72),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_65),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_133),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_101),
.A2(n_87),
.B1(n_66),
.B2(n_65),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_98),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_66),
.B1(n_47),
.B2(n_24),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_26),
.B(n_31),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_109),
.A2(n_25),
.B1(n_31),
.B2(n_29),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_143),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_146),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_143),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_116),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_148),
.C(n_150),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_113),
.C(n_107),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_106),
.B(n_94),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_164),
.B(n_171),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_106),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_94),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_49),
.C(n_32),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_158),
.B(n_142),
.Y(n_183)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_166),
.Y(n_189)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_120),
.A2(n_131),
.B1(n_141),
.B2(n_134),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_167),
.A2(n_170),
.B1(n_161),
.B2(n_171),
.Y(n_202)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_169),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_105),
.B1(n_91),
.B2(n_31),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_119),
.A2(n_23),
.B(n_27),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_172),
.A2(n_174),
.B1(n_122),
.B2(n_129),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_173),
.A2(n_137),
.B1(n_125),
.B2(n_142),
.Y(n_184)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_117),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_175),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_135),
.B(n_140),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_179),
.B(n_164),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_140),
.B(n_125),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_191),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_123),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_193),
.C(n_196),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_167),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_198),
.B1(n_160),
.B2(n_148),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_157),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_154),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_158),
.B(n_144),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_28),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_28),
.Y(n_197)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_155),
.A2(n_32),
.B1(n_28),
.B2(n_93),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_156),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_32),
.Y(n_200)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_32),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_28),
.C(n_47),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_202),
.A2(n_187),
.B1(n_195),
.B2(n_173),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_213),
.Y(n_230)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_207),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_178),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_170),
.Y(n_209)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_186),
.A2(n_163),
.B1(n_149),
.B2(n_169),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_179),
.Y(n_235)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_163),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_218),
.C(n_221),
.Y(n_229)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_219),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_189),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_200),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_28),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_189),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_224),
.B1(n_225),
.B2(n_186),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_7),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_223),
.B(n_177),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_183),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_184),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_225)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_227),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_225),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_197),
.Y(n_231)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_217),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_234),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_185),
.C(n_196),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_238),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_237),
.B(n_242),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_181),
.Y(n_238)
);

XNOR2x1_ASAP7_75t_SL g239 ( 
.A(n_206),
.B(n_176),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_182),
.B(n_204),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_208),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_215),
.B(n_182),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_226),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_246),
.B(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_205),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_207),
.B(n_222),
.C(n_224),
.Y(n_250)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_251),
.A2(n_252),
.B(n_255),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_201),
.B1(n_212),
.B2(n_218),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_257),
.A2(n_229),
.B1(n_234),
.B2(n_236),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_221),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_230),
.C(n_257),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_244),
.B(n_241),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_268),
.B(n_263),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_260),
.B(n_264),
.Y(n_273)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_192),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_235),
.Y(n_265)
);

OAI21x1_ASAP7_75t_L g280 ( 
.A1(n_265),
.A2(n_267),
.B(n_9),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_249),
.B(n_229),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_266),
.A2(n_254),
.B(n_245),
.Y(n_272)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_270),
.B1(n_261),
.B2(n_259),
.Y(n_276)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_276),
.B(n_12),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_270),
.A2(n_250),
.B1(n_256),
.B2(n_243),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_274),
.A2(n_279),
.B(n_7),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_279),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_253),
.B1(n_192),
.B2(n_230),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_260),
.C(n_10),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_267),
.A2(n_192),
.B1(n_258),
.B2(n_213),
.Y(n_279)
);

A2O1A1O1Ixp25_ASAP7_75t_L g287 ( 
.A1(n_280),
.A2(n_12),
.B(n_14),
.C(n_5),
.D(n_6),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_285),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_283),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_10),
.C(n_14),
.Y(n_283)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_287),
.A2(n_277),
.B1(n_13),
.B2(n_6),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_5),
.B(n_6),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_288),
.A2(n_274),
.B(n_12),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_292),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_289),
.Y(n_294)
);

NAND4xp25_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_296),
.C(n_293),
.D(n_15),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_282),
.B(n_284),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_295),
.B(n_15),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_15),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_299),
.B(n_3),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_4),
.C(n_298),
.Y(n_301)
);


endmodule