module fake_jpeg_27575_n_313 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_313);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_23),
.B1(n_21),
.B2(n_12),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_45),
.B1(n_46),
.B2(n_14),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_23),
.B1(n_21),
.B2(n_12),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_25),
.A2(n_23),
.B1(n_21),
.B2(n_13),
.Y(n_46)
);

AO22x2_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_24),
.B1(n_33),
.B2(n_31),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_51),
.B1(n_54),
.B2(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_53),
.Y(n_68)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_45),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_23),
.B1(n_26),
.B2(n_21),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_59),
.B1(n_18),
.B2(n_13),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_34),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_18),
.B1(n_14),
.B2(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_61),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_63),
.Y(n_69)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_15),
.B1(n_22),
.B2(n_13),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_28),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_15),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_44),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_75),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_81),
.B1(n_42),
.B2(n_33),
.Y(n_106)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_80),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_48),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_65),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_56),
.B1(n_55),
.B2(n_48),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_86),
.A2(n_89),
.B1(n_103),
.B2(n_106),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_53),
.B(n_50),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_98),
.B(n_82),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_48),
.B1(n_51),
.B2(n_54),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_90),
.B(n_89),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_50),
.C(n_53),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_97),
.C(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_53),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_96),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_73),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_48),
.B1(n_51),
.B2(n_50),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_95),
.A2(n_105),
.B1(n_106),
.B2(n_93),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_51),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_18),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_17),
.B(n_14),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_82),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_58),
.B1(n_49),
.B2(n_42),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_62),
.C(n_43),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_81),
.A2(n_34),
.B(n_33),
.C(n_31),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_137),
.B(n_138),
.Y(n_140)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_110),
.B(n_112),
.Y(n_154)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_114),
.Y(n_152)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_79),
.A3(n_84),
.B1(n_18),
.B2(n_17),
.Y(n_117)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_121),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_79),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_119),
.B(n_27),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_84),
.Y(n_126)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_96),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_128),
.A2(n_135),
.B(n_136),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_97),
.Y(n_129)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_84),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_128),
.B1(n_127),
.B2(n_110),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_95),
.A2(n_78),
.B1(n_67),
.B2(n_77),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_90),
.A2(n_78),
.B1(n_67),
.B2(n_77),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_90),
.A2(n_67),
.B1(n_77),
.B2(n_14),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_87),
.B(n_31),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_91),
.A2(n_17),
.B(n_15),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_105),
.B(n_11),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_141),
.A2(n_156),
.B(n_135),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_105),
.C(n_37),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_124),
.C(n_135),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_105),
.B1(n_77),
.B2(n_13),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_70),
.B1(n_19),
.B2(n_20),
.Y(n_186)
);

OA21x2_ASAP7_75t_L g146 ( 
.A1(n_138),
.A2(n_105),
.B(n_70),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_159),
.Y(n_188)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_70),
.B1(n_12),
.B2(n_30),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_148),
.A2(n_155),
.B1(n_163),
.B2(n_112),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_151),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_126),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_125),
.B(n_19),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_162),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_70),
.B1(n_30),
.B2(n_27),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_119),
.Y(n_156)
);

BUFx24_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_161),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_108),
.B(n_37),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_116),
.A2(n_70),
.B1(n_30),
.B2(n_27),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_165),
.B(n_16),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_129),
.B(n_19),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_134),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_176),
.C(n_192),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_166),
.Y(n_175)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_169),
.C(n_142),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_115),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_198),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_123),
.B1(n_118),
.B2(n_111),
.Y(n_178)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

NAND2xp33_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_117),
.Y(n_180)
);

AOI221xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_143),
.B1(n_164),
.B2(n_157),
.C(n_146),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_145),
.A2(n_111),
.B1(n_108),
.B2(n_121),
.Y(n_181)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_182),
.A2(n_185),
.B(n_141),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_184),
.B(n_139),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_161),
.A2(n_132),
.B1(n_135),
.B2(n_137),
.Y(n_185)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_189),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_37),
.C(n_16),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_37),
.C(n_16),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_195),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_140),
.B(n_19),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_140),
.C(n_167),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_197),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_19),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_16),
.C(n_20),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_158),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_156),
.A2(n_20),
.B1(n_16),
.B2(n_2),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_201),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_208),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_190),
.A2(n_156),
.B(n_144),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_210),
.Y(n_230)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_154),
.Y(n_213)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_194),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_216),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_170),
.Y(n_217)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_139),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_157),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_246)
);

BUFx4f_ASAP7_75t_SL g223 ( 
.A(n_179),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_146),
.B1(n_155),
.B2(n_163),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_200),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_224),
.B(n_159),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_212),
.A2(n_174),
.B1(n_148),
.B2(n_196),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_220),
.B1(n_212),
.B2(n_225),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_176),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_239),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_173),
.C(n_192),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_238),
.C(n_218),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_242),
.B1(n_225),
.B2(n_205),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_219),
.A2(n_197),
.B1(n_184),
.B2(n_173),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_235),
.A2(n_245),
.B1(n_203),
.B2(n_204),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_195),
.C(n_193),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_198),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_226),
.A2(n_159),
.B1(n_186),
.B2(n_8),
.Y(n_242)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_243),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_219),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_245)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_246),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_248),
.B(n_0),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_249),
.A2(n_235),
.B1(n_237),
.B2(n_223),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_253),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_252),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_218),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_202),
.C(n_221),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_262),
.C(n_239),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_213),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_256),
.Y(n_264)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_257),
.A2(n_234),
.B1(n_241),
.B2(n_245),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_208),
.B(n_210),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_260),
.B(n_261),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_229),
.B1(n_237),
.B2(n_227),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_228),
.A2(n_207),
.B(n_214),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_217),
.B(n_203),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_223),
.C(n_215),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_263),
.A2(n_268),
.B1(n_7),
.B2(n_10),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_266),
.B(n_274),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_271),
.C(n_247),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_250),
.C(n_254),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_258),
.A2(n_261),
.B(n_251),
.Y(n_272)
);

OAI321xp33_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_7),
.A3(n_10),
.B1(n_9),
.B2(n_4),
.C(n_6),
.Y(n_285)
);

NOR2x1_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_236),
.Y(n_273)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_255),
.A2(n_236),
.B(n_8),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_7),
.Y(n_283)
);

OAI21x1_ASAP7_75t_L g276 ( 
.A1(n_272),
.A2(n_248),
.B(n_253),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_276),
.B(n_283),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_267),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_278),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_247),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_271),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_284),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_287),
.C(n_269),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_7),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

AO22x1_ASAP7_75t_L g288 ( 
.A1(n_285),
.A2(n_275),
.B1(n_2),
.B2(n_3),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_265),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_292),
.Y(n_297)
);

A2O1A1O1Ixp25_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_273),
.B(n_266),
.C(n_9),
.D(n_10),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_0),
.B(n_2),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_16),
.C(n_20),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_296),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_10),
.B1(n_9),
.B2(n_3),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_279),
.C(n_16),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_299),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_20),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_20),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_293),
.B(n_3),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_301),
.A2(n_290),
.B(n_288),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_305),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_304),
.Y(n_306)
);

OAI311xp33_ASAP7_75t_L g308 ( 
.A1(n_306),
.A2(n_297),
.A3(n_298),
.B1(n_299),
.C1(n_302),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_307),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.C1(n_0),
.C2(n_16),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_4),
.B(n_6),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_4),
.B(n_6),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_6),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_312),
.Y(n_313)
);


endmodule