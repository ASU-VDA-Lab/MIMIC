module real_jpeg_25543_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_1),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_1),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_1),
.B(n_75),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g163 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_85),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_1),
.B(n_26),
.C(n_27),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_1),
.B(n_65),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_1),
.A2(n_41),
.B1(n_184),
.B2(n_191),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g76 ( 
.A(n_4),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_5),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_5),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_5),
.A2(n_67),
.B1(n_88),
.B2(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_67),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_67),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_7),
.A2(n_54),
.B1(n_62),
.B2(n_64),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_54),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_9),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_10),
.A2(n_79),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_10),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_10),
.A2(n_62),
.B1(n_64),
.B2(n_89),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_89),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_89),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_13),
.A2(n_62),
.B1(n_64),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_13),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_69),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_69),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_39),
.Y(n_49)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_15),
.Y(n_111)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_15),
.Y(n_185)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_15),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_129),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_112),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_20),
.B(n_112),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_92),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_50),
.B1(n_90),
.B2(n_91),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_22),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_34),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_24),
.B(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_24),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_24),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_24),
.B(n_85),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_25),
.B(n_197),
.Y(n_196)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AO22x1_ASAP7_75t_L g65 ( 
.A1(n_31),
.A2(n_32),
.B1(n_60),
.B2(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_31),
.B(n_60),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_32),
.A2(n_61),
.A3(n_64),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_32),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_53),
.B(n_55),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_35),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_35),
.A2(n_144),
.B(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_35),
.A2(n_143),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_35),
.A2(n_142),
.B1(n_143),
.B2(n_164),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_45),
.B(n_48),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_41),
.A2(n_48),
.B(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_41),
.A2(n_174),
.B(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_41),
.A2(n_181),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_42),
.A2(n_46),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_42),
.B(n_49),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_42),
.A2(n_180),
.B1(n_182),
.B2(n_183),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g176 ( 
.A(n_44),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.C(n_71),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_51),
.A2(n_52),
.B1(n_56),
.B2(n_115),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_53),
.Y(n_156)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_66),
.B1(n_68),
.B2(n_70),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_68),
.B(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_57),
.A2(n_66),
.B1(n_70),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_58),
.A2(n_65),
.B1(n_126),
.B2(n_135),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_65),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_62),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_64),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_77),
.B(n_84),
.C(n_105),
.Y(n_104)
);

HAxp5_ASAP7_75t_SL g135 ( 
.A(n_62),
.B(n_85),
.CON(n_135),
.SN(n_135)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_76),
.C(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_65),
.B(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_71),
.B(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_74),
.B1(n_81),
.B2(n_86),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_75),
.B1(n_87),
.B2(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_80),
.B(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_85),
.B(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_103),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_106),
.B1(n_107),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_111),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.C(n_118),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_113),
.B(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_116),
.B(n_118),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_124),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_122),
.B1(n_123),
.B2(n_149),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_119),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_208),
.B(n_212),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_158),
.B(n_207),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_145),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_132),
.B(n_145),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.C(n_141),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_133),
.B(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_176),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_140),
.B(n_141),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_146),
.B(n_153),
.C(n_157),
.Y(n_209)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_157),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_152),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_202),
.B(n_206),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_177),
.B(n_201),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_161),
.B(n_167),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_165),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_173),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_172),
.C(n_173),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_187),
.B(n_200),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_186),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_186),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_194),
.B(n_199),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_189),
.B(n_190),
.Y(n_199)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_203),
.B(n_204),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_209),
.B(n_210),
.Y(n_212)
);


endmodule