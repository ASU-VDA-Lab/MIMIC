module fake_netlist_1_422_n_16 (n_1, n_2, n_0, n_16);
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
CKINVDCx11_ASAP7_75t_R g3 ( .A(n_0), .Y(n_3) );
INVx2_ASAP7_75t_SL g4 ( .A(n_1), .Y(n_4) );
OAI21x1_ASAP7_75t_L g5 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_5) );
AND3x4_ASAP7_75t_L g6 ( .A(n_3), .B(n_0), .C(n_1), .Y(n_6) );
INVx2_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
HB1xp67_ASAP7_75t_L g8 ( .A(n_6), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_7), .B(n_4), .Y(n_9) );
AND2x4_ASAP7_75t_SL g10 ( .A(n_8), .B(n_6), .Y(n_10) );
OAI21xp5_ASAP7_75t_L g11 ( .A1(n_9), .A2(n_4), .B(n_3), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_10), .B(n_0), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
O2A1O1Ixp33_ASAP7_75t_L g14 ( .A1(n_11), .A2(n_1), .B(n_2), .C(n_8), .Y(n_14) );
INVx1_ASAP7_75t_SL g15 ( .A(n_13), .Y(n_15) );
OAI22xp5_ASAP7_75t_L g16 ( .A1(n_15), .A2(n_2), .B1(n_14), .B2(n_11), .Y(n_16) );
endmodule