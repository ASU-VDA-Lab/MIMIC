module fake_jpeg_17676_n_42 (n_3, n_2, n_1, n_0, n_4, n_5, n_42);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx5_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx4_ASAP7_75t_SL g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx10_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_4),
.Y(n_11)
);

AND2x2_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_3),
.Y(n_12)
);

CKINVDCx12_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_11),
.B(n_5),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_0),
.C(n_1),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_15),
.A2(n_3),
.B(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_19),
.Y(n_21)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_20),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_3),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_12),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_16),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_15),
.A2(n_8),
.B1(n_12),
.B2(n_10),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_6),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_6),
.C(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.C(n_23),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_36),
.A2(n_34),
.B1(n_32),
.B2(n_21),
.Y(n_38)
);

INVxp67_ASAP7_75t_SL g40 ( 
.A(n_38),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_28),
.B(n_4),
.Y(n_39)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_35),
.B(n_39),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_36),
.C(n_26),
.Y(n_42)
);


endmodule