module fake_jpeg_28640_n_532 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_532);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_532;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_55),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_28),
.B(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_57),
.B(n_81),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_62),
.Y(n_151)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_31),
.B(n_8),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_96),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_70),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_73),
.Y(n_148)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_28),
.B(n_8),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_83),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_89),
.Y(n_166)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_101),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_24),
.B(n_7),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_102),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_32),
.B(n_7),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_104),
.Y(n_109)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_106),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_25),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

INVx6_ASAP7_75t_SL g157 ( 
.A(n_107),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_30),
.B1(n_52),
.B2(n_51),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_118),
.A2(n_44),
.B1(n_30),
.B2(n_75),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_69),
.B(n_53),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_122),
.B(n_124),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_53),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_60),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_128),
.B(n_137),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_60),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_76),
.B(n_50),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_141),
.B(n_142),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_78),
.B(n_50),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_37),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_143),
.B(n_146),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_100),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_37),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_165),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_56),
.A2(n_43),
.B1(n_32),
.B2(n_40),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_20),
.B1(n_25),
.B2(n_27),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_58),
.B(n_40),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_163),
.B(n_156),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_61),
.B(n_43),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_66),
.B(n_20),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_35),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_170),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_171),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_112),
.Y(n_174)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_175),
.A2(n_198),
.B1(n_42),
.B2(n_154),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_27),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_176),
.B(n_183),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_157),
.A2(n_36),
.B1(n_26),
.B2(n_38),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_177),
.A2(n_184),
.B1(n_215),
.B2(n_217),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_108),
.A2(n_42),
.B(n_12),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_178),
.A2(n_181),
.B(n_42),
.Y(n_225)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_180),
.Y(n_241)
);

O2A1O1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_42),
.B(n_45),
.C(n_36),
.Y(n_181)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_120),
.B(n_144),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_149),
.A2(n_45),
.B1(n_41),
.B2(n_38),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_111),
.Y(n_185)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_186),
.Y(n_258)
);

AOI21xp33_ASAP7_75t_L g189 ( 
.A1(n_114),
.A2(n_109),
.B(n_120),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_189),
.B(n_166),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_113),
.A2(n_93),
.B1(n_87),
.B2(n_86),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_191),
.A2(n_203),
.B1(n_206),
.B2(n_213),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_110),
.Y(n_192)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_138),
.Y(n_194)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_194),
.Y(n_244)
);

CKINVDCx12_ASAP7_75t_R g195 ( 
.A(n_110),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_207),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_131),
.Y(n_196)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_196),
.Y(n_245)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_117),
.Y(n_199)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

BUFx24_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_201),
.Y(n_255)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_135),
.Y(n_202)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_202),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_133),
.A2(n_85),
.B1(n_80),
.B2(n_73),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_72),
.C(n_70),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_204),
.B(n_218),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_133),
.A2(n_67),
.B1(n_41),
.B2(n_26),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_209),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_211),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_125),
.B(n_52),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_121),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_214),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_148),
.A2(n_30),
.B1(n_51),
.B2(n_35),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_121),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_131),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_216),
.B(n_221),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_147),
.A2(n_52),
.B1(n_51),
.B2(n_35),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_126),
.B(n_44),
.C(n_51),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_115),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_219),
.B(n_220),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_123),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_132),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_148),
.B(n_44),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_134),
.Y(n_265)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_130),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_223),
.B(n_224),
.Y(n_233)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_169),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_225),
.A2(n_172),
.B1(n_158),
.B2(n_193),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_226),
.B(n_260),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_178),
.A2(n_118),
.B(n_140),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_232),
.B(n_261),
.C(n_181),
.Y(n_271)
);

AND2x4_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_42),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_256),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_183),
.B(n_51),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_239),
.B(n_187),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_176),
.A2(n_132),
.B1(n_167),
.B2(n_145),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_243),
.A2(n_246),
.B1(n_266),
.B2(n_209),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_204),
.A2(n_205),
.B1(n_174),
.B2(n_145),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_173),
.B(n_169),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_188),
.B(n_127),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_265),
.B(n_223),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_198),
.A2(n_167),
.B1(n_218),
.B2(n_154),
.Y(n_266)
);

OAI32xp33_ASAP7_75t_L g267 ( 
.A1(n_200),
.A2(n_134),
.A3(n_130),
.B1(n_52),
.B2(n_44),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_207),
.Y(n_280)
);

INVx13_ASAP7_75t_L g268 ( 
.A(n_242),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_268),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_269),
.A2(n_270),
.B1(n_253),
.B2(n_257),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_199),
.B1(n_202),
.B2(n_194),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_271),
.B(n_232),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_233),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_276),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_273),
.B(n_289),
.Y(n_319)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_275),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_234),
.Y(n_276)
);

INVx13_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_277),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_235),
.B(n_208),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_278),
.B(n_283),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_280),
.A2(n_294),
.B1(n_243),
.B2(n_250),
.Y(n_306)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

INVx13_ASAP7_75t_L g282 ( 
.A(n_228),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_290),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_235),
.B(n_224),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_229),
.Y(n_284)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_284),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_229),
.B(n_214),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_285),
.B(n_287),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_286),
.Y(n_309)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_244),
.Y(n_288)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_288),
.Y(n_324)
);

OAI221xp5_ASAP7_75t_L g289 ( 
.A1(n_226),
.A2(n_201),
.B1(n_192),
.B2(n_182),
.C(n_207),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_251),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_239),
.B(n_179),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_292),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_225),
.B(n_23),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_236),
.B(n_192),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_293),
.B(n_300),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_256),
.A2(n_119),
.B1(n_153),
.B2(n_164),
.Y(n_294)
);

INVx4_ASAP7_75t_SL g295 ( 
.A(n_230),
.Y(n_295)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_295),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_255),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_296),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_255),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_297),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_249),
.A2(n_220),
.B1(n_219),
.B2(n_129),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_298),
.A2(n_299),
.B(n_301),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_230),
.A2(n_129),
.B1(n_127),
.B2(n_197),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_238),
.B(n_164),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_231),
.A2(n_130),
.B1(n_123),
.B2(n_134),
.Y(n_301)
);

OR2x6_ASAP7_75t_L g302 ( 
.A(n_238),
.B(n_201),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_264),
.CI(n_238),
.CON(n_311),
.SN(n_311)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_227),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_237),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_264),
.C(n_261),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_304),
.B(n_317),
.C(n_302),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_306),
.A2(n_334),
.B1(n_309),
.B2(n_286),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_292),
.A2(n_264),
.B(n_246),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_310),
.A2(n_328),
.B(n_329),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_302),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_315),
.B(n_331),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_271),
.B(n_238),
.C(n_231),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_321),
.A2(n_326),
.B1(n_294),
.B2(n_272),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_274),
.B(n_267),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_323),
.B(n_274),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_269),
.A2(n_245),
.B1(n_180),
.B2(n_186),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_292),
.A2(n_263),
.B(n_250),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_302),
.A2(n_252),
.B(n_262),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_278),
.B(n_257),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_283),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_279),
.A2(n_252),
.B1(n_258),
.B2(n_245),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_284),
.Y(n_336)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_336),
.Y(n_354)
);

AND2x6_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_302),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_337),
.A2(n_348),
.B(n_287),
.Y(n_395)
);

CKINVDCx14_ASAP7_75t_R g386 ( 
.A(n_338),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_346),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_325),
.A2(n_302),
.B(n_279),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_340),
.B(n_341),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_290),
.Y(n_342)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_342),
.Y(n_389)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_320),
.Y(n_343)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_343),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_335),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_344),
.B(n_345),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_318),
.B(n_303),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_318),
.B(n_333),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_357),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_311),
.B(n_302),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_349),
.A2(n_361),
.B1(n_360),
.B2(n_338),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_335),
.Y(n_350)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_350),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_304),
.B(n_291),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_351),
.B(n_356),
.C(n_317),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_321),
.A2(n_323),
.B1(n_326),
.B2(n_279),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_355),
.B(n_365),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_316),
.B(n_273),
.Y(n_357)
);

MAJx2_ASAP7_75t_L g358 ( 
.A(n_304),
.B(n_279),
.C(n_300),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_325),
.Y(n_383)
);

AOI22x1_ASAP7_75t_L g359 ( 
.A1(n_310),
.A2(n_286),
.B1(n_289),
.B2(n_280),
.Y(n_359)
);

AO21x2_ASAP7_75t_L g392 ( 
.A1(n_359),
.A2(n_270),
.B(n_299),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_322),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_360),
.B(n_361),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_322),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_319),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_362),
.B(n_363),
.Y(n_399)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_314),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_327),
.B(n_293),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_364),
.B(n_368),
.Y(n_390)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_314),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_329),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_366),
.B(n_367),
.Y(n_398)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_336),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_312),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_370),
.C(n_374),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_351),
.B(n_356),
.C(n_353),
.Y(n_370)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_343),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_372),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_315),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_384),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_317),
.C(n_311),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_352),
.Y(n_375)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_375),
.Y(n_409)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_362),
.Y(n_377)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_377),
.Y(n_422)
);

OAI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_359),
.A2(n_306),
.B1(n_305),
.B2(n_328),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_379),
.A2(n_387),
.B1(n_355),
.B2(n_341),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_354),
.A2(n_305),
.B1(n_295),
.B2(n_298),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_380),
.A2(n_385),
.B1(n_346),
.B2(n_330),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_311),
.C(n_331),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_381),
.B(n_313),
.C(n_281),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_383),
.B(n_324),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_345),
.B(n_332),
.Y(n_384)
);

OAI21xp33_ASAP7_75t_SL g387 ( 
.A1(n_359),
.A2(n_332),
.B(n_334),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_392),
.A2(n_395),
.B(n_400),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_347),
.B(n_277),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_394),
.B(n_397),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_339),
.B(n_277),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_366),
.A2(n_301),
.B(n_330),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_401),
.A2(n_421),
.B1(n_428),
.B2(n_392),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_367),
.Y(n_403)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_403),
.Y(n_437)
);

OAI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_377),
.A2(n_365),
.B1(n_363),
.B2(n_354),
.Y(n_404)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_404),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_382),
.A2(n_337),
.B(n_348),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_405),
.B(n_424),
.Y(n_429)
);

MAJx2_ASAP7_75t_L g408 ( 
.A(n_374),
.B(n_348),
.C(n_341),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_408),
.B(n_425),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_340),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_410),
.B(n_417),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_391),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_412),
.B(n_418),
.Y(n_440)
);

XNOR2x1_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_392),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_398),
.A2(n_368),
.B(n_307),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_414),
.A2(n_400),
.B(n_396),
.Y(n_445)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_371),
.Y(n_415)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_415),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_386),
.B(n_307),
.Y(n_416)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_416),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_370),
.B(n_285),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_398),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_384),
.B(n_237),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_419),
.B(n_420),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_388),
.B(n_312),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_392),
.A2(n_324),
.B1(n_313),
.B2(n_320),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_390),
.B(n_385),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_426),
.B(n_376),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_369),
.B(n_288),
.C(n_275),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_427),
.B(n_381),
.C(n_373),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_392),
.A2(n_320),
.B1(n_295),
.B2(n_258),
.Y(n_428)
);

XOR2x1_ASAP7_75t_L g430 ( 
.A(n_405),
.B(n_395),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_430),
.B(n_432),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_431),
.B(n_433),
.C(n_438),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_427),
.B(n_382),
.C(n_378),
.Y(n_433)
);

XNOR2x1_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_378),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_434),
.B(n_268),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_435),
.A2(n_428),
.B1(n_421),
.B2(n_418),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_449),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_411),
.B(n_382),
.C(n_393),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_415),
.A2(n_389),
.B1(n_376),
.B2(n_396),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_444),
.A2(n_407),
.B1(n_410),
.B2(n_402),
.Y(n_459)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_445),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_411),
.B(n_372),
.C(n_240),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_451),
.C(n_228),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_406),
.B(n_262),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_406),
.B(n_254),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_450),
.B(n_425),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_240),
.C(n_254),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_429),
.B(n_409),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_452),
.B(n_453),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_446),
.B(n_416),
.Y(n_453)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_455),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_442),
.A2(n_401),
.B1(n_423),
.B2(n_403),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_456),
.B(n_458),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_457),
.B(n_468),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_448),
.A2(n_420),
.B1(n_414),
.B2(n_422),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_459),
.B(n_282),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_443),
.A2(n_407),
.B1(n_408),
.B2(n_241),
.Y(n_460)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_460),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_440),
.A2(n_241),
.B1(n_248),
.B2(n_247),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_461),
.A2(n_466),
.B(n_450),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_436),
.B(n_244),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_465),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_447),
.Y(n_466)
);

NOR3xp33_ASAP7_75t_SL g467 ( 
.A(n_430),
.B(n_268),
.C(n_282),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_467),
.B(n_470),
.Y(n_485)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_437),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_469),
.A2(n_438),
.B(n_431),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_471),
.A2(n_475),
.B(n_479),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_455),
.A2(n_432),
.B1(n_434),
.B2(n_449),
.Y(n_473)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_473),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_463),
.A2(n_433),
.B(n_451),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_457),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_462),
.B(n_439),
.C(n_441),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_439),
.C(n_441),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_480),
.A2(n_481),
.B(n_482),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_241),
.C(n_247),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_248),
.C(n_185),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_486),
.B(n_44),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_454),
.B(n_221),
.C(n_215),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_487),
.A2(n_166),
.B(n_190),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_454),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_490),
.B(n_494),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_485),
.B(n_463),
.Y(n_491)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_491),
.Y(n_508)
);

NOR2xp67_ASAP7_75t_L g492 ( 
.A(n_483),
.B(n_467),
.Y(n_492)
);

NOR2x1_ASAP7_75t_L g511 ( 
.A(n_492),
.B(n_6),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_480),
.A2(n_475),
.B(n_484),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_493),
.A2(n_496),
.B(n_6),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_474),
.A2(n_468),
.B(n_156),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_495),
.A2(n_482),
.B(n_487),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_485),
.B(n_196),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_498),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_476),
.B(n_52),
.Y(n_498)
);

FAx1_ASAP7_75t_SL g499 ( 
.A(n_476),
.B(n_119),
.CI(n_11),
.CON(n_499),
.SN(n_499)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_499),
.A2(n_500),
.B1(n_501),
.B2(n_486),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_477),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_502),
.B(n_472),
.C(n_481),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_505),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_491),
.A2(n_473),
.B(n_472),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_504),
.A2(n_507),
.B(n_513),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_506),
.B(n_15),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_488),
.B(n_0),
.C(n_1),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_SL g514 ( 
.A1(n_511),
.A2(n_496),
.B1(n_499),
.B2(n_2),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_512),
.A2(n_6),
.B(n_16),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_489),
.A2(n_6),
.B(n_16),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_514),
.A2(n_509),
.B(n_4),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_520),
.Y(n_523)
);

AOI322xp5_ASAP7_75t_L g517 ( 
.A1(n_508),
.A2(n_5),
.A3(n_15),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_17),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_517),
.B(n_518),
.Y(n_521)
);

AOI322xp5_ASAP7_75t_L g518 ( 
.A1(n_511),
.A2(n_5),
.A3(n_13),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_15),
.Y(n_518)
);

A2O1A1O1Ixp25_ASAP7_75t_L g522 ( 
.A1(n_519),
.A2(n_510),
.B(n_504),
.C(n_503),
.D(n_507),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_522),
.A2(n_524),
.B(n_515),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_525),
.B(n_526),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_521),
.B(n_509),
.C(n_10),
.Y(n_526)
);

AO21x1_ASAP7_75t_L g527 ( 
.A1(n_525),
.A2(n_523),
.B(n_10),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_527),
.B(n_10),
.C(n_12),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_529),
.A2(n_528),
.B(n_10),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_13),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_0),
.Y(n_532)
);


endmodule