module fake_aes_8508_n_14 (n_1, n_2, n_0, n_14);
input n_1;
input n_2;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
HB1xp67_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
BUFx10_ASAP7_75t_L g5 ( .A(n_4), .Y(n_5) );
OAI21x1_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_6), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_7), .B(n_5), .Y(n_9) );
NAND3x2_ASAP7_75t_L g10 ( .A(n_8), .B(n_5), .C(n_6), .Y(n_10) );
OAI22xp5_ASAP7_75t_L g11 ( .A1(n_9), .A2(n_8), .B1(n_1), .B2(n_2), .Y(n_11) );
OAI211xp5_ASAP7_75t_SL g12 ( .A1(n_10), .A2(n_0), .B(n_2), .C(n_9), .Y(n_12) );
INVxp67_ASAP7_75t_SL g13 ( .A(n_11), .Y(n_13) );
AOI21xp33_ASAP7_75t_SL g14 ( .A1(n_13), .A2(n_2), .B(n_12), .Y(n_14) );
endmodule