module fake_jpeg_30569_n_15 (n_3, n_2, n_1, n_0, n_4, n_15);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_15;

wire n_13;
wire n_11;
wire n_14;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

NAND2xp5_ASAP7_75t_SL g5 ( 
.A(n_3),
.B(n_4),
.Y(n_5)
);

INVx11_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_2),
.Y(n_7)
);

AOI22xp33_ASAP7_75t_L g8 ( 
.A1(n_2),
.A2(n_3),
.B1(n_0),
.B2(n_1),
.Y(n_8)
);

OAI22xp5_ASAP7_75t_L g9 ( 
.A1(n_8),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_9)
);

AOI22xp5_ASAP7_75t_SL g12 ( 
.A1(n_9),
.A2(n_8),
.B1(n_5),
.B2(n_7),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_7),
.B(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_12),
.B(n_9),
.C(n_6),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_13),
.A2(n_11),
.B(n_6),
.Y(n_14)
);

BUFx24_ASAP7_75t_SL g15 ( 
.A(n_14),
.Y(n_15)
);


endmodule