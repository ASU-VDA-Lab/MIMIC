module fake_netlist_6_118_n_1775 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1775);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1775;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_87),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_18),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_183),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_69),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_23),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_171),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_67),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_51),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_8),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_9),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_160),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_96),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_12),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_164),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_137),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_84),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_85),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_7),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_55),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_141),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_117),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_39),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_147),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_154),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_30),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_177),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_45),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_122),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_39),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_149),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

BUFx8_ASAP7_75t_SL g222 ( 
.A(n_106),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_127),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_2),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_120),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_116),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_179),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_112),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_36),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_14),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_19),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_123),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_49),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_102),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_110),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_78),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_71),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_145),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_124),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_150),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_17),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_32),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_158),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_136),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_10),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_64),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_111),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_105),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_81),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_58),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_169),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_157),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_36),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_156),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_10),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_89),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_68),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_9),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_114),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_103),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_148),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_50),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_130),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_2),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_107),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_21),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_75),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_73),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_82),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_151),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_128),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_133),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_168),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_152),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_47),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_27),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_37),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_46),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_37),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_125),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_62),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_26),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_180),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_18),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_42),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_181),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_6),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_19),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_21),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_22),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_42),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_35),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_162),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_4),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_91),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_109),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_54),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_108),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_61),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_49),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_135),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_3),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_92),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_48),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_182),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_43),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_27),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_153),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_12),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_83),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_97),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_95),
.Y(n_313)
);

BUFx8_ASAP7_75t_SL g314 ( 
.A(n_52),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_54),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_45),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_101),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_129),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_48),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_161),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_121),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_46),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_52),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_77),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_6),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_74),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_33),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_134),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_23),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_44),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_8),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_57),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_172),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_98),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g335 ( 
.A(n_175),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_144),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_99),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_35),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_22),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_132),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_146),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_76),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_1),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_86),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_56),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_38),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_30),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_57),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_31),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_143),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_63),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_115),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_113),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_26),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_138),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_72),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_53),
.Y(n_357)
);

BUFx5_ASAP7_75t_L g358 ( 
.A(n_88),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_15),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_25),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_14),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_0),
.Y(n_362)
);

BUFx5_ASAP7_75t_L g363 ( 
.A(n_142),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_79),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_7),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_66),
.Y(n_366)
);

INVx4_ASAP7_75t_R g367 ( 
.A(n_5),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_173),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_34),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_286),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_301),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_222),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_314),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_273),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_229),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_286),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_220),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_249),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_223),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_286),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_286),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_275),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_227),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_286),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_L g385 ( 
.A(n_288),
.B(n_0),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_286),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_284),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_201),
.B(n_3),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_317),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_219),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_226),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_286),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_228),
.Y(n_393)
);

INVxp33_ASAP7_75t_L g394 ( 
.A(n_232),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_226),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_233),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_235),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_250),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_286),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_236),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_238),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_250),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_239),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_241),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_216),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_320),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_244),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_248),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_216),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_253),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_258),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_252),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_255),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_353),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_216),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_257),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_289),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_216),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_260),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_261),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_262),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_266),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_268),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_270),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_349),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_271),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_216),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_272),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_307),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_307),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_307),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_307),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_274),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_296),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_307),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_300),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_358),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_358),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_254),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_254),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_201),
.B(n_4),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_306),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_312),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_280),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_341),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_344),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_280),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_292),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_263),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_350),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_278),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_352),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_355),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_358),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_354),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_356),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_189),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_185),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_292),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_303),
.B(n_5),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_189),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_195),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_305),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_224),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_305),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_425),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_391),
.B(n_309),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_375),
.B(n_343),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_395),
.B(n_213),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_370),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_405),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_370),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_437),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_405),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_464),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_402),
.B(n_213),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_376),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_409),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_409),
.B(n_309),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_457),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_376),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_415),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_415),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_388),
.B(n_304),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_441),
.B(n_265),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_418),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_398),
.B(n_277),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_398),
.B(n_277),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_418),
.B(n_304),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_427),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_427),
.B(n_429),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_380),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_380),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_429),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_381),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_381),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_458),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_461),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_437),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_430),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_431),
.B(n_335),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_431),
.Y(n_502)
);

INVx6_ASAP7_75t_L g503 ( 
.A(n_384),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_432),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_435),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_384),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_435),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_386),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_386),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_392),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_392),
.B(n_335),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_399),
.Y(n_512)
);

OR2x6_ASAP7_75t_L g513 ( 
.A(n_385),
.B(n_303),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_438),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_462),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_399),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_438),
.B(n_185),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_439),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_454),
.Y(n_519)
);

OR2x6_ASAP7_75t_L g520 ( 
.A(n_460),
.B(n_194),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_390),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_374),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_454),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_439),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_377),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_440),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_440),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_444),
.B(n_194),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_444),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_371),
.B(n_197),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_447),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_447),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_448),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_448),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_465),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_394),
.B(n_379),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_459),
.Y(n_537)
);

CKINVDCx8_ASAP7_75t_R g538 ( 
.A(n_417),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_416),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_459),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_463),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_463),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_509),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_517),
.B(n_383),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_485),
.A2(n_362),
.B1(n_251),
.B2(n_256),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_519),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_512),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_536),
.B(n_393),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_468),
.Y(n_549)
);

AND2x6_ASAP7_75t_L g550 ( 
.A(n_511),
.B(n_197),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_536),
.B(n_396),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_519),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_512),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_470),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_538),
.B(n_372),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_521),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_519),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_521),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_472),
.Y(n_559)
);

INVx1_ASAP7_75t_SL g560 ( 
.A(n_468),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_485),
.A2(n_362),
.B1(n_279),
.B2(n_290),
.Y(n_561)
);

AO22x2_ASAP7_75t_L g562 ( 
.A1(n_484),
.A2(n_264),
.B1(n_302),
.B2(n_287),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_470),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_484),
.A2(n_293),
.B1(n_295),
.B2(n_186),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_472),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g566 ( 
.A(n_466),
.B(n_451),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_523),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_472),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_517),
.B(n_397),
.Y(n_569)
);

NAND2xp33_ASAP7_75t_SL g570 ( 
.A(n_469),
.B(n_348),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_477),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_539),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_475),
.B(n_400),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_477),
.Y(n_574)
);

INVx5_ASAP7_75t_L g575 ( 
.A(n_470),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_477),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_481),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_475),
.B(n_401),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_475),
.B(n_403),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_502),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_479),
.B(n_465),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_481),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_467),
.B(n_404),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_467),
.B(n_407),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_498),
.A2(n_424),
.B1(n_428),
.B2(n_453),
.Y(n_585)
);

AND2x6_ASAP7_75t_L g586 ( 
.A(n_511),
.B(n_264),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_487),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_522),
.B(n_408),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_470),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_502),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_481),
.Y(n_591)
);

NAND3xp33_ASAP7_75t_L g592 ( 
.A(n_498),
.B(n_413),
.C(n_412),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_487),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_467),
.B(n_420),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_479),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_492),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_492),
.Y(n_597)
);

INVx5_ASAP7_75t_L g598 ( 
.A(n_470),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_511),
.B(n_422),
.Y(n_599)
);

INVxp67_ASAP7_75t_SL g600 ( 
.A(n_470),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_492),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_511),
.B(n_423),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_511),
.B(n_426),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_L g604 ( 
.A1(n_469),
.A2(n_302),
.B(n_287),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_493),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_493),
.Y(n_606)
);

AND2x6_ASAP7_75t_L g607 ( 
.A(n_489),
.B(n_340),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_520),
.B(n_433),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_515),
.A2(n_421),
.B1(n_434),
.B2(n_452),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_468),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_487),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_470),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_466),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_503),
.Y(n_614)
);

NOR3xp33_ASAP7_75t_L g615 ( 
.A(n_515),
.B(n_455),
.C(n_417),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_520),
.A2(n_308),
.B1(n_310),
.B2(n_315),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_523),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_493),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_495),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_479),
.Y(n_620)
);

INVx5_ASAP7_75t_L g621 ( 
.A(n_495),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_523),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_488),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_495),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_497),
.Y(n_625)
);

INVx1_ASAP7_75t_SL g626 ( 
.A(n_497),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_530),
.A2(n_445),
.B1(n_419),
.B2(n_450),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_495),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_488),
.Y(n_629)
);

BUFx10_ASAP7_75t_L g630 ( 
.A(n_539),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_488),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_523),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_497),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_495),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_506),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_506),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_508),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_508),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_508),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_523),
.Y(n_640)
);

AO21x2_ASAP7_75t_L g641 ( 
.A1(n_476),
.A2(n_193),
.B(n_188),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_495),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_510),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_495),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_520),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_479),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_520),
.B(n_442),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_510),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_520),
.B(n_443),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_503),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_522),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_503),
.Y(n_652)
);

OR2x2_ASAP7_75t_SL g653 ( 
.A(n_480),
.B(n_455),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_510),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_471),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_522),
.B(n_456),
.Y(n_656)
);

AND2x6_ASAP7_75t_L g657 ( 
.A(n_489),
.B(n_340),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_471),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_525),
.B(n_436),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_496),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_474),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_474),
.Y(n_662)
);

NAND3xp33_ASAP7_75t_L g663 ( 
.A(n_476),
.B(n_449),
.C(n_231),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_496),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_478),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_496),
.Y(n_666)
);

NOR2x1p5_ASAP7_75t_L g667 ( 
.A(n_525),
.B(n_373),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_496),
.Y(n_668)
);

INVx4_ASAP7_75t_L g669 ( 
.A(n_496),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_520),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_479),
.B(n_489),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_478),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_501),
.B(n_528),
.Y(n_673)
);

INVx1_ASAP7_75t_SL g674 ( 
.A(n_480),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_525),
.B(n_446),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_482),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_538),
.B(n_410),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_538),
.B(n_411),
.Y(n_678)
);

OR2x6_ASAP7_75t_L g679 ( 
.A(n_530),
.B(n_322),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_513),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_483),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_483),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_501),
.B(n_414),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_501),
.B(n_192),
.Y(n_684)
);

INVx5_ASAP7_75t_L g685 ( 
.A(n_496),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_496),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_530),
.A2(n_406),
.B1(n_389),
.B2(n_387),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_SL g688 ( 
.A(n_528),
.B(n_369),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_516),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_530),
.B(n_382),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_558),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_567),
.B(n_516),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_546),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_567),
.B(n_516),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_558),
.Y(n_695)
);

NOR3xp33_ASAP7_75t_L g696 ( 
.A(n_556),
.B(n_294),
.C(n_237),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_583),
.B(n_530),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_673),
.B(n_516),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_566),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_567),
.B(n_516),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_581),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_673),
.B(n_516),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_546),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_613),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_587),
.A2(n_530),
.B1(n_378),
.B2(n_513),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_673),
.B(n_516),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_566),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_581),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_674),
.B(n_513),
.Y(n_709)
);

BUFx4_ASAP7_75t_L g710 ( 
.A(n_572),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_552),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_604),
.A2(n_325),
.B1(n_330),
.B2(n_345),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_617),
.B(n_503),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_645),
.B(n_358),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_581),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_587),
.B(n_593),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_613),
.Y(n_717)
);

BUFx6f_ASAP7_75t_SL g718 ( 
.A(n_572),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_593),
.B(n_513),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_595),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_617),
.B(n_622),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_622),
.B(n_632),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_622),
.B(n_513),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_632),
.B(n_513),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_584),
.B(n_313),
.Y(n_725)
);

BUFx10_ASAP7_75t_L g726 ( 
.A(n_667),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_640),
.B(n_473),
.Y(n_727)
);

OR2x6_ASAP7_75t_L g728 ( 
.A(n_679),
.B(n_346),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_640),
.B(n_473),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_572),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_645),
.B(n_358),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_595),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_557),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_670),
.B(n_358),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_594),
.B(n_364),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_620),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_544),
.B(n_473),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_569),
.B(n_499),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_543),
.B(n_499),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_543),
.B(n_499),
.Y(n_740)
);

BUFx6f_ASAP7_75t_SL g741 ( 
.A(n_630),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_620),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_688),
.B(n_195),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_670),
.B(n_358),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_547),
.B(n_553),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_646),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_568),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_671),
.B(n_358),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_646),
.B(n_363),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_611),
.B(n_499),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_611),
.A2(n_629),
.B1(n_631),
.B2(n_623),
.Y(n_751)
);

OAI22x1_ASAP7_75t_R g752 ( 
.A1(n_549),
.A2(n_214),
.B1(n_211),
.B2(n_208),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_623),
.B(n_187),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_580),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_631),
.B(n_528),
.Y(n_755)
);

NAND3xp33_ASAP7_75t_L g756 ( 
.A(n_688),
.B(n_234),
.C(n_230),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_683),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_599),
.B(n_363),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_602),
.B(n_363),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_590),
.B(n_514),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_548),
.B(n_187),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_603),
.A2(n_336),
.B1(n_210),
.B2(n_209),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_662),
.Y(n_763)
);

NOR3xp33_ASAP7_75t_L g764 ( 
.A(n_585),
.B(n_243),
.C(n_242),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_608),
.B(n_363),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_684),
.B(n_514),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_662),
.B(n_514),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_L g768 ( 
.A1(n_679),
.A2(n_347),
.B1(n_359),
.B2(n_365),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_676),
.B(n_486),
.Y(n_769)
);

INVx8_ASAP7_75t_L g770 ( 
.A(n_679),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_676),
.B(n_486),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_681),
.B(n_682),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_568),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_681),
.B(n_490),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_682),
.B(n_490),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_655),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_550),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_655),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_647),
.B(n_363),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_570),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_651),
.B(n_263),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_658),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_625),
.B(n_196),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_649),
.B(n_363),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_600),
.B(n_494),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_680),
.A2(n_366),
.B1(n_297),
.B2(n_282),
.Y(n_786)
);

AOI22x1_ASAP7_75t_L g787 ( 
.A1(n_562),
.A2(n_366),
.B1(n_324),
.B2(n_218),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_571),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_551),
.B(n_190),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_658),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_571),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_592),
.B(n_190),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_562),
.A2(n_240),
.B1(n_212),
.B2(n_217),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_626),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_661),
.Y(n_795)
);

OR2x6_ASAP7_75t_L g796 ( 
.A(n_679),
.B(n_198),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_663),
.B(n_573),
.Y(n_797)
);

INVx8_ASAP7_75t_L g798 ( 
.A(n_607),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_661),
.Y(n_799)
);

INVx8_ASAP7_75t_L g800 ( 
.A(n_657),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_570),
.A2(n_337),
.B1(n_203),
.B2(n_204),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_657),
.B(n_500),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_665),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_657),
.B(n_500),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_657),
.B(n_641),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_574),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_680),
.B(n_205),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_545),
.A2(n_518),
.B(n_533),
.C(n_532),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_609),
.B(n_263),
.Y(n_809)
);

OR2x6_ASAP7_75t_L g810 ( 
.A(n_677),
.B(n_206),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_574),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_616),
.B(n_221),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_665),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_627),
.B(n_246),
.C(n_276),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_641),
.B(n_504),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_562),
.A2(n_245),
.B1(n_225),
.B2(n_247),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_672),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_641),
.B(n_504),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_550),
.A2(n_215),
.B1(n_200),
.B2(n_203),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_672),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_678),
.B(n_269),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_550),
.A2(n_586),
.B1(n_615),
.B2(n_578),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_579),
.B(n_200),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_633),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_560),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_642),
.B(n_505),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_562),
.A2(n_281),
.B1(n_299),
.B2(n_311),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_576),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_559),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_614),
.B(n_321),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_644),
.B(n_505),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_660),
.B(n_507),
.Y(n_832)
);

INVxp33_ASAP7_75t_L g833 ( 
.A(n_687),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_559),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_650),
.B(n_333),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_565),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_550),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_588),
.B(n_204),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_565),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_577),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_597),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_660),
.B(n_507),
.Y(n_842)
);

AND2x2_ASAP7_75t_SL g843 ( 
.A(n_561),
.B(n_564),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_721),
.A2(n_722),
.B(n_694),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_725),
.B(n_555),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_805),
.A2(n_601),
.B(n_597),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_695),
.B(n_690),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_691),
.B(n_659),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_704),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_699),
.B(n_675),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_692),
.A2(n_612),
.B(n_563),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_707),
.B(n_630),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_SL g853 ( 
.A1(n_714),
.A2(n_744),
.B(n_731),
.C(n_765),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_803),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_755),
.B(n_601),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_725),
.A2(n_652),
.B(n_342),
.C(n_351),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_772),
.B(n_636),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_803),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_735),
.B(n_824),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_748),
.A2(n_638),
.B(n_636),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_735),
.B(n_630),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_700),
.A2(n_612),
.B(n_563),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_794),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_713),
.A2(n_619),
.B(n_612),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_716),
.B(n_550),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_780),
.A2(n_808),
.B(n_807),
.C(n_765),
.Y(n_866)
);

OAI21xp33_ASAP7_75t_L g867 ( 
.A1(n_823),
.A2(n_838),
.B(n_789),
.Y(n_867)
);

OR2x2_ASAP7_75t_SL g868 ( 
.A(n_743),
.B(n_756),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_778),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_778),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_704),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_697),
.A2(n_586),
.B1(n_550),
.B2(n_656),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_776),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_697),
.B(n_586),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_732),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_717),
.B(n_653),
.Y(n_876)
);

O2A1O1Ixp5_ASAP7_75t_L g877 ( 
.A1(n_779),
.A2(n_689),
.B(n_686),
.C(n_664),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_763),
.B(n_586),
.Y(n_878)
);

NOR2xp67_ASAP7_75t_L g879 ( 
.A(n_825),
.B(n_638),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_727),
.A2(n_624),
.B(n_619),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_729),
.A2(n_624),
.B(n_619),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_753),
.B(n_586),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_833),
.B(n_653),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_766),
.A2(n_724),
.B(n_723),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_709),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_781),
.B(n_518),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_737),
.A2(n_634),
.B(n_624),
.Y(n_887)
);

BUFx8_ASAP7_75t_L g888 ( 
.A(n_718),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_753),
.B(n_586),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_833),
.B(n_549),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_782),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_790),
.Y(n_892)
);

AOI21xp33_ASAP7_75t_L g893 ( 
.A1(n_843),
.A2(n_643),
.B(n_639),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_745),
.B(n_738),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_757),
.B(n_610),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_797),
.A2(n_689),
.B1(n_686),
.B2(n_664),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_795),
.Y(n_897)
);

O2A1O1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_807),
.A2(n_648),
.B(n_654),
.C(n_635),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_698),
.A2(n_669),
.B(n_634),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_698),
.A2(n_669),
.B(n_634),
.Y(n_900)
);

INVx5_ASAP7_75t_L g901 ( 
.A(n_798),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_799),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_761),
.B(n_610),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_719),
.B(n_664),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_726),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_730),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_797),
.B(n_209),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_702),
.A2(n_669),
.B(n_628),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_754),
.B(n_666),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_R g910 ( 
.A(n_718),
.B(n_210),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_751),
.B(n_666),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_823),
.B(n_524),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_761),
.A2(n_689),
.B(n_686),
.C(n_637),
.Y(n_913)
);

AO22x1_ASAP7_75t_L g914 ( 
.A1(n_814),
.A2(n_319),
.B1(n_316),
.B2(n_323),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_720),
.A2(n_606),
.B1(n_582),
.B2(n_637),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_702),
.A2(n_706),
.B(n_750),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_789),
.B(n_215),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_701),
.B(n_591),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_734),
.A2(n_628),
.B(n_668),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_813),
.B(n_591),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_792),
.A2(n_606),
.B(n_596),
.C(n_635),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_705),
.B(n_792),
.Y(n_922)
);

CKINVDCx6p67_ASAP7_75t_R g923 ( 
.A(n_741),
.Y(n_923)
);

INVx4_ASAP7_75t_L g924 ( 
.A(n_732),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_708),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_817),
.B(n_605),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_820),
.B(n_769),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_771),
.B(n_618),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_774),
.B(n_554),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_822),
.B(n_318),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_802),
.A2(n_628),
.B(n_589),
.Y(n_931)
);

OAI21xp33_ASAP7_75t_L g932 ( 
.A1(n_712),
.A2(n_696),
.B(n_764),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_804),
.A2(n_589),
.B(n_554),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_715),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_693),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_783),
.B(n_318),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_815),
.A2(n_621),
.B(n_598),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_712),
.A2(n_337),
.B(n_328),
.C(n_326),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_809),
.B(n_326),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_775),
.B(n_534),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_703),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_810),
.B(n_524),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_798),
.A2(n_685),
.B(n_621),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_736),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_726),
.Y(n_945)
);

AND2x2_ASAP7_75t_SL g946 ( 
.A(n_801),
.B(n_367),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_818),
.A2(n_598),
.B(n_575),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_742),
.A2(n_746),
.B(n_759),
.C(n_758),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_810),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_728),
.B(n_526),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_762),
.B(n_334),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_798),
.A2(n_685),
.B(n_598),
.Y(n_952)
);

AND2x6_ASAP7_75t_L g953 ( 
.A(n_777),
.B(n_526),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_800),
.A2(n_685),
.B(n_598),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_829),
.B(n_534),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_834),
.B(n_534),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_836),
.B(n_534),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_839),
.B(n_534),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_841),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_800),
.A2(n_685),
.B(n_575),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_800),
.A2(n_685),
.B(n_575),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_785),
.A2(n_744),
.B(n_731),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_758),
.B(n_534),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_747),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_773),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_810),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_821),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_760),
.A2(n_575),
.B(n_491),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_759),
.B(n_534),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_821),
.B(n_334),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_821),
.B(n_527),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_784),
.A2(n_542),
.B(n_541),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_749),
.A2(n_542),
.B(n_540),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_749),
.A2(n_532),
.B(n_527),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_710),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_739),
.A2(n_533),
.B(n_531),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_812),
.A2(n_535),
.B1(n_191),
.B2(n_336),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_788),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_791),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_740),
.A2(n_368),
.B(n_531),
.C(n_529),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_777),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_819),
.A2(n_368),
.B1(n_535),
.B2(n_537),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_812),
.A2(n_535),
.B1(n_191),
.B2(n_360),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_826),
.A2(n_842),
.B(n_831),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_767),
.A2(n_832),
.B(n_806),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_837),
.A2(n_535),
.B(n_361),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_786),
.A2(n_191),
.B(n_211),
.C(n_208),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_837),
.A2(n_535),
.B(n_357),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_811),
.B(n_535),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_711),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_793),
.A2(n_827),
.B1(n_816),
.B2(n_770),
.Y(n_991)
);

AO21x1_ASAP7_75t_L g992 ( 
.A1(n_768),
.A2(n_11),
.B(n_13),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_770),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_828),
.B(n_840),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_733),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_830),
.Y(n_996)
);

OAI21xp33_ASAP7_75t_L g997 ( 
.A1(n_793),
.A2(n_339),
.B(n_338),
.Y(n_997)
);

INVx5_ASAP7_75t_L g998 ( 
.A(n_770),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_816),
.A2(n_291),
.B(n_259),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_835),
.A2(n_830),
.B(n_796),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_796),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_827),
.B(n_768),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_728),
.B(n_196),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_835),
.B(n_199),
.Y(n_1004)
);

OAI321xp33_ASAP7_75t_L g1005 ( 
.A1(n_796),
.A2(n_339),
.A3(n_338),
.B1(n_332),
.B2(n_331),
.C(n_329),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_787),
.A2(n_298),
.B(n_267),
.C(n_283),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_728),
.B(n_332),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_752),
.A2(n_285),
.B(n_329),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_741),
.B(n_331),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_725),
.A2(n_327),
.B(n_323),
.C(n_319),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_884),
.A2(n_70),
.B(n_184),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_867),
.B(n_327),
.Y(n_1012)
);

INVx4_ASAP7_75t_L g1013 ( 
.A(n_998),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_859),
.B(n_316),
.Y(n_1014)
);

AOI222xp33_ASAP7_75t_L g1015 ( 
.A1(n_903),
.A2(n_214),
.B1(n_207),
.B2(n_202),
.C1(n_199),
.C2(n_20),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_849),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_917),
.A2(n_207),
.B1(n_202),
.B2(n_178),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_959),
.Y(n_1018)
);

OA21x2_ASAP7_75t_L g1019 ( 
.A1(n_846),
.A2(n_166),
.B(n_163),
.Y(n_1019)
);

INVx4_ASAP7_75t_L g1020 ( 
.A(n_998),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_894),
.A2(n_159),
.B(n_140),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_R g1022 ( 
.A(n_906),
.B(n_139),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_922),
.A2(n_11),
.B(n_13),
.C(n_16),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_981),
.Y(n_1024)
);

INVxp33_ASAP7_75t_SL g1025 ( 
.A(n_890),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_874),
.A2(n_889),
.B(n_882),
.Y(n_1026)
);

BUFx4f_ASAP7_75t_L g1027 ( 
.A(n_923),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_888),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_888),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_845),
.A2(n_16),
.B(n_17),
.C(n_20),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_912),
.B(n_24),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_993),
.Y(n_1032)
);

CKINVDCx6p67_ASAP7_75t_R g1033 ( 
.A(n_905),
.Y(n_1033)
);

BUFx10_ASAP7_75t_L g1034 ( 
.A(n_883),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_854),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_865),
.A2(n_119),
.B(n_118),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_855),
.B(n_104),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_844),
.A2(n_100),
.B(n_94),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_886),
.B(n_24),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_993),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_932),
.A2(n_93),
.B1(n_90),
.B2(n_80),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_927),
.B(n_25),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_962),
.A2(n_65),
.B(n_28),
.Y(n_1043)
);

OAI21xp33_ASAP7_75t_L g1044 ( 
.A1(n_939),
.A2(n_28),
.B(n_29),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_871),
.B(n_847),
.Y(n_1045)
);

BUFx12f_ASAP7_75t_L g1046 ( 
.A(n_945),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_936),
.B(n_29),
.Y(n_1047)
);

INVx5_ASAP7_75t_L g1048 ( 
.A(n_981),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_853),
.A2(n_929),
.B(n_887),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_929),
.A2(n_60),
.B(n_32),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_981),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_855),
.B(n_31),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_863),
.Y(n_1053)
);

OAI21xp33_ASAP7_75t_L g1054 ( 
.A1(n_970),
.A2(n_33),
.B(n_34),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_875),
.B(n_38),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_910),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_991),
.B(n_40),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_857),
.A2(n_40),
.B(n_41),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_857),
.A2(n_60),
.B(n_43),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_848),
.B(n_41),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_850),
.Y(n_1061)
);

NAND2x1p5_ASAP7_75t_L g1062 ( 
.A(n_998),
.B(n_47),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_875),
.B(n_51),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_984),
.A2(n_53),
.B(n_55),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_916),
.A2(n_58),
.B(n_59),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_861),
.A2(n_59),
.B1(n_885),
.B2(n_895),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_R g1067 ( 
.A(n_998),
.B(n_993),
.Y(n_1067)
);

INVxp67_ASAP7_75t_L g1068 ( 
.A(n_852),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_879),
.B(n_946),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_949),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_876),
.B(n_907),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_899),
.A2(n_900),
.B(n_862),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_858),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_851),
.A2(n_933),
.B(n_931),
.Y(n_1074)
);

XOR2x2_ASAP7_75t_SL g1075 ( 
.A(n_1002),
.B(n_1007),
.Y(n_1075)
);

OAI22x1_ASAP7_75t_L g1076 ( 
.A1(n_966),
.A2(n_967),
.B1(n_1002),
.B2(n_1001),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_868),
.A2(n_872),
.B1(n_1010),
.B2(n_938),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_934),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_1003),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_924),
.B(n_950),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_950),
.Y(n_1081)
);

AO32x1_ASAP7_75t_L g1082 ( 
.A1(n_891),
.A2(n_902),
.A3(n_897),
.B1(n_892),
.B2(n_873),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_965),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_1001),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_866),
.A2(n_996),
.B(n_1000),
.C(n_999),
.Y(n_1085)
);

BUFx4f_ASAP7_75t_SL g1086 ( 
.A(n_975),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_948),
.A2(n_987),
.B(n_925),
.C(n_893),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_928),
.A2(n_901),
.B1(n_925),
.B2(n_977),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_920),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_924),
.B(n_971),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_893),
.A2(n_980),
.B(n_942),
.C(n_930),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_1005),
.A2(n_951),
.B(n_1008),
.C(n_1007),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_997),
.B(n_1009),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_937),
.A2(n_947),
.B(n_864),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_944),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_901),
.A2(n_911),
.B1(n_1004),
.B2(n_896),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_856),
.A2(n_1004),
.B(n_1006),
.C(n_992),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_920),
.Y(n_1098)
);

AOI21x1_ASAP7_75t_L g1099 ( 
.A1(n_940),
.A2(n_957),
.B(n_956),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_870),
.A2(n_990),
.B1(n_941),
.B2(n_935),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_965),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_877),
.A2(n_913),
.B(n_921),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_914),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_953),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_964),
.B(n_995),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_869),
.B(n_978),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_979),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_974),
.B(n_983),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_878),
.A2(n_880),
.B(n_881),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_926),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_940),
.A2(n_904),
.B(n_908),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_901),
.B(n_976),
.Y(n_1112)
);

INVx5_ASAP7_75t_L g1113 ( 
.A(n_953),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_919),
.A2(n_901),
.B(n_985),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_994),
.B(n_918),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_909),
.B(n_994),
.Y(n_1116)
);

INVx6_ASAP7_75t_L g1117 ( 
.A(n_953),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_898),
.A2(n_988),
.B(n_986),
.C(n_860),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_989),
.Y(n_1119)
);

OAI21xp33_ASAP7_75t_L g1120 ( 
.A1(n_982),
.A2(n_958),
.B(n_956),
.Y(n_1120)
);

AOI21x1_ASAP7_75t_L g1121 ( 
.A1(n_955),
.A2(n_958),
.B(n_957),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_915),
.A2(n_955),
.B1(n_969),
.B2(n_963),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_953),
.B(n_989),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_953),
.Y(n_1124)
);

BUFx12f_ASAP7_75t_L g1125 ( 
.A(n_973),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_972),
.B(n_968),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_943),
.A2(n_952),
.B1(n_954),
.B2(n_960),
.Y(n_1127)
);

OAI21xp33_ASAP7_75t_L g1128 ( 
.A1(n_961),
.A2(n_556),
.B(n_939),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_849),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_859),
.B(n_558),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_894),
.B(n_855),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_858),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_894),
.B(n_855),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_871),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_894),
.B(n_855),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_859),
.B(n_556),
.Y(n_1136)
);

NAND2xp33_ASAP7_75t_R g1137 ( 
.A(n_890),
.B(n_539),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_894),
.B(n_855),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_894),
.B(n_855),
.Y(n_1139)
);

BUFx8_ASAP7_75t_L g1140 ( 
.A(n_949),
.Y(n_1140)
);

BUFx12f_ASAP7_75t_SL g1141 ( 
.A(n_852),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_894),
.B(n_855),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_894),
.B(n_855),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_859),
.B(n_556),
.Y(n_1144)
);

NAND2x1p5_ASAP7_75t_L g1145 ( 
.A(n_998),
.B(n_901),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_993),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_867),
.A2(n_917),
.B(n_922),
.C(n_845),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_849),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_884),
.A2(n_722),
.B(n_721),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_959),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_867),
.A2(n_1002),
.B1(n_991),
.B2(n_843),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_849),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_858),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_884),
.A2(n_722),
.B(n_721),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_R g1155 ( 
.A(n_906),
.B(n_539),
.Y(n_1155)
);

INVx1_ASAP7_75t_SL g1156 ( 
.A(n_849),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_849),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1094),
.A2(n_1085),
.A3(n_1151),
.B(n_1049),
.Y(n_1158)
);

AND2x6_ASAP7_75t_L g1159 ( 
.A(n_1124),
.B(n_1123),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1136),
.B(n_1144),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1131),
.B(n_1133),
.Y(n_1161)
);

NAND3xp33_ASAP7_75t_L g1162 ( 
.A(n_1047),
.B(n_1147),
.C(n_1015),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_1129),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1092),
.A2(n_1151),
.B(n_1015),
.C(n_1044),
.Y(n_1164)
);

OAI22x1_ASAP7_75t_L g1165 ( 
.A1(n_1066),
.A2(n_1071),
.B1(n_1069),
.B2(n_1103),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1150),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_SL g1167 ( 
.A1(n_1131),
.A2(n_1135),
.B(n_1133),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_SL g1168 ( 
.A1(n_1025),
.A2(n_1057),
.B1(n_1093),
.B2(n_1079),
.Y(n_1168)
);

AO32x2_ASAP7_75t_L g1169 ( 
.A1(n_1077),
.A2(n_1096),
.A3(n_1122),
.B1(n_1088),
.B2(n_1075),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_1130),
.B(n_1014),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1078),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_L g1172 ( 
.A(n_1017),
.B(n_1054),
.C(n_1064),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1156),
.B(n_1157),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1135),
.B(n_1138),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1077),
.A2(n_1061),
.B1(n_1060),
.B2(n_1108),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1114),
.A2(n_1026),
.B(n_1154),
.Y(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1012),
.A2(n_1031),
.B(n_1023),
.C(n_1039),
.Y(n_1177)
);

AOI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1112),
.A2(n_1121),
.B(n_1099),
.Y(n_1178)
);

INVxp67_ASAP7_75t_L g1179 ( 
.A(n_1016),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_1030),
.B(n_1128),
.C(n_1091),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1084),
.B(n_1080),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1035),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1045),
.B(n_1068),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1138),
.B(n_1139),
.Y(n_1184)
);

BUFx8_ASAP7_75t_L g1185 ( 
.A(n_1046),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_1134),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1139),
.B(n_1142),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_SL g1188 ( 
.A1(n_1142),
.A2(n_1143),
.B(n_1087),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1081),
.B(n_1034),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1097),
.A2(n_1143),
.B(n_1043),
.C(n_1065),
.Y(n_1190)
);

INVxp67_ASAP7_75t_SL g1191 ( 
.A(n_1148),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1115),
.B(n_1089),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1116),
.A2(n_1042),
.B(n_1041),
.C(n_1120),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1149),
.A2(n_1127),
.B(n_1111),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1013),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1098),
.B(n_1110),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1105),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1152),
.B(n_1141),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1096),
.A2(n_1037),
.B(n_1052),
.C(n_1059),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1073),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1053),
.B(n_1034),
.Y(n_1201)
);

OA21x2_ASAP7_75t_L g1202 ( 
.A1(n_1102),
.A2(n_1126),
.B(n_1118),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_SL g1203 ( 
.A1(n_1088),
.A2(n_1145),
.B(n_1127),
.Y(n_1203)
);

NAND3xp33_ASAP7_75t_L g1204 ( 
.A(n_1137),
.B(n_1058),
.C(n_1050),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1055),
.A2(n_1063),
.B(n_1090),
.C(n_1107),
.Y(n_1205)
);

OAI22x1_ASAP7_75t_L g1206 ( 
.A1(n_1062),
.A2(n_1070),
.B1(n_1104),
.B2(n_1095),
.Y(n_1206)
);

BUFx16f_ASAP7_75t_R g1207 ( 
.A(n_1140),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1083),
.B(n_1101),
.Y(n_1208)
);

AOI221x1_ASAP7_75t_L g1209 ( 
.A1(n_1076),
.A2(n_1011),
.B1(n_1038),
.B2(n_1036),
.C(n_1021),
.Y(n_1209)
);

OAI22x1_ASAP7_75t_L g1210 ( 
.A1(n_1062),
.A2(n_1106),
.B1(n_1019),
.B2(n_1056),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_1119),
.A2(n_1082),
.A3(n_1132),
.B(n_1153),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1100),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1024),
.B(n_1051),
.Y(n_1213)
);

AOI221xp5_ASAP7_75t_SL g1214 ( 
.A1(n_1051),
.A2(n_1146),
.B1(n_1040),
.B2(n_1032),
.C(n_1082),
.Y(n_1214)
);

AO31x2_ASAP7_75t_L g1215 ( 
.A1(n_1082),
.A2(n_1013),
.A3(n_1020),
.B(n_1125),
.Y(n_1215)
);

BUFx2_ASAP7_75t_SL g1216 ( 
.A(n_1032),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1113),
.A2(n_1048),
.B(n_1020),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1113),
.A2(n_1117),
.A3(n_1048),
.B(n_1067),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1117),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1027),
.A2(n_1040),
.B(n_1032),
.C(n_1146),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_1117),
.A2(n_1040),
.A3(n_1140),
.B(n_1022),
.Y(n_1221)
);

NAND3xp33_ASAP7_75t_L g1222 ( 
.A(n_1028),
.B(n_1029),
.C(n_1155),
.Y(n_1222)
);

INVxp67_ASAP7_75t_L g1223 ( 
.A(n_1027),
.Y(n_1223)
);

AOI211x1_ASAP7_75t_L g1224 ( 
.A1(n_1033),
.A2(n_1151),
.B(n_867),
.C(n_992),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1086),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1046),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1130),
.B(n_558),
.Y(n_1227)
);

BUFx10_ASAP7_75t_L g1228 ( 
.A(n_1136),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1018),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1094),
.A2(n_1085),
.A3(n_1151),
.B(n_1049),
.Y(n_1230)
);

OA21x2_ASAP7_75t_L g1231 ( 
.A1(n_1102),
.A2(n_1094),
.B(n_1026),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1131),
.B(n_1133),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1047),
.A2(n_867),
.B(n_845),
.C(n_917),
.Y(n_1233)
);

O2A1O1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1047),
.A2(n_867),
.B(n_845),
.C(n_917),
.Y(n_1234)
);

AOI221x1_ASAP7_75t_L g1235 ( 
.A1(n_1047),
.A2(n_867),
.B1(n_1151),
.B2(n_1044),
.C(n_1077),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1155),
.Y(n_1236)
);

NAND2xp33_ASAP7_75t_L g1237 ( 
.A(n_1067),
.B(n_867),
.Y(n_1237)
);

BUFx2_ASAP7_75t_SL g1238 ( 
.A(n_1134),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1109),
.A2(n_1072),
.B(n_1074),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1109),
.A2(n_1072),
.B(n_1074),
.Y(n_1240)
);

AOI211x1_ASAP7_75t_L g1241 ( 
.A1(n_1151),
.A2(n_867),
.B(n_992),
.C(n_1057),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1131),
.B(n_1133),
.Y(n_1242)
);

AOI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1112),
.A2(n_1114),
.B(n_1121),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1109),
.A2(n_1072),
.B(n_1074),
.Y(n_1244)
);

AO21x2_ASAP7_75t_L g1245 ( 
.A1(n_1094),
.A2(n_1102),
.B(n_1049),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1109),
.A2(n_1072),
.B(n_1074),
.Y(n_1246)
);

NAND3xp33_ASAP7_75t_SL g1247 ( 
.A(n_1015),
.B(n_867),
.C(n_521),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1013),
.Y(n_1248)
);

INVx5_ASAP7_75t_L g1249 ( 
.A(n_1117),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1151),
.A2(n_1133),
.B1(n_1135),
.B2(n_1131),
.Y(n_1250)
);

NOR4xp25_ASAP7_75t_L g1251 ( 
.A(n_1054),
.B(n_867),
.C(n_1147),
.D(n_1044),
.Y(n_1251)
);

OR2x6_ASAP7_75t_L g1252 ( 
.A(n_1070),
.B(n_993),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1109),
.A2(n_1072),
.B(n_1074),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1129),
.Y(n_1254)
);

AOI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1047),
.A2(n_867),
.B1(n_1151),
.B2(n_917),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1131),
.B(n_1133),
.Y(n_1256)
);

AOI221x1_ASAP7_75t_L g1257 ( 
.A1(n_1047),
.A2(n_867),
.B1(n_1151),
.B2(n_1044),
.C(n_1077),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1085),
.A2(n_1151),
.B(n_1026),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_1094),
.A2(n_1085),
.A3(n_1151),
.B(n_1049),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1032),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_SL g1261 ( 
.A1(n_1085),
.A2(n_991),
.B(n_1131),
.Y(n_1261)
);

INVx1_ASAP7_75t_SL g1262 ( 
.A(n_1156),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1131),
.B(n_1133),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1134),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1085),
.A2(n_1151),
.B(n_1026),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1147),
.A2(n_867),
.B(n_1047),
.C(n_917),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1018),
.Y(n_1267)
);

AO22x2_ASAP7_75t_L g1268 ( 
.A1(n_1151),
.A2(n_1077),
.B1(n_922),
.B2(n_1057),
.Y(n_1268)
);

BUFx10_ASAP7_75t_L g1269 ( 
.A(n_1136),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1018),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1109),
.A2(n_1072),
.B(n_1074),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1013),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1109),
.A2(n_1072),
.B(n_1074),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1136),
.B(n_1144),
.Y(n_1274)
);

AO31x2_ASAP7_75t_L g1275 ( 
.A1(n_1094),
.A2(n_1085),
.A3(n_1151),
.B(n_1049),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1018),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1130),
.B(n_558),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1131),
.B(n_1133),
.Y(n_1278)
);

O2A1O1Ixp33_ASAP7_75t_SL g1279 ( 
.A1(n_1085),
.A2(n_1057),
.B(n_1151),
.C(n_867),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1130),
.B(n_558),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1129),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1109),
.A2(n_1072),
.B(n_1074),
.Y(n_1282)
);

AO21x1_ASAP7_75t_L g1283 ( 
.A1(n_1151),
.A2(n_1147),
.B(n_1077),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1085),
.A2(n_1151),
.B(n_1026),
.Y(n_1284)
);

AO31x2_ASAP7_75t_L g1285 ( 
.A1(n_1094),
.A2(n_1085),
.A3(n_1151),
.B(n_1049),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_SL g1286 ( 
.A1(n_1097),
.A2(n_866),
.B(n_1043),
.Y(n_1286)
);

INVx6_ASAP7_75t_L g1287 ( 
.A(n_1249),
.Y(n_1287)
);

INVx6_ASAP7_75t_L g1288 ( 
.A(n_1249),
.Y(n_1288)
);

CKINVDCx11_ASAP7_75t_R g1289 ( 
.A(n_1207),
.Y(n_1289)
);

NOR2x1_ASAP7_75t_L g1290 ( 
.A(n_1167),
.B(n_1222),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1249),
.B(n_1195),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1236),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1162),
.A2(n_1247),
.B1(n_1160),
.B2(n_1274),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1162),
.A2(n_1255),
.B1(n_1172),
.B2(n_1168),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1255),
.A2(n_1172),
.B1(n_1168),
.B2(n_1283),
.Y(n_1295)
);

BUFx12f_ASAP7_75t_L g1296 ( 
.A(n_1185),
.Y(n_1296)
);

OAI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1235),
.A2(n_1257),
.B1(n_1165),
.B2(n_1170),
.Y(n_1297)
);

BUFx12f_ASAP7_75t_L g1298 ( 
.A(n_1185),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1226),
.Y(n_1299)
);

BUFx12f_ASAP7_75t_L g1300 ( 
.A(n_1281),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_SL g1301 ( 
.A1(n_1164),
.A2(n_1234),
.B(n_1233),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1173),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1174),
.B(n_1256),
.Y(n_1303)
);

INVx8_ASAP7_75t_L g1304 ( 
.A(n_1252),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1268),
.A2(n_1228),
.B1(n_1269),
.B2(n_1180),
.Y(n_1305)
);

BUFx12f_ASAP7_75t_L g1306 ( 
.A(n_1264),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1229),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1268),
.A2(n_1204),
.B1(n_1180),
.B2(n_1175),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1174),
.B(n_1256),
.Y(n_1309)
);

BUFx12f_ASAP7_75t_L g1310 ( 
.A(n_1252),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1161),
.B(n_1184),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1204),
.A2(n_1280),
.B1(n_1237),
.B2(n_1269),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1218),
.Y(n_1313)
);

BUFx10_ASAP7_75t_L g1314 ( 
.A(n_1201),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_SL g1315 ( 
.A1(n_1228),
.A2(n_1284),
.B1(n_1265),
.B2(n_1258),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1266),
.A2(n_1183),
.B1(n_1198),
.B2(n_1189),
.Y(n_1316)
);

CKINVDCx11_ASAP7_75t_R g1317 ( 
.A(n_1207),
.Y(n_1317)
);

CKINVDCx11_ASAP7_75t_R g1318 ( 
.A(n_1262),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1171),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1225),
.Y(n_1320)
);

CKINVDCx11_ASAP7_75t_R g1321 ( 
.A(n_1262),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1250),
.A2(n_1284),
.B1(n_1265),
.B2(n_1258),
.Y(n_1322)
);

OAI22x1_ASAP7_75t_L g1323 ( 
.A1(n_1191),
.A2(n_1181),
.B1(n_1182),
.B2(n_1270),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1187),
.B(n_1232),
.Y(n_1324)
);

BUFx4f_ASAP7_75t_SL g1325 ( 
.A(n_1225),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1238),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1163),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1242),
.A2(n_1263),
.B1(n_1278),
.B2(n_1241),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1254),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1250),
.A2(n_1181),
.B1(n_1277),
.B2(n_1227),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1267),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1286),
.A2(n_1192),
.B1(n_1245),
.B2(n_1202),
.Y(n_1332)
);

CKINVDCx11_ASAP7_75t_R g1333 ( 
.A(n_1252),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1276),
.Y(n_1334)
);

NAND2x1p5_ASAP7_75t_L g1335 ( 
.A(n_1195),
.B(n_1248),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1196),
.B(n_1188),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1200),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1197),
.Y(n_1338)
);

OAI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1179),
.A2(n_1222),
.B1(n_1212),
.B2(n_1206),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1223),
.A2(n_1209),
.B1(n_1208),
.B2(n_1210),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1211),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1241),
.B(n_1251),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1205),
.B(n_1219),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1193),
.A2(n_1261),
.B1(n_1224),
.B2(n_1190),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1159),
.A2(n_1245),
.B1(n_1202),
.B2(n_1231),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_1216),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1213),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1251),
.A2(n_1279),
.B1(n_1159),
.B2(n_1199),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1224),
.A2(n_1220),
.B1(n_1177),
.B2(n_1203),
.Y(n_1349)
);

BUFx8_ASAP7_75t_L g1350 ( 
.A(n_1260),
.Y(n_1350)
);

BUFx2_ASAP7_75t_SL g1351 ( 
.A(n_1248),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1169),
.A2(n_1194),
.B1(n_1176),
.B2(n_1272),
.Y(n_1352)
);

INVx3_ASAP7_75t_SL g1353 ( 
.A(n_1272),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1218),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_1217),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1221),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1169),
.A2(n_1243),
.B1(n_1178),
.B2(n_1214),
.Y(n_1357)
);

CKINVDCx6p67_ASAP7_75t_R g1358 ( 
.A(n_1221),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1221),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1169),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1158),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1239),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_SL g1363 ( 
.A1(n_1230),
.A2(n_1259),
.B1(n_1275),
.B2(n_1285),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_SL g1364 ( 
.A1(n_1240),
.A2(n_1282),
.B1(n_1273),
.B2(n_1271),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1244),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1230),
.B(n_1285),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1215),
.Y(n_1367)
);

INVx4_ASAP7_75t_L g1368 ( 
.A(n_1246),
.Y(n_1368)
);

CKINVDCx14_ASAP7_75t_R g1369 ( 
.A(n_1259),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1253),
.Y(n_1370)
);

INVx6_ASAP7_75t_L g1371 ( 
.A(n_1185),
.Y(n_1371)
);

INVx4_ASAP7_75t_L g1372 ( 
.A(n_1249),
.Y(n_1372)
);

BUFx10_ASAP7_75t_L g1373 ( 
.A(n_1201),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1166),
.Y(n_1374)
);

OAI21xp33_ASAP7_75t_L g1375 ( 
.A1(n_1160),
.A2(n_1274),
.B(n_867),
.Y(n_1375)
);

BUFx8_ASAP7_75t_SL g1376 ( 
.A(n_1225),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1174),
.B(n_1256),
.Y(n_1377)
);

INVx6_ASAP7_75t_L g1378 ( 
.A(n_1249),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1173),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1162),
.A2(n_1255),
.B1(n_1274),
.B2(n_1160),
.Y(n_1380)
);

BUFx12f_ASAP7_75t_L g1381 ( 
.A(n_1185),
.Y(n_1381)
);

BUFx8_ASAP7_75t_L g1382 ( 
.A(n_1281),
.Y(n_1382)
);

OAI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1247),
.A2(n_1162),
.B1(n_1274),
.B2(n_1160),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1174),
.B(n_1256),
.Y(n_1384)
);

INVx1_ASAP7_75t_SL g1385 ( 
.A(n_1173),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1166),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1186),
.Y(n_1387)
);

BUFx2_ASAP7_75t_SL g1388 ( 
.A(n_1225),
.Y(n_1388)
);

INVxp67_ASAP7_75t_L g1389 ( 
.A(n_1163),
.Y(n_1389)
);

BUFx8_ASAP7_75t_L g1390 ( 
.A(n_1281),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1162),
.A2(n_1247),
.B1(n_867),
.B2(n_1160),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1162),
.A2(n_1255),
.B1(n_1274),
.B2(n_1160),
.Y(n_1392)
);

BUFx10_ASAP7_75t_L g1393 ( 
.A(n_1201),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1166),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1162),
.A2(n_1247),
.B1(n_867),
.B2(n_1160),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1162),
.A2(n_1247),
.B1(n_867),
.B2(n_1160),
.Y(n_1396)
);

CKINVDCx6p67_ASAP7_75t_R g1397 ( 
.A(n_1186),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1166),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1160),
.A2(n_903),
.B1(n_1274),
.B2(n_1247),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1162),
.A2(n_1255),
.B1(n_1274),
.B2(n_1160),
.Y(n_1400)
);

INVx4_ASAP7_75t_L g1401 ( 
.A(n_1249),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1341),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1338),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1369),
.B(n_1315),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1327),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1366),
.B(n_1360),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1361),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1322),
.B(n_1308),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1290),
.B(n_1319),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1380),
.A2(n_1400),
.B1(n_1392),
.B2(n_1383),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1363),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1323),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1304),
.Y(n_1413)
);

BUFx12f_ASAP7_75t_L g1414 ( 
.A(n_1289),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1367),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1342),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1342),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1293),
.B(n_1380),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1346),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1295),
.B(n_1294),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1331),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1334),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1337),
.Y(n_1423)
);

AO21x2_ASAP7_75t_L g1424 ( 
.A1(n_1352),
.A2(n_1357),
.B(n_1340),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1357),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1359),
.B(n_1336),
.Y(n_1426)
);

A2O1A1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1301),
.A2(n_1375),
.B(n_1399),
.C(n_1396),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1304),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1354),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1336),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1352),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1348),
.Y(n_1432)
);

BUFx2_ASAP7_75t_SL g1433 ( 
.A(n_1355),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1307),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1370),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1344),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1344),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1350),
.Y(n_1438)
);

AOI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1349),
.A2(n_1328),
.B(n_1309),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1345),
.A2(n_1313),
.B(n_1349),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1333),
.Y(n_1441)
);

INVx4_ASAP7_75t_L g1442 ( 
.A(n_1287),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1301),
.A2(n_1362),
.B(n_1328),
.Y(n_1443)
);

AOI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1303),
.A2(n_1377),
.B(n_1309),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1332),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1362),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1374),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1386),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_1350),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_1376),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1356),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_SL g1452 ( 
.A(n_1292),
.B(n_1296),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1313),
.B(n_1394),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1365),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1365),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1365),
.Y(n_1456)
);

OAI21xp33_ASAP7_75t_SL g1457 ( 
.A1(n_1391),
.A2(n_1395),
.B(n_1324),
.Y(n_1457)
);

AO21x2_ASAP7_75t_L g1458 ( 
.A1(n_1297),
.A2(n_1339),
.B(n_1343),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1335),
.A2(n_1312),
.B(n_1398),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1327),
.Y(n_1460)
);

BUFx2_ASAP7_75t_SL g1461 ( 
.A(n_1314),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1358),
.Y(n_1462)
);

OR2x6_ASAP7_75t_L g1463 ( 
.A(n_1368),
.B(n_1388),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1311),
.B(n_1324),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1384),
.B(n_1330),
.Y(n_1465)
);

NOR2x1_ASAP7_75t_L g1466 ( 
.A(n_1311),
.B(n_1401),
.Y(n_1466)
);

CKINVDCx20_ASAP7_75t_R g1467 ( 
.A(n_1325),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1302),
.B(n_1379),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1384),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1364),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1347),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1305),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1385),
.B(n_1318),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1351),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1385),
.B(n_1316),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1329),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1389),
.B(n_1353),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1321),
.B(n_1320),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1326),
.A2(n_1310),
.B1(n_1287),
.B2(n_1288),
.Y(n_1479)
);

INVx4_ASAP7_75t_L g1480 ( 
.A(n_1288),
.Y(n_1480)
);

AO21x2_ASAP7_75t_L g1481 ( 
.A1(n_1291),
.A2(n_1378),
.B(n_1288),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1387),
.B(n_1401),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1372),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1382),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1299),
.Y(n_1485)
);

OR2x2_ASAP7_75t_SL g1486 ( 
.A(n_1371),
.B(n_1317),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1314),
.A2(n_1373),
.B(n_1393),
.Y(n_1487)
);

BUFx12f_ASAP7_75t_L g1488 ( 
.A(n_1298),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1467),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1433),
.B(n_1300),
.Y(n_1490)
);

AO32x2_ASAP7_75t_L g1491 ( 
.A1(n_1479),
.A2(n_1373),
.A3(n_1393),
.B1(n_1382),
.B2(n_1390),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1406),
.B(n_1397),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1406),
.B(n_1306),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1410),
.A2(n_1371),
.B1(n_1381),
.B2(n_1427),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1457),
.B(n_1418),
.Y(n_1495)
);

AO32x2_ASAP7_75t_L g1496 ( 
.A1(n_1413),
.A2(n_1428),
.A3(n_1480),
.B1(n_1442),
.B2(n_1424),
.Y(n_1496)
);

OAI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1420),
.A2(n_1408),
.B(n_1466),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1420),
.A2(n_1408),
.B(n_1459),
.Y(n_1498)
);

A2O1A1Ixp33_ASAP7_75t_L g1499 ( 
.A1(n_1475),
.A2(n_1436),
.B(n_1437),
.C(n_1432),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1476),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1468),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1432),
.A2(n_1472),
.B1(n_1464),
.B2(n_1437),
.Y(n_1502)
);

A2O1A1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1436),
.A2(n_1404),
.B(n_1472),
.C(n_1445),
.Y(n_1503)
);

AO32x2_ASAP7_75t_L g1504 ( 
.A1(n_1413),
.A2(n_1428),
.A3(n_1442),
.B1(n_1480),
.B2(n_1424),
.Y(n_1504)
);

NAND4xp25_ASAP7_75t_L g1505 ( 
.A(n_1473),
.B(n_1465),
.C(n_1430),
.D(n_1425),
.Y(n_1505)
);

A2O1A1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1440),
.A2(n_1412),
.B(n_1411),
.C(n_1451),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1471),
.B(n_1451),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1458),
.A2(n_1426),
.B1(n_1411),
.B2(n_1412),
.Y(n_1508)
);

NOR2x1_ASAP7_75t_SL g1509 ( 
.A(n_1463),
.B(n_1481),
.Y(n_1509)
);

INVxp67_ASAP7_75t_L g1510 ( 
.A(n_1405),
.Y(n_1510)
);

OR2x6_ASAP7_75t_L g1511 ( 
.A(n_1463),
.B(n_1462),
.Y(n_1511)
);

OR2x6_ASAP7_75t_L g1512 ( 
.A(n_1463),
.B(n_1462),
.Y(n_1512)
);

O2A1O1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1458),
.A2(n_1460),
.B(n_1482),
.C(n_1403),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1426),
.B(n_1476),
.Y(n_1514)
);

AOI21xp33_ASAP7_75t_L g1515 ( 
.A1(n_1458),
.A2(n_1424),
.B(n_1470),
.Y(n_1515)
);

A2O1A1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1487),
.A2(n_1431),
.B(n_1409),
.C(n_1459),
.Y(n_1516)
);

AND2x4_ASAP7_75t_SL g1517 ( 
.A(n_1485),
.B(n_1441),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1421),
.B(n_1422),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1414),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1423),
.B(n_1477),
.Y(n_1520)
);

AO22x1_ASAP7_75t_SL g1521 ( 
.A1(n_1416),
.A2(n_1417),
.B1(n_1474),
.B2(n_1469),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1469),
.B(n_1434),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1447),
.B(n_1448),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1402),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1486),
.A2(n_1417),
.B1(n_1416),
.B2(n_1439),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1486),
.A2(n_1461),
.B1(n_1441),
.B2(n_1438),
.Y(n_1526)
);

AO21x2_ASAP7_75t_L g1527 ( 
.A1(n_1446),
.A2(n_1407),
.B(n_1455),
.Y(n_1527)
);

AO21x1_ASAP7_75t_L g1528 ( 
.A1(n_1415),
.A2(n_1483),
.B(n_1453),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1444),
.A2(n_1443),
.B(n_1446),
.Y(n_1529)
);

BUFx4f_ASAP7_75t_SL g1530 ( 
.A(n_1450),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1495),
.A2(n_1494),
.B1(n_1502),
.B2(n_1505),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1524),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1509),
.B(n_1454),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1529),
.B(n_1429),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1527),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1500),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1494),
.A2(n_1441),
.B1(n_1419),
.B2(n_1484),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1527),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1502),
.A2(n_1441),
.B1(n_1419),
.B2(n_1488),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1521),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1518),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1523),
.Y(n_1542)
);

INVx4_ASAP7_75t_L g1543 ( 
.A(n_1511),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1522),
.B(n_1498),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1496),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1521),
.Y(n_1546)
);

BUFx12f_ASAP7_75t_L g1547 ( 
.A(n_1519),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1528),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1498),
.B(n_1510),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1496),
.B(n_1435),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1496),
.B(n_1456),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1512),
.B(n_1456),
.Y(n_1552)
);

AO21x2_ASAP7_75t_L g1553 ( 
.A1(n_1535),
.A2(n_1515),
.B(n_1506),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1551),
.B(n_1504),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1532),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1532),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1533),
.B(n_1512),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1540),
.B(n_1513),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1545),
.B(n_1514),
.Y(n_1559)
);

INVx5_ASAP7_75t_SL g1560 ( 
.A(n_1552),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1551),
.B(n_1504),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1551),
.B(n_1504),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1533),
.Y(n_1563)
);

OAI31xp33_ASAP7_75t_L g1564 ( 
.A1(n_1531),
.A2(n_1503),
.A3(n_1525),
.B(n_1499),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1533),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1540),
.B(n_1516),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1546),
.B(n_1520),
.Y(n_1567)
);

CKINVDCx16_ASAP7_75t_R g1568 ( 
.A(n_1546),
.Y(n_1568)
);

AO21x2_ASAP7_75t_L g1569 ( 
.A1(n_1538),
.A2(n_1525),
.B(n_1497),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1550),
.B(n_1508),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1538),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1544),
.B(n_1505),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1547),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1544),
.B(n_1507),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1559),
.B(n_1549),
.Y(n_1575)
);

INVx4_ASAP7_75t_L g1576 ( 
.A(n_1573),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1555),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1565),
.B(n_1543),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1555),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1555),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1554),
.B(n_1548),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1571),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1563),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1554),
.B(n_1548),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1554),
.B(n_1541),
.Y(n_1585)
);

NAND2x1p5_ASAP7_75t_L g1586 ( 
.A(n_1557),
.B(n_1543),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1559),
.B(n_1549),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1554),
.B(n_1541),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1561),
.B(n_1541),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1566),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1571),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1556),
.Y(n_1592)
);

NAND4xp25_ASAP7_75t_L g1593 ( 
.A(n_1564),
.B(n_1531),
.C(n_1539),
.D(n_1537),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1559),
.B(n_1534),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1556),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1572),
.B(n_1542),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1572),
.B(n_1542),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1561),
.B(n_1562),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1572),
.B(n_1534),
.Y(n_1599)
);

NAND2x1p5_ASAP7_75t_L g1600 ( 
.A(n_1557),
.B(n_1543),
.Y(n_1600)
);

AOI221xp5_ASAP7_75t_L g1601 ( 
.A1(n_1593),
.A2(n_1558),
.B1(n_1566),
.B2(n_1564),
.C(n_1570),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1590),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1598),
.B(n_1568),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1599),
.B(n_1558),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1599),
.B(n_1574),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1582),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1582),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1590),
.B(n_1567),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1596),
.B(n_1597),
.Y(n_1609)
);

CKINVDCx16_ASAP7_75t_R g1610 ( 
.A(n_1576),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1596),
.B(n_1567),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1597),
.B(n_1536),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1598),
.B(n_1568),
.Y(n_1613)
);

NAND2x1_ASAP7_75t_L g1614 ( 
.A(n_1578),
.B(n_1563),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1576),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1585),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1576),
.B(n_1573),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1575),
.B(n_1574),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1591),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1598),
.B(n_1568),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1575),
.B(n_1536),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1591),
.Y(n_1622)
);

NAND3xp33_ASAP7_75t_SL g1623 ( 
.A(n_1586),
.B(n_1539),
.C(n_1537),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1577),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1593),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1581),
.B(n_1560),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1577),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1581),
.B(n_1560),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1579),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1579),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1580),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1580),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1592),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1581),
.B(n_1560),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1587),
.B(n_1570),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1592),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1578),
.B(n_1557),
.Y(n_1637)
);

AND3x2_ASAP7_75t_L g1638 ( 
.A(n_1578),
.B(n_1452),
.C(n_1490),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1584),
.B(n_1570),
.Y(n_1639)
);

INVxp67_ASAP7_75t_L g1640 ( 
.A(n_1584),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1595),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1606),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1624),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1601),
.B(n_1584),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1627),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1625),
.A2(n_1569),
.B1(n_1553),
.B2(n_1576),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1603),
.B(n_1586),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1602),
.B(n_1588),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1604),
.B(n_1594),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1603),
.B(n_1586),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1614),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1606),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1607),
.B(n_1588),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1613),
.B(n_1586),
.Y(n_1654)
);

INVxp67_ASAP7_75t_SL g1655 ( 
.A(n_1613),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1620),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1629),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1630),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1631),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1619),
.B(n_1589),
.Y(n_1660)
);

INVxp67_ASAP7_75t_L g1661 ( 
.A(n_1617),
.Y(n_1661)
);

INVx1_ASAP7_75t_SL g1662 ( 
.A(n_1615),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1608),
.B(n_1570),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1620),
.B(n_1578),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1626),
.B(n_1628),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1622),
.B(n_1589),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1616),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1604),
.B(n_1594),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1617),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1610),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1626),
.B(n_1600),
.Y(n_1671)
);

INVx1_ASAP7_75t_SL g1672 ( 
.A(n_1638),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1611),
.B(n_1612),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1632),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1633),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1636),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1616),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1637),
.B(n_1578),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1643),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1643),
.Y(n_1680)
);

OR2x6_ASAP7_75t_L g1681 ( 
.A(n_1661),
.B(n_1669),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1645),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1645),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1657),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1657),
.Y(n_1685)
);

INVxp67_ASAP7_75t_SL g1686 ( 
.A(n_1642),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1670),
.B(n_1547),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1662),
.B(n_1609),
.Y(n_1688)
);

INVxp67_ASAP7_75t_SL g1689 ( 
.A(n_1655),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1658),
.Y(n_1690)
);

INVx1_ASAP7_75t_SL g1691 ( 
.A(n_1672),
.Y(n_1691)
);

OAI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1644),
.A2(n_1672),
.B1(n_1656),
.B2(n_1623),
.Y(n_1692)
);

OAI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1644),
.A2(n_1639),
.B1(n_1635),
.B2(n_1605),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1658),
.Y(n_1694)
);

AOI211xp5_ASAP7_75t_SL g1695 ( 
.A1(n_1656),
.A2(n_1526),
.B(n_1640),
.C(n_1628),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_SL g1696 ( 
.A1(n_1646),
.A2(n_1641),
.B(n_1634),
.C(n_1621),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1662),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1656),
.A2(n_1569),
.B1(n_1553),
.B2(n_1634),
.Y(n_1698)
);

INVx1_ASAP7_75t_SL g1699 ( 
.A(n_1665),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1659),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1642),
.B(n_1609),
.Y(n_1701)
);

INVxp67_ASAP7_75t_SL g1702 ( 
.A(n_1642),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1663),
.A2(n_1569),
.B(n_1553),
.Y(n_1703)
);

NOR2x1_ASAP7_75t_L g1704 ( 
.A(n_1652),
.B(n_1441),
.Y(n_1704)
);

AOI211x1_ASAP7_75t_L g1705 ( 
.A1(n_1692),
.A2(n_1693),
.B(n_1703),
.C(n_1688),
.Y(n_1705)
);

XNOR2xp5_ASAP7_75t_L g1706 ( 
.A(n_1691),
.B(n_1517),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1697),
.B(n_1673),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1689),
.B(n_1652),
.Y(n_1708)
);

OAI322xp33_ASAP7_75t_L g1709 ( 
.A1(n_1699),
.A2(n_1652),
.A3(n_1668),
.B1(n_1649),
.B2(n_1666),
.C1(n_1660),
.C2(n_1653),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1681),
.B(n_1665),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1704),
.A2(n_1664),
.B1(n_1654),
.B2(n_1647),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1681),
.B(n_1687),
.Y(n_1712)
);

INVxp67_ASAP7_75t_L g1713 ( 
.A(n_1681),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1695),
.B(n_1664),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1701),
.B(n_1547),
.Y(n_1715)
);

NOR2xp67_ASAP7_75t_L g1716 ( 
.A(n_1679),
.B(n_1651),
.Y(n_1716)
);

AOI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1696),
.A2(n_1674),
.B1(n_1659),
.B2(n_1676),
.C(n_1675),
.Y(n_1717)
);

NAND2x1_ASAP7_75t_L g1718 ( 
.A(n_1680),
.B(n_1651),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1686),
.B(n_1664),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1686),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1702),
.B(n_1649),
.Y(n_1721)
);

AOI211x1_ASAP7_75t_SL g1722 ( 
.A1(n_1702),
.A2(n_1677),
.B(n_1667),
.C(n_1653),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1682),
.B(n_1547),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1683),
.Y(n_1724)
);

INVx1_ASAP7_75t_SL g1725 ( 
.A(n_1684),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1705),
.A2(n_1698),
.B1(n_1700),
.B2(n_1694),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1710),
.A2(n_1664),
.B1(n_1650),
.B2(n_1647),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1720),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1713),
.B(n_1685),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1708),
.B(n_1690),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1706),
.B(n_1488),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1721),
.Y(n_1732)
);

NOR2xp67_ASAP7_75t_L g1733 ( 
.A(n_1711),
.B(n_1651),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1718),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1712),
.B(n_1650),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1731),
.B(n_1707),
.Y(n_1736)
);

NOR3xp33_ASAP7_75t_L g1737 ( 
.A(n_1726),
.B(n_1715),
.C(n_1714),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1732),
.B(n_1719),
.Y(n_1738)
);

OAI211xp5_ASAP7_75t_L g1739 ( 
.A1(n_1726),
.A2(n_1717),
.B(n_1725),
.C(n_1724),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1735),
.B(n_1724),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1733),
.B(n_1716),
.Y(n_1741)
);

AOI211xp5_ASAP7_75t_L g1742 ( 
.A1(n_1729),
.A2(n_1723),
.B(n_1709),
.C(n_1725),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1728),
.B(n_1722),
.Y(n_1743)
);

INVx2_ASAP7_75t_SL g1744 ( 
.A(n_1734),
.Y(n_1744)
);

AOI221xp5_ASAP7_75t_L g1745 ( 
.A1(n_1739),
.A2(n_1737),
.B1(n_1742),
.B2(n_1743),
.C(n_1744),
.Y(n_1745)
);

NOR4xp25_ASAP7_75t_L g1746 ( 
.A(n_1738),
.B(n_1740),
.C(n_1741),
.D(n_1730),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1736),
.B(n_1727),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1737),
.A2(n_1654),
.B1(n_1671),
.B2(n_1678),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1744),
.B(n_1674),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1745),
.A2(n_1746),
.B1(n_1747),
.B2(n_1749),
.C(n_1748),
.Y(n_1750)
);

OAI211xp5_ASAP7_75t_SL g1751 ( 
.A1(n_1745),
.A2(n_1478),
.B(n_1651),
.C(n_1648),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1746),
.B(n_1668),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1749),
.Y(n_1753)
);

AOI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1745),
.A2(n_1675),
.B1(n_1676),
.B2(n_1667),
.C(n_1677),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1749),
.Y(n_1755)
);

NAND3x1_ASAP7_75t_SL g1756 ( 
.A(n_1750),
.B(n_1414),
.C(n_1671),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1752),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1755),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1753),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1754),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_L g1761 ( 
.A(n_1757),
.B(n_1751),
.C(n_1677),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1760),
.B(n_1648),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1758),
.B(n_1660),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1763),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1764),
.A2(n_1761),
.B1(n_1762),
.B2(n_1759),
.Y(n_1765)
);

INVx1_ASAP7_75t_SL g1766 ( 
.A(n_1765),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_SL g1767 ( 
.A1(n_1765),
.A2(n_1756),
.B1(n_1530),
.B2(n_1449),
.Y(n_1767)
);

OA21x2_ASAP7_75t_L g1768 ( 
.A1(n_1766),
.A2(n_1667),
.B(n_1678),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_SL g1769 ( 
.A1(n_1767),
.A2(n_1438),
.B1(n_1449),
.B2(n_1678),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1769),
.A2(n_1678),
.B1(n_1666),
.B2(n_1637),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1770),
.B(n_1768),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_SL g1772 ( 
.A1(n_1771),
.A2(n_1493),
.B(n_1492),
.Y(n_1772)
);

OAI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1772),
.A2(n_1614),
.B1(n_1489),
.B2(n_1605),
.Y(n_1773)
);

OAI221xp5_ASAP7_75t_R g1774 ( 
.A1(n_1773),
.A2(n_1637),
.B1(n_1491),
.B2(n_1583),
.C(n_1618),
.Y(n_1774)
);

AOI211xp5_ASAP7_75t_L g1775 ( 
.A1(n_1774),
.A2(n_1482),
.B(n_1501),
.C(n_1618),
.Y(n_1775)
);


endmodule