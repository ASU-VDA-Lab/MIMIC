module real_jpeg_13318_n_11 (n_5, n_4, n_8, n_0, n_39, n_40, n_1, n_2, n_38, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_39;
input n_40;
input n_1;
input n_2;
input n_38;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_17;
wire n_21;
wire n_33;
wire n_35;
wire n_29;
wire n_31;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_36;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_L g36 ( 
.A(n_0),
.B(n_1),
.C(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

NAND3xp33_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_4),
.C(n_14),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_2),
.A2(n_4),
.B(n_14),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_3),
.B(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_5),
.A2(n_14),
.B(n_38),
.Y(n_22)
);

NAND3xp33_ASAP7_75t_L g26 ( 
.A(n_5),
.B(n_14),
.C(n_40),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_7),
.A2(n_9),
.B(n_14),
.Y(n_19)
);

NAND3xp33_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_9),
.C(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_8),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_8),
.A2(n_28),
.B(n_29),
.Y(n_27)
);

NOR3xp33_ASAP7_75t_L g30 ( 
.A(n_8),
.B(n_28),
.C(n_29),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_8),
.A2(n_33),
.B(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_17),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_15),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_32),
.B(n_35),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B(n_31),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_27),
.B(n_30),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B(n_26),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_39),
.Y(n_25)
);


endmodule