module fake_jpeg_30029_n_188 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_188);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_1),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx6p67_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_13),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_17),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_21),
.B1(n_24),
.B2(n_20),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_41),
.B1(n_39),
.B2(n_23),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_62),
.Y(n_79)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_14),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_28),
.B1(n_15),
.B2(n_18),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_39),
.B1(n_24),
.B2(n_20),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_27),
.Y(n_58)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_22),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_14),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_37),
.B1(n_31),
.B2(n_33),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_78),
.B1(n_80),
.B2(n_93),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_42),
.B(n_19),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_52),
.C(n_2),
.Y(n_111)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_87),
.Y(n_99)
);

AO22x2_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_33),
.B1(n_31),
.B2(n_39),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_59),
.B(n_56),
.C(n_52),
.Y(n_104)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_85),
.B(n_55),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_39),
.B1(n_35),
.B2(n_24),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_41),
.B(n_34),
.C(n_35),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_88),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_91),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_25),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_49),
.A2(n_34),
.B1(n_21),
.B2(n_19),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_94),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_75),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_100),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_46),
.B(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_71),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_85),
.B1(n_68),
.B2(n_94),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_75),
.A2(n_49),
.B1(n_54),
.B2(n_18),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_96),
.B1(n_104),
.B2(n_85),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_52),
.B(n_2),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_111),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_52),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_66),
.C(n_85),
.Y(n_132)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_120),
.A2(n_126),
.B(n_132),
.Y(n_138)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_124),
.B(n_130),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_72),
.B(n_68),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_79),
.B(n_117),
.Y(n_139)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_125),
.B(n_131),
.C(n_127),
.D(n_130),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_68),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_131),
.Y(n_136)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_68),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_110),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_134),
.A2(n_117),
.B1(n_95),
.B2(n_104),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_113),
.C(n_99),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_98),
.C(n_69),
.Y(n_159)
);

AOI221xp5_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_120),
.B1(n_119),
.B2(n_115),
.C(n_98),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_144),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_107),
.Y(n_141)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_127),
.C(n_138),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_154),
.C(n_155),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_120),
.B1(n_134),
.B2(n_132),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_151),
.A2(n_157),
.B1(n_158),
.B2(n_106),
.Y(n_168)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_136),
.A2(n_120),
.B(n_123),
.C(n_133),
.D(n_121),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_136),
.C(n_139),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_102),
.C(n_114),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_102),
.C(n_97),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_119),
.B1(n_115),
.B2(n_108),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_146),
.C(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_163),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_167),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_140),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_146),
.B(n_140),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_157),
.B(n_159),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_150),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_151),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_108),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_166),
.A2(n_165),
.B1(n_164),
.B2(n_161),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_82),
.C(n_88),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_84),
.B1(n_100),
.B2(n_3),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_5),
.B(n_6),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_171),
.A2(n_1),
.B(n_3),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_172),
.A2(n_174),
.B1(n_4),
.B2(n_5),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_160),
.C(n_2),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_177),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_179),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_3),
.C(n_4),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_169),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_170),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_181),
.C(n_7),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_171),
.B(n_8),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_184),
.A2(n_7),
.B(n_9),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_186),
.C(n_7),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_9),
.Y(n_188)
);


endmodule