module real_jpeg_32006_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_648;
wire n_95;
wire n_541;
wire n_441;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_669;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_611;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_653;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_412;
wire n_155;
wire n_405;
wire n_586;
wire n_572;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_642;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g210 ( 
.A(n_0),
.Y(n_210)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_0),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g258 ( 
.A(n_0),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_0),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_1),
.A2(n_131),
.B(n_134),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_1),
.B(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_1),
.Y(n_236)
);

OAI32xp33_ASAP7_75t_L g431 ( 
.A1(n_1),
.A2(n_100),
.A3(n_432),
.B1(n_436),
.B2(n_439),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_1),
.A2(n_236),
.B1(n_473),
.B2(n_478),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_1),
.B(n_117),
.Y(n_531)
);

OAI22xp33_ASAP7_75t_SL g565 ( 
.A1(n_1),
.A2(n_209),
.B1(n_552),
.B2(n_566),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_2),
.A2(n_184),
.B1(n_187),
.B2(n_191),
.Y(n_183)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_2),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_2),
.A2(n_191),
.B1(n_213),
.B2(n_217),
.Y(n_212)
);

AO22x1_ASAP7_75t_L g319 ( 
.A1(n_2),
.A2(n_191),
.B1(n_320),
.B2(n_322),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_2),
.A2(n_138),
.B1(n_191),
.B2(n_408),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_3),
.A2(n_21),
.B(n_22),
.Y(n_20)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_5),
.A2(n_138),
.B1(n_141),
.B2(n_142),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_5),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_5),
.A2(n_141),
.B1(n_199),
.B2(n_202),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_5),
.A2(n_141),
.B1(n_509),
.B2(n_511),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_5),
.A2(n_141),
.B1(n_553),
.B2(n_555),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_6),
.A2(n_226),
.B1(n_227),
.B2(n_231),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_6),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_6),
.A2(n_226),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_6),
.A2(n_226),
.B1(n_362),
.B2(n_364),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_SL g610 ( 
.A1(n_6),
.A2(n_226),
.B1(n_611),
.B2(n_612),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_7),
.A2(n_52),
.B1(n_56),
.B2(n_59),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_7),
.A2(n_59),
.B1(n_262),
.B2(n_339),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_7),
.A2(n_59),
.B1(n_391),
.B2(n_393),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g648 ( 
.A1(n_7),
.A2(n_59),
.B1(n_649),
.B2(n_653),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_8),
.A2(n_173),
.B1(n_176),
.B2(n_180),
.Y(n_172)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_8),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_8),
.A2(n_180),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_8),
.A2(n_180),
.B1(n_370),
.B2(n_372),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_8),
.A2(n_180),
.B1(n_448),
.B2(n_451),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_9),
.A2(n_120),
.B1(n_121),
.B2(n_125),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_9),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_9),
.A2(n_120),
.B1(n_313),
.B2(n_315),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_9),
.A2(n_120),
.B1(n_176),
.B2(n_429),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_9),
.A2(n_120),
.B1(n_279),
.B2(n_521),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_10),
.A2(n_261),
.B1(n_262),
.B2(n_265),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_10),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_10),
.A2(n_261),
.B1(n_273),
.B2(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_10),
.A2(n_261),
.B1(n_400),
.B2(n_402),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_SL g641 ( 
.A1(n_10),
.A2(n_52),
.B1(n_261),
.B2(n_642),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_11),
.A2(n_63),
.B1(n_67),
.B2(n_71),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_11),
.A2(n_71),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_11),
.A2(n_71),
.B1(n_177),
.B2(n_274),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_11),
.A2(n_71),
.B1(n_474),
.B2(n_622),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_13),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_13),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_14),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_14),
.Y(n_220)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_14),
.Y(n_234)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_14),
.Y(n_525)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_15),
.Y(n_151)
);

CKINVDCx11_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_16),
.B(n_678),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_17),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_17),
.A2(n_87),
.B1(n_138),
.B2(n_289),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_17),
.A2(n_87),
.B1(n_274),
.B2(n_483),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_SL g539 ( 
.A1(n_17),
.A2(n_87),
.B1(n_540),
.B2(n_543),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_18),
.Y(n_110)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_18),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_18),
.Y(n_160)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_19),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_19),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_72),
.B(n_677),
.Y(n_22)
);

INVxp67_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_60),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_26),
.B(n_680),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_38),
.B(n_51),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_27),
.A2(n_38),
.B1(n_51),
.B2(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_27),
.A2(n_38),
.B1(n_130),
.B2(n_137),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_27),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_27),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_27),
.A2(n_38),
.B1(n_288),
.B2(n_312),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_27),
.A2(n_38),
.B1(n_312),
.B2(n_368),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g639 ( 
.A1(n_27),
.A2(n_38),
.B1(n_640),
.B2(n_641),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_SL g666 ( 
.A1(n_27),
.A2(n_38),
.B1(n_62),
.B2(n_641),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_28)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_29),
.Y(n_401)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_30),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_30),
.Y(n_477)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_39),
.A2(n_286),
.B1(n_287),
.B2(n_293),
.Y(n_285)
);

AO22x1_ASAP7_75t_L g406 ( 
.A1(n_39),
.A2(n_286),
.B1(n_369),
.B2(n_407),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_39),
.A2(n_286),
.B1(n_407),
.B2(n_610),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_43),
.Y(n_140)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_43),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_43),
.Y(n_314)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_46),
.Y(n_243)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_47),
.Y(n_133)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_48),
.Y(n_136)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_50),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_54),
.Y(n_144)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_55),
.Y(n_247)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_60),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_61),
.B(n_669),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_61),
.B(n_669),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_66),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_66),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_70),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_596),
.B(n_670),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_420),
.B(n_587),
.Y(n_74)
);

NAND4xp25_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_305),
.C(n_378),
.D(n_412),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_268),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_77),
.B(n_268),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_194),
.C(n_237),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_78),
.B(n_584),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_128),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_79),
.B(n_192),
.C(n_193),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_91),
.B1(n_117),
.B2(n_118),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g196 ( 
.A1(n_81),
.A2(n_92),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_86),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_86),
.Y(n_652)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_90),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_91),
.A2(n_117),
.B1(n_319),
.B2(n_325),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_91),
.A2(n_117),
.B1(n_319),
.B2(n_325),
.Y(n_344)
);

AOI22x1_ASAP7_75t_L g360 ( 
.A1(n_91),
.A2(n_117),
.B1(n_319),
.B2(n_361),
.Y(n_360)
);

AOI22x1_ASAP7_75t_L g398 ( 
.A1(n_91),
.A2(n_117),
.B1(n_361),
.B2(n_399),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_91),
.A2(n_117),
.B(n_665),
.Y(n_664)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_92),
.A2(n_119),
.B1(n_197),
.B2(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_92),
.A2(n_197),
.B1(n_198),
.B2(n_472),
.Y(n_471)
);

OA22x2_ASAP7_75t_L g620 ( 
.A1(n_92),
.A2(n_197),
.B1(n_621),
.B2(n_626),
.Y(n_620)
);

OA22x2_ASAP7_75t_L g647 ( 
.A1(n_92),
.A2(n_197),
.B1(n_621),
.B2(n_648),
.Y(n_647)
);

AO21x2_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_100),
.B(n_108),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_101),
.Y(n_297)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_102),
.Y(n_240)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_102),
.Y(n_625)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_103),
.Y(n_253)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_111),
.B1(n_113),
.B2(n_115),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_114),
.Y(n_438)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_117),
.Y(n_197)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_124),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_145),
.B1(n_192),
.B2(n_193),
.Y(n_128)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_134),
.Y(n_254)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_137),
.Y(n_293)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_138),
.Y(n_611)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_140),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_172),
.B1(n_181),
.B2(n_183),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_146),
.A2(n_181),
.B1(n_183),
.B2(n_272),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_146),
.A2(n_181),
.B1(n_272),
.B2(n_332),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_146),
.A2(n_181),
.B1(n_332),
.B2(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_146),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_146),
.A2(n_172),
.B1(n_426),
.B2(n_427),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_146),
.A2(n_181),
.B1(n_482),
.B2(n_507),
.Y(n_532)
);

AO21x2_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_156),
.B(n_164),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g618 ( 
.A(n_147),
.Y(n_618)
);

NAND2xp67_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_165),
.B1(n_168),
.B2(n_170),
.Y(n_164)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_150),
.Y(n_500)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_155),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_156),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_159),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_160),
.Y(n_335)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_160),
.Y(n_396)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

INVxp33_ASAP7_75t_SL g619 ( 
.A(n_164),
.Y(n_619)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_167),
.Y(n_216)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_169),
.Y(n_280)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_179),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_181),
.Y(n_397)
);

AOI21x1_ASAP7_75t_L g616 ( 
.A1(n_181),
.A2(n_390),
.B(n_617),
.Y(n_616)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_186),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_190),
.Y(n_392)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_190),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_195),
.B(n_237),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_206),
.C(n_235),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_196),
.B(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_205),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_206),
.A2(n_207),
.B1(n_235),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_212),
.B1(n_221),
.B2(n_225),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_208),
.A2(n_225),
.B1(n_256),
.B2(n_259),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_208),
.A2(n_352),
.B(n_353),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_208),
.A2(n_212),
.B1(n_447),
.B2(n_455),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_208),
.A2(n_538),
.B1(n_544),
.B2(n_545),
.Y(n_537)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_209),
.A2(n_260),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_209),
.A2(n_278),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_209),
.A2(n_520),
.B1(n_526),
.B2(n_529),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_209),
.A2(n_539),
.B1(n_552),
.B2(n_559),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_216),
.Y(n_493)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx2_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_219),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_220),
.Y(n_498)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_220),
.Y(n_558)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_223),
.Y(n_570)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_224),
.Y(n_562)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_231),
.Y(n_279)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_232),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_233),
.Y(n_554)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_234),
.Y(n_264)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_234),
.Y(n_450)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_234),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_234),
.Y(n_542)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_235),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_236),
.B(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_236),
.B(n_502),
.Y(n_501)
);

OA21x2_ASAP7_75t_SL g513 ( 
.A1(n_236),
.A2(n_501),
.B(n_514),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g563 ( 
.A(n_236),
.B(n_426),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_236),
.B(n_569),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_255),
.B1(n_266),
.B2(n_267),
.Y(n_237)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

OAI32xp33_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_241),
.A3(n_244),
.B1(n_248),
.B2(n_254),
.Y(n_238)
);

OAI32xp33_ASAP7_75t_L g304 ( 
.A1(n_239),
.A2(n_241),
.A3(n_244),
.B1(n_248),
.B2(n_254),
.Y(n_304)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_256),
.Y(n_277)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx8_ASAP7_75t_L g337 ( 
.A(n_258),
.Y(n_337)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_265),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_267),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_267),
.B(n_304),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_282),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_281),
.Y(n_269)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_270),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_276),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_271),
.B(n_276),
.Y(n_309)
);

BUFx6f_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_281),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_282),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_303),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_294),
.B2(n_295),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_285),
.Y(n_328)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_294),
.B(n_327),
.C(n_328),
.Y(n_326)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_296),
.Y(n_325)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_300),
.Y(n_365)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_301),
.Y(n_403)
);

INVx8_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_302),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_340),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_306),
.A2(n_340),
.B1(n_413),
.B2(n_589),
.Y(n_590)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_306),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_326),
.C(n_329),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_307),
.B(n_330),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_343),
.C(n_344),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_318),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_311),
.Y(n_343)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_314),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_326),
.Y(n_418)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_336),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_331),
.B(n_336),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_337),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_338),
.Y(n_353)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_340),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_355),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_345),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_345),
.C(n_356),
.Y(n_379)
);

OAI21x1_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_350),
.B(n_354),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NAND2xp33_ASAP7_75t_SL g604 ( 
.A(n_347),
.B(n_350),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_348),
.B(n_351),
.Y(n_354)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_349),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_SL g603 ( 
.A1(n_350),
.A2(n_604),
.B(n_605),
.Y(n_603)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2x1_ASAP7_75t_L g405 ( 
.A(n_354),
.B(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_376),
.B2(n_377),
.Y(n_356)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_357),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_358),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_366),
.B2(n_367),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_376),
.C(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_367),
.Y(n_382)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_375),
.Y(n_645)
);

A2O1A1Ixp33_ASAP7_75t_L g587 ( 
.A1(n_378),
.A2(n_588),
.B(n_590),
.C(n_591),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_379),
.B(n_380),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_383),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_381),
.B(n_600),
.C(n_601),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_385),
.B1(n_405),
.B2(n_411),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_384),
.Y(n_600)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_398),
.B(n_404),
.Y(n_385)
);

NAND2x1p5_ASAP7_75t_L g404 ( 
.A(n_386),
.B(n_398),
.Y(n_404)
);

AOI22x1_ASAP7_75t_SL g386 ( 
.A1(n_387),
.A2(n_388),
.B1(n_389),
.B2(n_397),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_388),
.A2(n_397),
.B1(n_428),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_388),
.Y(n_512)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx4f_ASAP7_75t_L g510 ( 
.A(n_394),
.Y(n_510)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_396),
.Y(n_517)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_397),
.Y(n_426)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_399),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_404),
.B(n_607),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_404),
.B(n_603),
.C(n_632),
.Y(n_631)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_405),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_405),
.Y(n_601)
);

INVxp67_ASAP7_75t_SL g605 ( 
.A(n_406),
.Y(n_605)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_417),
.Y(n_412)
);

OAI21xp33_ASAP7_75t_L g588 ( 
.A1(n_413),
.A2(n_417),
.B(n_589),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.C(n_416),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.Y(n_417)
);

AOI21x1_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_582),
.B(n_586),
.Y(n_420)
);

OAI21x1_ASAP7_75t_SL g421 ( 
.A1(n_422),
.A2(n_487),
.B(n_581),
.Y(n_421)
);

AOI211xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_461),
.B(n_466),
.C(n_467),
.Y(n_422)
);

A2O1A1Ixp33_ASAP7_75t_L g581 ( 
.A1(n_423),
.A2(n_461),
.B(n_466),
.C(n_467),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_424),
.B(n_463),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_430),
.B1(n_459),
.B2(n_460),
.Y(n_424)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_425),
.B(n_459),
.C(n_462),
.Y(n_585)
);

OAI22x1_ASAP7_75t_L g506 ( 
.A1(n_426),
.A2(n_507),
.B1(n_512),
.B2(n_513),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_430),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_445),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_431),
.A2(n_445),
.B1(n_446),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_431),
.Y(n_469)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_443),
.Y(n_505)
);

INVx5_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_444),
.Y(n_486)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_447),
.Y(n_529)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_453),
.Y(n_571)
);

BUFx12f_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_458),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_458),
.Y(n_547)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_470),
.C(n_480),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_468),
.B(n_578),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_470),
.A2(n_471),
.B1(n_480),
.B2(n_579),
.Y(n_578)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_480),
.Y(n_579)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_486),
.Y(n_485)
);

AOI21x1_ASAP7_75t_L g487 ( 
.A1(n_488),
.A2(n_575),
.B(n_580),
.Y(n_487)
);

OAI21x1_ASAP7_75t_SL g488 ( 
.A1(n_489),
.A2(n_535),
.B(n_574),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_518),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_490),
.B(n_518),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_506),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g548 ( 
.A(n_491),
.B(n_506),
.Y(n_548)
);

AO21x1_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_494),
.B(n_495),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_494),
.A2(n_618),
.B(n_619),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_496),
.A2(n_499),
.B(n_501),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_530),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_519),
.B(n_532),
.C(n_533),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_520),
.Y(n_544)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_531),
.A2(n_532),
.B1(n_533),
.B2(n_534),
.Y(n_530)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_531),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_532),
.Y(n_534)
);

AOI21x1_ASAP7_75t_L g535 ( 
.A1(n_536),
.A2(n_549),
.B(n_573),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_548),
.Y(n_536)
);

NOR2xp67_ASAP7_75t_L g573 ( 
.A(n_537),
.B(n_548),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx3_ASAP7_75t_SL g545 ( 
.A(n_546),
.Y(n_545)
);

INVx8_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_550),
.A2(n_564),
.B(n_572),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_551),
.B(n_563),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_551),
.B(n_563),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_560),
.Y(n_566)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_562),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_565),
.B(n_567),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g567 ( 
.A(n_568),
.B(n_571),
.Y(n_567)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_576),
.B(n_577),
.Y(n_575)
);

NOR2xp67_ASAP7_75t_SL g580 ( 
.A(n_576),
.B(n_577),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_583),
.B(n_585),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_583),
.B(n_585),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_592),
.B(n_595),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_593),
.B(n_594),
.Y(n_592)
);

NAND3xp33_ASAP7_75t_L g596 ( 
.A(n_597),
.B(n_656),
.C(n_668),
.Y(n_596)
);

NOR2xp67_ASAP7_75t_SL g597 ( 
.A(n_598),
.B(n_629),
.Y(n_597)
);

NOR2xp67_ASAP7_75t_L g598 ( 
.A(n_599),
.B(n_602),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_599),
.B(n_602),
.Y(n_673)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_603),
.B(n_606),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_607),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_608),
.B(n_614),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_609),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_610),
.Y(n_640)
);

INVx4_ASAP7_75t_SL g612 ( 
.A(n_613),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_615),
.A2(n_620),
.B(n_627),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g660 ( 
.A(n_615),
.B(n_639),
.C(n_661),
.Y(n_660)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_616),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_616),
.B(n_635),
.C(n_636),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_SL g646 ( 
.A(n_616),
.B(n_647),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_620),
.B(n_628),
.Y(n_627)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_620),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_623),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_624),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

AOI21x1_ASAP7_75t_SL g672 ( 
.A1(n_630),
.A2(n_673),
.B(n_674),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_631),
.B(n_633),
.Y(n_630)
);

NOR2xp67_ASAP7_75t_SL g674 ( 
.A(n_631),
.B(n_633),
.Y(n_674)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_634),
.B(n_637),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g667 ( 
.A(n_634),
.B(n_635),
.C(n_638),
.Y(n_667)
);

XNOR2xp5_ASAP7_75t_L g637 ( 
.A(n_635),
.B(n_638),
.Y(n_637)
);

XNOR2x1_ASAP7_75t_L g638 ( 
.A(n_639),
.B(n_646),
.Y(n_638)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_643),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_644),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_645),
.Y(n_644)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_647),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_648),
.Y(n_665)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_651),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_652),
.Y(n_651)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_654),
.Y(n_653)
);

INVx8_ASAP7_75t_L g654 ( 
.A(n_655),
.Y(n_654)
);

INVxp33_ASAP7_75t_SL g656 ( 
.A(n_657),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_SL g671 ( 
.A1(n_657),
.A2(n_672),
.B(n_675),
.Y(n_671)
);

NOR2x1_ASAP7_75t_R g657 ( 
.A(n_658),
.B(n_667),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_658),
.B(n_667),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_SL g658 ( 
.A1(n_659),
.A2(n_660),
.B1(n_662),
.B2(n_663),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_659),
.B(n_664),
.C(n_666),
.Y(n_669)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_660),
.Y(n_659)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_663),
.Y(n_662)
);

XOR2xp5_ASAP7_75t_L g663 ( 
.A(n_664),
.B(n_666),
.Y(n_663)
);

AOI21xp33_ASAP7_75t_SL g670 ( 
.A1(n_668),
.A2(n_671),
.B(n_676),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_679),
.Y(n_678)
);


endmodule