module fake_jpeg_16300_n_38 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx12_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_15),
.B(n_18),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_1),
.Y(n_16)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_16),
.B(n_17),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_1),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_8),
.A2(n_6),
.B1(n_2),
.B2(n_3),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_14),
.B(n_15),
.Y(n_21)
);

NOR2x1p5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_26),
.B1(n_8),
.B2(n_13),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_17),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_16),
.C(n_18),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_7),
.C(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_19),
.B(n_12),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_29),
.C(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_35),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_32),
.B(n_11),
.C(n_19),
.Y(n_38)
);


endmodule