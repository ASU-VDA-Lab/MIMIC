module fake_netlist_1_7857_n_28 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_28);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
CKINVDCx20_ASAP7_75t_R g8 ( .A(n_7), .Y(n_8) );
NOR2xp33_ASAP7_75t_R g9 ( .A(n_2), .B(n_6), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_3), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_5), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_0), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_12), .B(n_1), .Y(n_16) );
INVx5_ASAP7_75t_L g17 ( .A(n_9), .Y(n_17) );
BUFx3_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_16), .A2(n_10), .B(n_11), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_17), .Y(n_21) );
NAND2x1p5_ASAP7_75t_L g22 ( .A(n_18), .B(n_17), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_20), .B(n_8), .Y(n_23) );
OR2x2_ASAP7_75t_L g24 ( .A(n_22), .B(n_19), .Y(n_24) );
NOR2xp33_ASAP7_75t_R g25 ( .A(n_24), .B(n_21), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_23), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
endmodule