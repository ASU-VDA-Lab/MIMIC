module real_jpeg_6236_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_1),
.B(n_261),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_1),
.A2(n_120),
.B(n_260),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_1),
.B(n_193),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_1),
.B(n_370),
.C(n_373),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_L g375 ( 
.A1(n_1),
.A2(n_45),
.B1(n_376),
.B2(n_377),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_1),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_1),
.B(n_90),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_1),
.A2(n_143),
.B1(n_413),
.B2(n_421),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_2),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_2),
.A2(n_48),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_2),
.A2(n_48),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_2),
.A2(n_48),
.B1(n_94),
.B2(n_187),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_3),
.A2(n_65),
.B1(n_70),
.B2(n_71),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_3),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_3),
.A2(n_70),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_3),
.A2(n_70),
.B1(n_226),
.B2(n_229),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_3),
.A2(n_70),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_4),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_5),
.A2(n_173),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_5),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_5),
.A2(n_106),
.B1(n_255),
.B2(n_292),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_5),
.A2(n_292),
.B1(n_388),
.B2(n_390),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g401 ( 
.A1(n_5),
.A2(n_292),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_6),
.A2(n_45),
.B1(n_59),
.B2(n_61),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_6),
.A2(n_61),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_6),
.A2(n_61),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_6),
.A2(n_61),
.B1(n_144),
.B2(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_7),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_18)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_9),
.A2(n_92),
.B1(n_93),
.B2(n_97),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_9),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_9),
.A2(n_92),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_9),
.A2(n_92),
.B1(n_195),
.B2(n_198),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_9),
.A2(n_92),
.B1(n_274),
.B2(n_276),
.Y(n_273)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_10),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_10),
.Y(n_151)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_10),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_10),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_10),
.Y(n_308)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_11),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_11),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_11),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_11),
.Y(n_139)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_11),
.Y(n_258)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_14),
.Y(n_118)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_14),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_14),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_14),
.Y(n_133)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_14),
.Y(n_136)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_14),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_14),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_14),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g234 ( 
.A(n_14),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_14),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_15),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_15),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_15),
.A2(n_97),
.B1(n_235),
.B2(n_282),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_15),
.A2(n_145),
.B1(n_235),
.B2(n_396),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_15),
.A2(n_165),
.B1(n_235),
.B2(n_453),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_16),
.A2(n_173),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_16),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_16),
.A2(n_72),
.B1(n_289),
.B2(n_339),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_16),
.A2(n_165),
.B1(n_289),
.B2(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_16),
.A2(n_289),
.B1(n_414),
.B2(n_416),
.Y(n_413)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_17),
.Y(n_372)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_201),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_199),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_176),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_27),
.B(n_176),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_27),
.B(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_27),
.B(n_203),
.Y(n_482)
);

FAx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_98),
.CI(n_141),
.CON(n_27),
.SN(n_27)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_28),
.A2(n_29),
.B(n_62),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_62),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_51),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_30),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_44),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_31),
.A2(n_44),
.B(n_52),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_31),
.A2(n_52),
.B1(n_57),
.B2(n_225),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_31),
.B(n_376),
.Y(n_411)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_32),
.B(n_58),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_32),
.A2(n_53),
.B1(n_163),
.B2(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_32),
.A2(n_53),
.B1(n_375),
.B2(n_378),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_32),
.A2(n_53),
.B1(n_378),
.B2(n_387),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_32),
.A2(n_53),
.B1(n_387),
.B2(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_41),
.B1(n_46),
.B2(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_35),
.Y(n_373)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_37),
.Y(n_217)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_40),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_40),
.Y(n_275)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_44),
.A2(n_52),
.B(n_168),
.Y(n_295)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_49),
.Y(n_445)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_52),
.A2(n_162),
.B(n_168),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_52),
.A2(n_465),
.B(n_466),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_55),
.Y(n_392)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_56),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_56),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_56),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_56),
.Y(n_389)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_75),
.B1(n_90),
.B2(n_91),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_64),
.A2(n_76),
.B(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_84),
.B1(n_86),
.B2(n_88),
.Y(n_83)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_69),
.Y(n_285)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_69),
.Y(n_341)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_73),
.A2(n_96),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_74),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_74),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g450 ( 
.A(n_74),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_91),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_75),
.B(n_105),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_75),
.A2(n_185),
.B(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_75),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_75),
.A2(n_90),
.B1(n_338),
.B2(n_449),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_83),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_76),
.B(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_76),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_76),
.A2(n_300),
.B1(n_301),
.B2(n_337),
.Y(n_336)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_81),
.B2(n_82),
.Y(n_76)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_77),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_77),
.Y(n_377)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_78),
.Y(n_444)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_80),
.Y(n_438)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_96),
.Y(n_442)
);

OAI32xp33_ASAP7_75t_L g433 ( 
.A1(n_97),
.A2(n_434),
.A3(n_436),
.B1(n_439),
.B2(n_443),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_111),
.B2(n_140),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_109),
.B2(n_110),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_101),
.A2(n_110),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_102),
.B(n_110),
.C(n_111),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_104),
.A2(n_186),
.B(n_301),
.Y(n_319)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_106),
.Y(n_255)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_111),
.A2(n_140),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_116),
.B(n_123),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_112),
.B(n_125),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_112),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_112),
.A2(n_130),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_112),
.A2(n_130),
.B1(n_232),
.B2(n_291),
.Y(n_320)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_115),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_118),
.Y(n_251)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_128),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_129),
.A2(n_170),
.B(n_175),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_129),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_129),
.A2(n_193),
.B1(n_287),
.B2(n_290),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_130),
.A2(n_232),
.B(n_237),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_160),
.B(n_169),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_142),
.A2(n_169),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_142),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_142),
.A2(n_161),
.B1(n_206),
.B2(n_350),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_150),
.B(n_152),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_143),
.B(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_143),
.A2(n_263),
.B1(n_269),
.B2(n_273),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_143),
.A2(n_273),
.B(n_305),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_143),
.A2(n_218),
.B(n_395),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_143),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_143),
.A2(n_307),
.B1(n_401),
.B2(n_413),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_143),
.A2(n_152),
.B(n_305),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.Y(n_143)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_144),
.Y(n_265)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_147),
.Y(n_278)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_149),
.Y(n_333)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_149),
.Y(n_425)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

INVx3_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_158),
.Y(n_415)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_159),
.Y(n_268)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_159),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_161),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_170),
.B(n_193),
.Y(n_237)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx8_ASAP7_75t_L g293 ( 
.A(n_172),
.Y(n_293)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_191),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_190),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_240),
.B(n_481),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.C(n_209),
.Y(n_203)
);

FAx1_ASAP7_75t_SL g358 ( 
.A(n_204),
.B(n_208),
.CI(n_209),
.CON(n_358),
.SN(n_358)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_230),
.C(n_238),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_210),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_222),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_211),
.A2(n_222),
.B1(n_223),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_211),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_218),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_213),
.A2(n_264),
.B(n_330),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_214),
.Y(n_309)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

INVx5_ASAP7_75t_L g421 ( 
.A(n_220),
.Y(n_421)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_226),
.Y(n_453)
);

INVx5_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_228),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_230),
.A2(n_231),
.B1(n_238),
.B2(n_239),
.Y(n_352)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_359),
.B(n_475),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_344),
.C(n_356),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_323),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_243),
.A2(n_477),
.B(n_478),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_311),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_244),
.B(n_311),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_294),
.C(n_303),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_245),
.B(n_343),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_279),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_246),
.B(n_280),
.C(n_286),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_262),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_247),
.B(n_262),
.Y(n_326)
);

OAI32xp33_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_251),
.A3(n_252),
.B1(n_254),
.B2(n_259),
.Y(n_247)
);

INVx4_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_251),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVxp33_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_267),
.Y(n_396)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx6_ASAP7_75t_L g402 ( 
.A(n_276),
.Y(n_402)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_277),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_286),
.Y(n_279)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_287),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_294),
.B(n_303),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.C(n_299),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g325 ( 
.A(n_295),
.B(n_296),
.CI(n_299),
.CON(n_325),
.SN(n_325)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_310),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_310),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_309),
.Y(n_305)
);

INVx3_ASAP7_75t_SL g306 ( 
.A(n_307),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_308),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_312),
.B(n_314),
.C(n_316),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_316),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_322),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_321),
.C(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_342),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_324),
.B(n_342),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.C(n_327),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_325),
.B(n_473),
.Y(n_472)
);

BUFx24_ASAP7_75t_SL g483 ( 
.A(n_325),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_326),
.B(n_327),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_334),
.C(n_336),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_328),
.A2(n_329),
.B1(n_334),
.B2(n_335),
.Y(n_460)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx8_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_336),
.B(n_460),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

A2O1A1O1Ixp25_ASAP7_75t_L g475 ( 
.A1(n_344),
.A2(n_356),
.B(n_476),
.C(n_479),
.D(n_480),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_355),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_345),
.B(n_355),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_346),
.B(n_349),
.C(n_354),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_351),
.B1(n_353),
.B2(n_354),
.Y(n_348)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_349),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_351),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_357),
.B(n_358),
.Y(n_480)
);

BUFx24_ASAP7_75t_SL g485 ( 
.A(n_358),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_470),
.B(n_474),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_361),
.A2(n_455),
.B(n_469),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_429),
.B(n_454),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_363),
.A2(n_397),
.B(n_428),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_382),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_364),
.B(n_382),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_374),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_365),
.B(n_374),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_369),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_376),
.B(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_376),
.B(n_440),
.Y(n_439)
);

OAI21xp33_ASAP7_75t_SL g449 ( 
.A1(n_376),
.A2(n_439),
.B(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_381),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_394),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_385),
.B1(n_386),
.B2(n_393),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_384),
.B(n_393),
.C(n_394),
.Y(n_430)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_386),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_395),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_409),
.B(n_427),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_408),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_399),
.B(n_408),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_400),
.A2(n_404),
.B1(n_405),
.B2(n_406),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_402),
.B(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_410),
.A2(n_419),
.B(n_426),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_411),
.B(n_412),
.Y(n_426)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx4_ASAP7_75t_SL g416 ( 
.A(n_417),
.Y(n_416)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_420),
.B(n_422),
.Y(n_419)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_431),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_447),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_448),
.C(n_451),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_446),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_433),
.B(n_446),
.Y(n_463)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx6_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_451),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_452),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_456),
.B(n_457),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_458),
.A2(n_459),
.B1(n_461),
.B2(n_462),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_464),
.C(n_467),
.Y(n_471)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_463),
.A2(n_464),
.B1(n_467),
.B2(n_468),
.Y(n_462)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_463),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_464),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_472),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_471),
.B(n_472),
.Y(n_474)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);


endmodule