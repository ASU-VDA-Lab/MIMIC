module fake_netlist_6_2357_n_2336 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_521, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_533, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_546, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2336);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_533;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_546;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2336;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2129;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_572;
wire n_813;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2207;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_2073;
wire n_2273;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2193;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_690;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_2178;
wire n_950;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_1139;
wire n_872;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_2069;
wire n_2307;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2204;
wire n_1520;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_1905;
wire n_2016;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_621;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_2083;
wire n_1931;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_2287;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_2318;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_2233;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g549 ( 
.A(n_315),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_31),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_21),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_403),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_381),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_21),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_123),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_384),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_0),
.Y(n_557)
);

INVxp67_ASAP7_75t_SL g558 ( 
.A(n_540),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_404),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_183),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_46),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_427),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_406),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_267),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_220),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_367),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_305),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_140),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_333),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_432),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_101),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_335),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_2),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_537),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_261),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_472),
.Y(n_576)
);

CKINVDCx14_ASAP7_75t_R g577 ( 
.A(n_217),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_441),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_437),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_394),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_18),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_22),
.Y(n_582)
);

BUFx5_ASAP7_75t_L g583 ( 
.A(n_309),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_452),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_489),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_174),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_503),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_155),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_372),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_494),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_239),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_229),
.Y(n_592)
);

CKINVDCx16_ASAP7_75t_R g593 ( 
.A(n_108),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_341),
.Y(n_594)
);

CKINVDCx14_ASAP7_75t_R g595 ( 
.A(n_295),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_224),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_397),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_188),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_52),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_28),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_209),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_7),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_61),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_341),
.Y(n_604)
);

BUFx8_ASAP7_75t_SL g605 ( 
.A(n_490),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_396),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_497),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_322),
.Y(n_608)
);

CKINVDCx16_ASAP7_75t_R g609 ( 
.A(n_473),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_469),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_156),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_51),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_501),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_293),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_376),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_251),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_211),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_519),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_63),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_251),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_4),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_434),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_402),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_356),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_498),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_157),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_122),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_281),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_121),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_228),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_96),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_202),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_529),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_31),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_137),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_148),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_89),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_217),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_99),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_407),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_496),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_315),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_420),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_330),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_121),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_425),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_438),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_75),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_203),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_392),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_412),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_105),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_36),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_495),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_274),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_510),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_479),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_443),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_350),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_46),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_33),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_302),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_7),
.Y(n_663)
);

BUFx5_ASAP7_75t_L g664 ( 
.A(n_29),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_92),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_340),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_321),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_255),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_262),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_263),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_483),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_271),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_199),
.Y(n_673)
);

INVx1_ASAP7_75t_SL g674 ( 
.A(n_373),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_16),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_461),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_182),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_440),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_335),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_542),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_141),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_340),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_465),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_211),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_376),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_39),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_117),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_76),
.Y(n_688)
);

BUFx10_ASAP7_75t_L g689 ( 
.A(n_411),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_331),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_309),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_387),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_53),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_428),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_64),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_319),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_42),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_439),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_200),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_306),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_175),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_395),
.Y(n_702)
);

BUFx5_ASAP7_75t_L g703 ( 
.A(n_522),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_233),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_385),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_38),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_457),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_0),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_525),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_209),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_254),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_163),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_239),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_356),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_324),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_185),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_224),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_347),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_358),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_463),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_386),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_327),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_50),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_297),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_47),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_291),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_347),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_230),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_471),
.Y(n_729)
);

BUFx2_ASAP7_75t_SL g730 ( 
.A(n_81),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_82),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_41),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_231),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_173),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_28),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_189),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_366),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_388),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_108),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_143),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_160),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_77),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_486),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_405),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_442),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_287),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_20),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_366),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_444),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_543),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_349),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_91),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_168),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_6),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_245),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_213),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_448),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_367),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_98),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_125),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_583),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_753),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_583),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_583),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_583),
.Y(n_765)
);

INVxp67_ASAP7_75t_SL g766 ( 
.A(n_694),
.Y(n_766)
);

BUFx10_ASAP7_75t_L g767 ( 
.A(n_628),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_583),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_583),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_583),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_560),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_664),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_664),
.Y(n_773)
);

INVxp33_ASAP7_75t_SL g774 ( 
.A(n_730),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_554),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_689),
.Y(n_776)
);

CKINVDCx16_ASAP7_75t_R g777 ( 
.A(n_593),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_664),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_577),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_664),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_664),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_664),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_664),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_644),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_644),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_644),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_644),
.Y(n_787)
);

INVxp33_ASAP7_75t_L g788 ( 
.A(n_549),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_701),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_701),
.Y(n_790)
);

CKINVDCx14_ASAP7_75t_R g791 ( 
.A(n_577),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_703),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_560),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_604),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_604),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_714),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_714),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_746),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_746),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_701),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_595),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_701),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_554),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_718),
.Y(n_804)
);

INVxp33_ASAP7_75t_SL g805 ( 
.A(n_551),
.Y(n_805)
);

NOR2xp67_ASAP7_75t_L g806 ( 
.A(n_694),
.B(n_1),
.Y(n_806)
);

INVxp33_ASAP7_75t_SL g807 ( 
.A(n_555),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_718),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_718),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_718),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_616),
.Y(n_811)
);

INVxp67_ASAP7_75t_SL g812 ( 
.A(n_694),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_737),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_595),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_737),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_557),
.Y(n_816)
);

INVxp33_ASAP7_75t_L g817 ( 
.A(n_550),
.Y(n_817)
);

INVxp33_ASAP7_75t_L g818 ( 
.A(n_553),
.Y(n_818)
);

INVxp67_ASAP7_75t_SL g819 ( 
.A(n_737),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_737),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_616),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_556),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_566),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_575),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_588),
.Y(n_825)
);

INVxp33_ASAP7_75t_L g826 ( 
.A(n_592),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_596),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_603),
.Y(n_828)
);

INVxp33_ASAP7_75t_L g829 ( 
.A(n_614),
.Y(n_829)
);

CKINVDCx16_ASAP7_75t_R g830 ( 
.A(n_609),
.Y(n_830)
);

INVxp33_ASAP7_75t_SL g831 ( 
.A(n_561),
.Y(n_831)
);

INVxp33_ASAP7_75t_L g832 ( 
.A(n_615),
.Y(n_832)
);

INVxp67_ASAP7_75t_SL g833 ( 
.A(n_562),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_564),
.Y(n_834)
);

INVxp67_ASAP7_75t_SL g835 ( 
.A(n_570),
.Y(n_835)
);

NOR2xp67_ASAP7_75t_L g836 ( 
.A(n_755),
.B(n_1),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_626),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_601),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_601),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_627),
.Y(n_840)
);

CKINVDCx16_ASAP7_75t_R g841 ( 
.A(n_650),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_611),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_565),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_634),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_567),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_635),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_649),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_636),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_637),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_638),
.Y(n_850)
);

INVxp67_ASAP7_75t_SL g851 ( 
.A(n_574),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_568),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_703),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_563),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_703),
.Y(n_855)
);

CKINVDCx16_ASAP7_75t_R g856 ( 
.A(n_650),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_611),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_662),
.Y(n_858)
);

INVx5_ASAP7_75t_L g859 ( 
.A(n_854),
.Y(n_859)
);

INVx4_ASAP7_75t_L g860 ( 
.A(n_854),
.Y(n_860)
);

INVx4_ASAP7_75t_L g861 ( 
.A(n_854),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_762),
.A2(n_749),
.B1(n_654),
.B2(n_671),
.Y(n_862)
);

INVx5_ASAP7_75t_L g863 ( 
.A(n_854),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_854),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_784),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_784),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_785),
.Y(n_867)
);

BUFx8_ASAP7_75t_L g868 ( 
.A(n_776),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_766),
.B(n_641),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_768),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_785),
.Y(n_871)
);

INVx5_ASAP7_75t_L g872 ( 
.A(n_768),
.Y(n_872)
);

BUFx8_ASAP7_75t_L g873 ( 
.A(n_776),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_786),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_786),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_791),
.B(n_662),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_819),
.B(n_607),
.Y(n_877)
);

NOR2xp67_ASAP7_75t_L g878 ( 
.A(n_816),
.B(n_843),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_779),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_787),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_787),
.Y(n_881)
);

INVx5_ASAP7_75t_L g882 ( 
.A(n_769),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_816),
.Y(n_883)
);

INVx6_ASAP7_75t_L g884 ( 
.A(n_767),
.Y(n_884)
);

CKINVDCx11_ASAP7_75t_R g885 ( 
.A(n_771),
.Y(n_885)
);

OA21x2_ASAP7_75t_L g886 ( 
.A1(n_764),
.A2(n_559),
.B(n_552),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_767),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_830),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_812),
.B(n_607),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_789),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_794),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_833),
.B(n_552),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_789),
.Y(n_893)
);

OAI22x1_ASAP7_75t_SL g894 ( 
.A1(n_771),
.A2(n_687),
.B1(n_697),
.B2(n_649),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_790),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_790),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_841),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_800),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_835),
.B(n_851),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_769),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_802),
.Y(n_901)
);

INVx5_ASAP7_75t_L g902 ( 
.A(n_770),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_770),
.Y(n_903)
);

BUFx8_ASAP7_75t_SL g904 ( 
.A(n_793),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_804),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_856),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_808),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_779),
.B(n_559),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_795),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_809),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_761),
.Y(n_911)
);

AND2x6_ASAP7_75t_L g912 ( 
.A(n_764),
.B(n_563),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_843),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_763),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_810),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_801),
.B(n_623),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_813),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_806),
.B(n_623),
.Y(n_918)
);

AND2x6_ASAP7_75t_L g919 ( 
.A(n_778),
.B(n_563),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_815),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_820),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_778),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_845),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_792),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_904),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_922),
.Y(n_926)
);

CKINVDCx20_ASAP7_75t_R g927 ( 
.A(n_885),
.Y(n_927)
);

CKINVDCx16_ASAP7_75t_R g928 ( 
.A(n_862),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_897),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_922),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_911),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_897),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_906),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_906),
.Y(n_934)
);

OAI21x1_ASAP7_75t_L g935 ( 
.A1(n_886),
.A2(n_772),
.B(n_765),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_876),
.B(n_801),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_918),
.B(n_822),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_900),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_888),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_911),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_914),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_888),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_900),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_868),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_908),
.B(n_847),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_918),
.B(n_823),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_868),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_864),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_914),
.Y(n_949)
);

BUFx10_ASAP7_75t_L g950 ( 
.A(n_884),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_864),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_864),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_868),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_918),
.B(n_824),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_864),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_903),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_891),
.Y(n_957)
);

OA21x2_ASAP7_75t_L g958 ( 
.A1(n_892),
.A2(n_773),
.B(n_780),
.Y(n_958)
);

CKINVDCx16_ASAP7_75t_R g959 ( 
.A(n_879),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_873),
.Y(n_960)
);

NAND2xp33_ASAP7_75t_R g961 ( 
.A(n_913),
.B(n_845),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_891),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_903),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_909),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_887),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_913),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_899),
.B(n_877),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_909),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_893),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_893),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_870),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_898),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_873),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_898),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_873),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_864),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_901),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_879),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_886),
.A2(n_889),
.B(n_869),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_859),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_859),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_859),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_870),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_886),
.A2(n_781),
.B(n_780),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_907),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_907),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_915),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_883),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_884),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_859),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_915),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_870),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_884),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_923),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_894),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_878),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_877),
.B(n_825),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_860),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_874),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_894),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_887),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_860),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_899),
.B(n_814),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_865),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_916),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_874),
.Y(n_1006)
);

AND2x2_ASAP7_75t_SL g1007 ( 
.A(n_877),
.B(n_729),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_899),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_865),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_860),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_1007),
.B(n_563),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_SL g1012 ( 
.A1(n_1007),
.A2(n_811),
.B1(n_821),
.B2(n_793),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_972),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_1008),
.B(n_585),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_1008),
.A2(n_651),
.B1(n_671),
.B2(n_654),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_983),
.Y(n_1016)
);

INVx4_ASAP7_75t_L g1017 ( 
.A(n_950),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_938),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_983),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_978),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_974),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_967),
.B(n_585),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_977),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_938),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_943),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_925),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_943),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_983),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_945),
.B(n_805),
.Y(n_1029)
);

INVx4_ASAP7_75t_L g1030 ( 
.A(n_998),
.Y(n_1030)
);

AND3x2_ASAP7_75t_L g1031 ( 
.A(n_1001),
.B(n_803),
.C(n_775),
.Y(n_1031)
);

AND2x6_ASAP7_75t_L g1032 ( 
.A(n_1003),
.B(n_729),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_985),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_936),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_958),
.A2(n_886),
.B1(n_693),
.B2(n_710),
.Y(n_1035)
);

AO21x2_ASAP7_75t_L g1036 ( 
.A1(n_979),
.A2(n_558),
.B(n_576),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_986),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_956),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_987),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_956),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_991),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_948),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_963),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_926),
.B(n_852),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_932),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_969),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1005),
.A2(n_678),
.B1(n_749),
.B2(n_651),
.Y(n_1047)
);

INVxp33_ASAP7_75t_L g1048 ( 
.A(n_937),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_997),
.B(n_585),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_930),
.B(n_852),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_958),
.A2(n_693),
.B1(n_710),
.B2(n_686),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_965),
.B(n_805),
.Y(n_1052)
);

OAI22xp33_ASAP7_75t_SL g1053 ( 
.A1(n_928),
.A2(n_807),
.B1(n_831),
.B2(n_774),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_970),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_996),
.B(n_807),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_997),
.B(n_585),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_1005),
.B(n_831),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_997),
.B(n_834),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_925),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_989),
.B(n_613),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_963),
.Y(n_1061)
);

NAND3xp33_ASAP7_75t_L g1062 ( 
.A(n_961),
.B(n_840),
.C(n_836),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_957),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_984),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_984),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_978),
.Y(n_1066)
);

BUFx10_ASAP7_75t_L g1067 ( 
.A(n_939),
.Y(n_1067)
);

NOR2x1p5_ASAP7_75t_L g1068 ( 
.A(n_989),
.B(n_993),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_962),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_931),
.B(n_865),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_964),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_968),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_940),
.B(n_865),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_999),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_950),
.Y(n_1075)
);

AO21x2_ASAP7_75t_L g1076 ( 
.A1(n_979),
.A2(n_580),
.B(n_579),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_999),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_939),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_950),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1006),
.Y(n_1080)
);

BUFx4f_ASAP7_75t_L g1081 ( 
.A(n_929),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_958),
.A2(n_712),
.B1(n_725),
.B2(n_686),
.Y(n_1082)
);

NOR2x1p5_ASAP7_75t_L g1083 ( 
.A(n_993),
.B(n_796),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_998),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_SL g1085 ( 
.A1(n_995),
.A2(n_821),
.B1(n_811),
.B2(n_687),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_SL g1086 ( 
.A(n_946),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_1006),
.Y(n_1087)
);

OAI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_959),
.A2(n_697),
.B1(n_742),
.B2(n_717),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_948),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_935),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_935),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_954),
.A2(n_725),
.B1(n_728),
.B2(n_712),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_954),
.B(n_613),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_941),
.B(n_865),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_954),
.B(n_613),
.Y(n_1095)
);

INVx6_ASAP7_75t_L g1096 ( 
.A(n_948),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_971),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_988),
.B(n_777),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_949),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_998),
.B(n_613),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_951),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_971),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_992),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_1002),
.B(n_703),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_933),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1002),
.B(n_866),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_951),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_1002),
.Y(n_1108)
);

CKINVDCx6p67_ASAP7_75t_R g1109 ( 
.A(n_927),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_992),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1004),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_948),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_942),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_948),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1010),
.B(n_1009),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_932),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_952),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_952),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_1010),
.B(n_774),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_955),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_976),
.B(n_866),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_942),
.Y(n_1122)
);

NAND3xp33_ASAP7_75t_L g1123 ( 
.A(n_933),
.B(n_798),
.C(n_797),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_976),
.Y(n_1124)
);

INVx4_ASAP7_75t_L g1125 ( 
.A(n_955),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_976),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_955),
.Y(n_1127)
);

OR2x6_ASAP7_75t_L g1128 ( 
.A(n_944),
.B(n_799),
.Y(n_1128)
);

INVx5_ASAP7_75t_L g1129 ( 
.A(n_980),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_955),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_955),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_934),
.A2(n_678),
.B1(n_587),
.B2(n_590),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_980),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_980),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_980),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_980),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_994),
.Y(n_1137)
);

AND2x6_ASAP7_75t_L g1138 ( 
.A(n_981),
.B(n_584),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_1034),
.Y(n_1139)
);

NOR2x1p5_ASAP7_75t_L g1140 ( 
.A(n_1109),
.B(n_944),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1046),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1054),
.Y(n_1142)
);

NOR2xp67_ASAP7_75t_L g1143 ( 
.A(n_1105),
.B(n_947),
.Y(n_1143)
);

OR2x6_ASAP7_75t_L g1144 ( 
.A(n_1113),
.B(n_728),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1058),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_1081),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1119),
.B(n_781),
.Y(n_1147)
);

INVxp33_ASAP7_75t_L g1148 ( 
.A(n_1098),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_1081),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1030),
.B(n_934),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1013),
.Y(n_1151)
);

XNOR2xp5_ASAP7_75t_L g1152 ( 
.A(n_1012),
.B(n_927),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1119),
.B(n_782),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1030),
.B(n_782),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1030),
.B(n_783),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1108),
.B(n_783),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1029),
.B(n_994),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_1072),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1108),
.B(n_880),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1021),
.Y(n_1160)
);

INVxp67_ASAP7_75t_L g1161 ( 
.A(n_1020),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1047),
.B(n_966),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1084),
.B(n_606),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_1066),
.B(n_1015),
.Y(n_1164)
);

NOR2xp67_ASAP7_75t_L g1165 ( 
.A(n_1062),
.B(n_953),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1055),
.B(n_966),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1018),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1075),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1084),
.B(n_702),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1052),
.B(n_767),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1024),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1023),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1055),
.B(n_953),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_L g1174 ( 
.A(n_1052),
.B(n_1000),
.C(n_995),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1051),
.B(n_1082),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1048),
.B(n_960),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1044),
.B(n_1050),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1057),
.B(n_960),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1051),
.B(n_880),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1025),
.Y(n_1180)
);

INVxp67_ASAP7_75t_L g1181 ( 
.A(n_1057),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1033),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1027),
.Y(n_1183)
);

INVxp67_ASAP7_75t_L g1184 ( 
.A(n_1123),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1037),
.Y(n_1185)
);

BUFx5_ASAP7_75t_L g1186 ( 
.A(n_1133),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1082),
.B(n_881),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1016),
.B(n_881),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_1026),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1039),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1016),
.B(n_890),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1019),
.B(n_890),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1132),
.B(n_973),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1041),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1075),
.B(n_973),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1019),
.B(n_1028),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1079),
.B(n_975),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1028),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1092),
.A2(n_742),
.B1(n_717),
.B2(n_731),
.Y(n_1199)
);

NOR2xp67_ASAP7_75t_L g1200 ( 
.A(n_1122),
.B(n_975),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1063),
.B(n_1000),
.Y(n_1201)
);

OR2x6_ASAP7_75t_L g1202 ( 
.A(n_1137),
.B(n_731),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1083),
.B(n_788),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1027),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1099),
.B(n_709),
.Y(n_1205)
);

INVxp33_ASAP7_75t_L g1206 ( 
.A(n_1085),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1079),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1038),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1011),
.B(n_720),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_SL g1210 ( 
.A(n_1026),
.B(n_605),
.Y(n_1210)
);

BUFx4_ASAP7_75t_L g1211 ( 
.A(n_1045),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_SL g1212 ( 
.A(n_1059),
.B(n_605),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1038),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1011),
.B(n_750),
.Y(n_1214)
);

NAND2xp33_ASAP7_75t_L g1215 ( 
.A(n_1032),
.B(n_703),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1017),
.B(n_578),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1069),
.B(n_648),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1067),
.B(n_817),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1040),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1071),
.B(n_895),
.Y(n_1220)
);

INVxp33_ASAP7_75t_L g1221 ( 
.A(n_1014),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1097),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1074),
.B(n_895),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1097),
.Y(n_1224)
);

BUFx2_ASAP7_75t_R g1225 ( 
.A(n_1078),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1078),
.B(n_674),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1074),
.B(n_896),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1017),
.B(n_597),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1092),
.B(n_610),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1067),
.B(n_1068),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1102),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1087),
.B(n_896),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1088),
.B(n_675),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1043),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1077),
.B(n_792),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1045),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1102),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_1116),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1088),
.B(n_759),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_1128),
.Y(n_1240)
);

AO221x1_ASAP7_75t_L g1241 ( 
.A1(n_1101),
.A2(n_668),
.B1(n_681),
.B2(n_663),
.C(n_659),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1014),
.B(n_618),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1103),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1080),
.B(n_853),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1043),
.B(n_853),
.Y(n_1245)
);

INVxp33_ASAP7_75t_L g1246 ( 
.A(n_1116),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1067),
.B(n_818),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1061),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1103),
.Y(n_1249)
);

INVx2_ASAP7_75t_SL g1250 ( 
.A(n_1031),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1060),
.B(n_622),
.Y(n_1251)
);

NAND3xp33_ASAP7_75t_L g1252 ( 
.A(n_1060),
.B(n_571),
.C(n_569),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1061),
.B(n_855),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1053),
.B(n_826),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1086),
.B(n_1059),
.Y(n_1255)
);

INVx2_ASAP7_75t_SL g1256 ( 
.A(n_1128),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1042),
.B(n_625),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1035),
.B(n_855),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1035),
.B(n_866),
.Y(n_1259)
);

INVxp67_ASAP7_75t_L g1260 ( 
.A(n_1128),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1110),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1086),
.B(n_829),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1032),
.B(n_866),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1042),
.B(n_633),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1111),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1117),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1042),
.B(n_640),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1042),
.B(n_643),
.Y(n_1268)
);

NOR3xp33_ASAP7_75t_L g1269 ( 
.A(n_1049),
.B(n_828),
.C(n_827),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1032),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1117),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1049),
.B(n_832),
.Y(n_1272)
);

OR2x6_ASAP7_75t_L g1273 ( 
.A(n_1056),
.B(n_602),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1089),
.B(n_646),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1124),
.Y(n_1275)
);

NAND3xp33_ASAP7_75t_L g1276 ( 
.A(n_1093),
.B(n_573),
.C(n_572),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1064),
.B(n_867),
.Y(n_1277)
);

BUFx8_ASAP7_75t_L g1278 ( 
.A(n_1138),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1093),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1101),
.Y(n_1280)
);

INVx4_ASAP7_75t_L g1281 ( 
.A(n_1089),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1089),
.B(n_647),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1126),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1107),
.Y(n_1284)
);

BUFx5_ASAP7_75t_L g1285 ( 
.A(n_1136),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1089),
.B(n_656),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1112),
.B(n_657),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1118),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1112),
.B(n_658),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1095),
.B(n_581),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1112),
.B(n_676),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1112),
.B(n_680),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1118),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1115),
.B(n_582),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1104),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1104),
.B(n_586),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1022),
.A2(n_691),
.B(n_685),
.C(n_684),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1130),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1065),
.B(n_867),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1076),
.B(n_837),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1130),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1131),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1131),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1076),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1070),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1073),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1094),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1127),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1121),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_1036),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1114),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1100),
.B(n_589),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1100),
.B(n_1106),
.Y(n_1313)
);

NOR3xp33_ASAP7_75t_L g1314 ( 
.A(n_1120),
.B(n_846),
.C(n_844),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1141),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1142),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1151),
.Y(n_1317)
);

OAI221xp5_ASAP7_75t_L g1318 ( 
.A1(n_1233),
.A2(n_598),
.B1(n_599),
.B2(n_594),
.C(n_591),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1181),
.B(n_1114),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1177),
.A2(n_698),
.B1(n_707),
.B2(n_683),
.Y(n_1320)
);

OR2x6_ASAP7_75t_L g1321 ( 
.A(n_1146),
.B(n_1096),
.Y(n_1321)
);

OAI221xp5_ASAP7_75t_L g1322 ( 
.A1(n_1239),
.A2(n_612),
.B1(n_617),
.B2(n_608),
.C(n_600),
.Y(n_1322)
);

AO22x2_ASAP7_75t_L g1323 ( 
.A1(n_1199),
.A2(n_695),
.B1(n_696),
.B2(n_692),
.Y(n_1323)
);

AO22x2_ASAP7_75t_L g1324 ( 
.A1(n_1199),
.A2(n_715),
.B1(n_716),
.B2(n_713),
.Y(n_1324)
);

BUFx8_ASAP7_75t_L g1325 ( 
.A(n_1250),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1160),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1167),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1168),
.B(n_1120),
.Y(n_1328)
);

AO22x1_ASAP7_75t_L g1329 ( 
.A1(n_1206),
.A2(n_620),
.B1(n_621),
.B2(n_619),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1145),
.B(n_848),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1172),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1182),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1185),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_1168),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1296),
.A2(n_743),
.B1(n_745),
.B2(n_744),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1238),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1190),
.Y(n_1337)
);

AO22x2_ASAP7_75t_L g1338 ( 
.A1(n_1164),
.A2(n_733),
.B1(n_734),
.B2(n_724),
.Y(n_1338)
);

OR2x6_ASAP7_75t_L g1339 ( 
.A(n_1149),
.B(n_1096),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1294),
.B(n_1090),
.Y(n_1340)
);

NAND2x1p5_ASAP7_75t_L g1341 ( 
.A(n_1168),
.B(n_1125),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1171),
.Y(n_1342)
);

AO22x2_ASAP7_75t_L g1343 ( 
.A1(n_1304),
.A2(n_739),
.B1(n_740),
.B2(n_735),
.Y(n_1343)
);

AO22x2_ASAP7_75t_L g1344 ( 
.A1(n_1174),
.A2(n_748),
.B1(n_752),
.B2(n_747),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1194),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1189),
.Y(n_1346)
);

NAND2x1_ASAP7_75t_L g1347 ( 
.A(n_1281),
.B(n_1096),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1222),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1224),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1231),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1237),
.Y(n_1351)
);

INVxp33_ASAP7_75t_SL g1352 ( 
.A(n_1157),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1147),
.B(n_1091),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1243),
.Y(n_1354)
);

NAND2x1p5_ASAP7_75t_L g1355 ( 
.A(n_1207),
.B(n_1134),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1249),
.Y(n_1356)
);

NAND2x1p5_ASAP7_75t_L g1357 ( 
.A(n_1207),
.B(n_1134),
.Y(n_1357)
);

NAND2x1p5_ASAP7_75t_L g1358 ( 
.A(n_1281),
.B(n_1135),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1139),
.Y(n_1359)
);

OAI221xp5_ASAP7_75t_L g1360 ( 
.A1(n_1254),
.A2(n_630),
.B1(n_631),
.B2(n_629),
.C(n_624),
.Y(n_1360)
);

CKINVDCx16_ASAP7_75t_R g1361 ( 
.A(n_1210),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1180),
.Y(n_1362)
);

OAI221xp5_ASAP7_75t_L g1363 ( 
.A1(n_1162),
.A2(n_642),
.B1(n_645),
.B2(n_639),
.C(n_632),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1311),
.B(n_1158),
.Y(n_1364)
);

BUFx8_ASAP7_75t_L g1365 ( 
.A(n_1230),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1183),
.Y(n_1366)
);

AO22x2_ASAP7_75t_L g1367 ( 
.A1(n_1170),
.A2(n_756),
.B1(n_758),
.B2(n_754),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1204),
.Y(n_1368)
);

AO22x2_ASAP7_75t_L g1369 ( 
.A1(n_1175),
.A2(n_1236),
.B1(n_1256),
.B2(n_1310),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1265),
.B(n_1135),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1208),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1213),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1225),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1178),
.Y(n_1374)
);

AO22x2_ASAP7_75t_L g1375 ( 
.A1(n_1300),
.A2(n_1036),
.B1(n_850),
.B2(n_849),
.Y(n_1375)
);

CKINVDCx14_ASAP7_75t_R g1376 ( 
.A(n_1152),
.Y(n_1376)
);

BUFx8_ASAP7_75t_L g1377 ( 
.A(n_1218),
.Y(n_1377)
);

AO22x2_ASAP7_75t_L g1378 ( 
.A1(n_1240),
.A2(n_839),
.B1(n_842),
.B2(n_838),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1247),
.B(n_838),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1255),
.Y(n_1380)
);

AO22x2_ASAP7_75t_L g1381 ( 
.A1(n_1260),
.A2(n_842),
.B1(n_857),
.B2(n_839),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1153),
.B(n_757),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1219),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1234),
.Y(n_1384)
);

INVxp67_ASAP7_75t_L g1385 ( 
.A(n_1203),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1248),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1272),
.B(n_857),
.Y(n_1387)
);

OAI221xp5_ASAP7_75t_L g1388 ( 
.A1(n_1184),
.A2(n_655),
.B1(n_660),
.B2(n_653),
.C(n_652),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1261),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1266),
.Y(n_1390)
);

AO22x2_ASAP7_75t_L g1391 ( 
.A1(n_1150),
.A2(n_858),
.B1(n_4),
.B2(n_2),
.Y(n_1391)
);

OAI221xp5_ASAP7_75t_L g1392 ( 
.A1(n_1193),
.A2(n_666),
.B1(n_667),
.B2(n_665),
.C(n_661),
.Y(n_1392)
);

AO22x2_ASAP7_75t_L g1393 ( 
.A1(n_1279),
.A2(n_858),
.B1(n_6),
.B2(n_3),
.Y(n_1393)
);

AO22x2_ASAP7_75t_L g1394 ( 
.A1(n_1176),
.A2(n_8),
.B1(n_3),
.B2(n_5),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1275),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1305),
.B(n_1138),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1271),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1161),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1306),
.B(n_1138),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1217),
.B(n_669),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1220),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1221),
.B(n_689),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1298),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1303),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1307),
.B(n_1138),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1283),
.Y(n_1406)
);

OAI221xp5_ASAP7_75t_L g1407 ( 
.A1(n_1226),
.A2(n_673),
.B1(n_677),
.B2(n_672),
.C(n_670),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1173),
.B(n_679),
.Y(n_1408)
);

AO22x2_ASAP7_75t_L g1409 ( 
.A1(n_1252),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1148),
.B(n_689),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1301),
.Y(n_1411)
);

NAND2x1p5_ASAP7_75t_L g1412 ( 
.A(n_1311),
.B(n_1198),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1166),
.B(n_682),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1302),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1188),
.Y(n_1415)
);

CKINVDCx16_ASAP7_75t_R g1416 ( 
.A(n_1212),
.Y(n_1416)
);

NAND2x1p5_ASAP7_75t_L g1417 ( 
.A(n_1198),
.B(n_1129),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1188),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1202),
.Y(n_1419)
);

NAND2x1p5_ASAP7_75t_L g1420 ( 
.A(n_1200),
.B(n_1129),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1309),
.B(n_688),
.Y(n_1421)
);

AO22x2_ASAP7_75t_L g1422 ( 
.A1(n_1295),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1191),
.Y(n_1423)
);

NAND2x1p5_ASAP7_75t_L g1424 ( 
.A(n_1270),
.B(n_1129),
.Y(n_1424)
);

NAND2x1p5_ASAP7_75t_L g1425 ( 
.A(n_1143),
.B(n_1129),
.Y(n_1425)
);

AO22x2_ASAP7_75t_L g1426 ( 
.A1(n_1195),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1191),
.Y(n_1427)
);

BUFx8_ASAP7_75t_L g1428 ( 
.A(n_1211),
.Y(n_1428)
);

NAND2x1p5_ASAP7_75t_L g1429 ( 
.A(n_1280),
.B(n_861),
.Y(n_1429)
);

OAI221xp5_ASAP7_75t_L g1430 ( 
.A1(n_1201),
.A2(n_700),
.B1(n_704),
.B2(n_699),
.C(n_690),
.Y(n_1430)
);

AO22x2_ASAP7_75t_L g1431 ( 
.A1(n_1197),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1290),
.B(n_705),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1192),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1288),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1192),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1308),
.Y(n_1436)
);

AO22x2_ASAP7_75t_L g1437 ( 
.A1(n_1209),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1312),
.A2(n_919),
.B1(n_912),
.B2(n_910),
.Y(n_1438)
);

NAND2x1p5_ASAP7_75t_L g1439 ( 
.A(n_1284),
.B(n_861),
.Y(n_1439)
);

INVxp67_ASAP7_75t_L g1440 ( 
.A(n_1262),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1144),
.B(n_706),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1293),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1165),
.B(n_389),
.Y(n_1443)
);

OAI221xp5_ASAP7_75t_L g1444 ( 
.A1(n_1202),
.A2(n_1144),
.B1(n_1314),
.B2(n_1269),
.C(n_1229),
.Y(n_1444)
);

AO22x2_ASAP7_75t_L g1445 ( 
.A1(n_1214),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1445)
);

CKINVDCx6p67_ASAP7_75t_R g1446 ( 
.A(n_1202),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1140),
.B(n_390),
.Y(n_1447)
);

NAND2x1p5_ASAP7_75t_L g1448 ( 
.A(n_1196),
.B(n_861),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_1144),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1235),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1278),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1313),
.B(n_708),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1273),
.B(n_711),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1235),
.Y(n_1454)
);

NAND2x1p5_ASAP7_75t_L g1455 ( 
.A(n_1196),
.B(n_1216),
.Y(n_1455)
);

AO22x2_ASAP7_75t_L g1456 ( 
.A1(n_1242),
.A2(n_22),
.B1(n_19),
.B2(n_20),
.Y(n_1456)
);

NAND2x1p5_ASAP7_75t_L g1457 ( 
.A(n_1228),
.B(n_867),
.Y(n_1457)
);

NAND2x1p5_ASAP7_75t_L g1458 ( 
.A(n_1257),
.B(n_871),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1154),
.B(n_719),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1273),
.B(n_391),
.Y(n_1460)
);

NAND2x1p5_ASAP7_75t_L g1461 ( 
.A(n_1264),
.B(n_871),
.Y(n_1461)
);

AO22x2_ASAP7_75t_L g1462 ( 
.A1(n_1251),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1462)
);

NAND2x1p5_ASAP7_75t_L g1463 ( 
.A(n_1267),
.B(n_871),
.Y(n_1463)
);

AO22x2_ASAP7_75t_L g1464 ( 
.A1(n_1259),
.A2(n_1276),
.B1(n_1241),
.B2(n_1187),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1244),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1244),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1245),
.Y(n_1467)
);

AO22x2_ASAP7_75t_L g1468 ( 
.A1(n_1259),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1468)
);

INVxp67_ASAP7_75t_L g1469 ( 
.A(n_1205),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1155),
.B(n_721),
.Y(n_1470)
);

AND2x2_ASAP7_75t_SL g1471 ( 
.A(n_1215),
.B(n_26),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1156),
.B(n_722),
.Y(n_1472)
);

AO22x2_ASAP7_75t_L g1473 ( 
.A1(n_1179),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_L g1474 ( 
.A(n_1273),
.B(n_726),
.C(n_723),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1253),
.Y(n_1475)
);

AND2x6_ASAP7_75t_L g1476 ( 
.A(n_1258),
.B(n_981),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1223),
.Y(n_1477)
);

AOI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1268),
.A2(n_919),
.B1(n_912),
.B2(n_910),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1227),
.Y(n_1479)
);

OAI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1297),
.A2(n_736),
.B1(n_738),
.B2(n_732),
.C(n_727),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1232),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1277),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1274),
.A2(n_919),
.B1(n_912),
.B2(n_910),
.Y(n_1483)
);

BUFx8_ASAP7_75t_L g1484 ( 
.A(n_1246),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1186),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1299),
.Y(n_1486)
);

CKINVDCx10_ASAP7_75t_R g1487 ( 
.A(n_1361),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1352),
.B(n_1163),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1408),
.B(n_1169),
.Y(n_1489)
);

NAND3xp33_ASAP7_75t_L g1490 ( 
.A(n_1432),
.B(n_1286),
.C(n_1282),
.Y(n_1490)
);

OAI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1340),
.A2(n_1187),
.B(n_1179),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1398),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1315),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1353),
.A2(n_1159),
.B(n_1263),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1379),
.B(n_1287),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1334),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1316),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1363),
.A2(n_1291),
.B1(n_1292),
.B2(n_1289),
.Y(n_1498)
);

OR2x6_ASAP7_75t_SL g1499 ( 
.A(n_1346),
.B(n_741),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1387),
.B(n_1186),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1469),
.B(n_1285),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_1334),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1317),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1401),
.B(n_1285),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1400),
.B(n_1413),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1382),
.A2(n_919),
.B(n_912),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1326),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1459),
.B(n_1285),
.Y(n_1508)
);

O2A1O1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1360),
.A2(n_760),
.B(n_751),
.C(n_32),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1470),
.B(n_1285),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1452),
.A2(n_919),
.B(n_912),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1450),
.A2(n_924),
.B(n_863),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1330),
.B(n_1285),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1472),
.B(n_1285),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1385),
.B(n_905),
.Y(n_1515)
);

AO21x1_ASAP7_75t_L g1516 ( 
.A1(n_1455),
.A2(n_27),
.B(n_30),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1328),
.Y(n_1517)
);

OAI321xp33_ASAP7_75t_L g1518 ( 
.A1(n_1318),
.A2(n_33),
.A3(n_35),
.B1(n_30),
.B2(n_32),
.C(n_34),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1454),
.A2(n_924),
.B(n_863),
.Y(n_1519)
);

AOI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1375),
.A2(n_1464),
.B(n_1399),
.Y(n_1520)
);

CKINVDCx8_ASAP7_75t_R g1521 ( 
.A(n_1373),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1415),
.B(n_34),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1418),
.B(n_36),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1423),
.B(n_37),
.Y(n_1524)
);

O2A1O1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1392),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_1525)
);

A2O1A1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1444),
.A2(n_910),
.B(n_917),
.C(n_905),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1465),
.A2(n_882),
.B(n_872),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1336),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1331),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1427),
.B(n_40),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1332),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1440),
.B(n_40),
.Y(n_1532)
);

BUFx12f_ASAP7_75t_L g1533 ( 
.A(n_1428),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1466),
.A2(n_882),
.B(n_872),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1396),
.A2(n_919),
.B(n_912),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1328),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1433),
.B(n_1435),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1467),
.A2(n_882),
.B(n_872),
.Y(n_1538)
);

O2A1O1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1322),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1477),
.B(n_43),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1374),
.A2(n_919),
.B1(n_910),
.B2(n_917),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_SL g1542 ( 
.A(n_1471),
.B(n_44),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1475),
.A2(n_902),
.B(n_882),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1333),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1479),
.B(n_44),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1359),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1482),
.A2(n_875),
.B(n_871),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1336),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1380),
.B(n_905),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1347),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1416),
.B(n_905),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1481),
.B(n_45),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1405),
.A2(n_902),
.B(n_393),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1337),
.Y(n_1554)
);

O2A1O1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1430),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1421),
.B(n_48),
.Y(n_1556)
);

BUFx8_ASAP7_75t_L g1557 ( 
.A(n_1419),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1486),
.A2(n_990),
.B(n_982),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1345),
.B(n_49),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1377),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1389),
.B(n_50),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1449),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1485),
.A2(n_990),
.B(n_982),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1323),
.B(n_51),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1419),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_1428),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1323),
.B(n_52),
.Y(n_1567)
);

NAND2x1p5_ASAP7_75t_L g1568 ( 
.A(n_1347),
.B(n_871),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1377),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1369),
.Y(n_1570)
);

INVx2_ASAP7_75t_SL g1571 ( 
.A(n_1325),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1367),
.B(n_920),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1348),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1441),
.B(n_1370),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1436),
.A2(n_920),
.B1(n_921),
.B2(n_875),
.Y(n_1575)
);

A2O1A1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1335),
.A2(n_920),
.B(n_921),
.C(n_875),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1406),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1457),
.A2(n_982),
.B(n_981),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1349),
.Y(n_1579)
);

A2O1A1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1480),
.A2(n_920),
.B(n_921),
.C(n_875),
.Y(n_1580)
);

O2A1O1Ixp5_ASAP7_75t_L g1581 ( 
.A1(n_1319),
.A2(n_1402),
.B(n_1410),
.C(n_1350),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1458),
.A2(n_1463),
.B(n_1461),
.Y(n_1582)
);

CKINVDCx10_ASAP7_75t_R g1583 ( 
.A(n_1484),
.Y(n_1583)
);

A2O1A1Ixp33_ASAP7_75t_L g1584 ( 
.A1(n_1474),
.A2(n_921),
.B(n_875),
.C(n_55),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1376),
.A2(n_982),
.B1(n_56),
.B2(n_53),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1370),
.B(n_54),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1407),
.B(n_54),
.Y(n_1587)
);

OA21x2_ASAP7_75t_L g1588 ( 
.A1(n_1395),
.A2(n_399),
.B(n_398),
.Y(n_1588)
);

OAI21xp33_ASAP7_75t_L g1589 ( 
.A1(n_1324),
.A2(n_56),
.B(n_57),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1324),
.B(n_57),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1388),
.B(n_1453),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1351),
.B(n_58),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1448),
.A2(n_401),
.B(n_400),
.Y(n_1593)
);

O2A1O1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1442),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1354),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1356),
.B(n_62),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1369),
.B(n_63),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1439),
.A2(n_409),
.B(n_408),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1411),
.Y(n_1599)
);

INVx5_ASAP7_75t_L g1600 ( 
.A(n_1476),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1414),
.A2(n_413),
.B(n_410),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1443),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1434),
.B(n_65),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1460),
.B(n_66),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1329),
.B(n_67),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1341),
.A2(n_415),
.B(n_414),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1327),
.B(n_67),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1438),
.A2(n_417),
.B(n_416),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1460),
.B(n_68),
.Y(n_1609)
);

NAND3xp33_ASAP7_75t_L g1610 ( 
.A(n_1320),
.B(n_68),
.C(n_69),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1358),
.A2(n_1417),
.B(n_1366),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1342),
.B(n_69),
.Y(n_1612)
);

O2A1O1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1443),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1429),
.A2(n_419),
.B(n_418),
.Y(n_1614)
);

NOR2xp67_ASAP7_75t_L g1615 ( 
.A(n_1451),
.B(n_421),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1362),
.A2(n_423),
.B(n_422),
.Y(n_1616)
);

AOI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1368),
.A2(n_1372),
.B(n_1371),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1344),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1446),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1383),
.Y(n_1620)
);

O2A1O1Ixp5_ASAP7_75t_L g1621 ( 
.A1(n_1384),
.A2(n_77),
.B(n_74),
.C(n_76),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1386),
.A2(n_426),
.B(n_424),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1412),
.A2(n_430),
.B(n_429),
.Y(n_1623)
);

AOI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1343),
.A2(n_548),
.B(n_433),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1447),
.B(n_78),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_1365),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1390),
.A2(n_435),
.B(n_431),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1367),
.B(n_78),
.Y(n_1628)
);

NAND3xp33_ASAP7_75t_L g1629 ( 
.A(n_1397),
.B(n_79),
.C(n_80),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1378),
.B(n_79),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1403),
.A2(n_1404),
.B(n_1424),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1355),
.A2(n_1357),
.B(n_1339),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1378),
.B(n_80),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1364),
.B(n_81),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1321),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1381),
.B(n_1344),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1365),
.B(n_1420),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1381),
.B(n_83),
.Y(n_1638)
);

NAND2x1_ASAP7_75t_L g1639 ( 
.A(n_1321),
.B(n_436),
.Y(n_1639)
);

INVx4_ASAP7_75t_L g1640 ( 
.A(n_1425),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1476),
.B(n_445),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1478),
.A2(n_447),
.B(n_446),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1483),
.A2(n_450),
.B(n_449),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1338),
.B(n_84),
.Y(n_1644)
);

O2A1O1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1489),
.A2(n_1338),
.B(n_1409),
.C(n_1426),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1488),
.B(n_1343),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1517),
.B(n_451),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1493),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1591),
.A2(n_1391),
.B1(n_1431),
.B2(n_1426),
.Y(n_1649)
);

INVxp67_ASAP7_75t_L g1650 ( 
.A(n_1492),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1507),
.Y(n_1651)
);

AO21x1_ASAP7_75t_L g1652 ( 
.A1(n_1542),
.A2(n_1468),
.B(n_1473),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1505),
.A2(n_1431),
.B1(n_1394),
.B2(n_1456),
.Y(n_1653)
);

A2O1A1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1509),
.A2(n_1462),
.B(n_1456),
.C(n_1394),
.Y(n_1654)
);

BUFx12f_ASAP7_75t_L g1655 ( 
.A(n_1533),
.Y(n_1655)
);

A2O1A1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1587),
.A2(n_1462),
.B(n_1409),
.C(n_1393),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1542),
.A2(n_1393),
.B1(n_1445),
.B2(n_1437),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1547),
.A2(n_1468),
.B(n_1422),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1495),
.B(n_1437),
.Y(n_1659)
);

OAI21xp33_ASAP7_75t_L g1660 ( 
.A1(n_1556),
.A2(n_1589),
.B(n_1610),
.Y(n_1660)
);

INVx5_ASAP7_75t_L g1661 ( 
.A(n_1496),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1537),
.B(n_1445),
.Y(n_1662)
);

CKINVDCx14_ASAP7_75t_R g1663 ( 
.A(n_1566),
.Y(n_1663)
);

INVx6_ASAP7_75t_L g1664 ( 
.A(n_1557),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1513),
.B(n_85),
.Y(n_1665)
);

INVxp67_ASAP7_75t_SL g1666 ( 
.A(n_1500),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1528),
.B(n_85),
.Y(n_1667)
);

O2A1O1Ixp33_ASAP7_75t_L g1668 ( 
.A1(n_1525),
.A2(n_88),
.B(n_86),
.C(n_87),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1529),
.Y(n_1669)
);

INVx8_ASAP7_75t_L g1670 ( 
.A(n_1496),
.Y(n_1670)
);

AOI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1494),
.A2(n_454),
.B(n_453),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1554),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1501),
.B(n_86),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1508),
.A2(n_547),
.B(n_456),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1562),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1625),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1546),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1510),
.A2(n_458),
.B(n_455),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1546),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1610),
.A2(n_94),
.B1(n_90),
.B2(n_93),
.Y(n_1680)
);

AND2x6_ASAP7_75t_L g1681 ( 
.A(n_1641),
.B(n_459),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_SL g1682 ( 
.A(n_1521),
.B(n_460),
.Y(n_1682)
);

INVx1_ASAP7_75t_SL g1683 ( 
.A(n_1548),
.Y(n_1683)
);

NAND2xp33_ASAP7_75t_L g1684 ( 
.A(n_1517),
.B(n_1562),
.Y(n_1684)
);

O2A1O1Ixp33_ASAP7_75t_L g1685 ( 
.A1(n_1539),
.A2(n_95),
.B(n_93),
.C(n_94),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1574),
.B(n_96),
.Y(n_1686)
);

INVx4_ASAP7_75t_L g1687 ( 
.A(n_1496),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1514),
.A2(n_546),
.B(n_464),
.Y(n_1688)
);

A2O1A1Ixp33_ASAP7_75t_SL g1689 ( 
.A1(n_1518),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1604),
.B(n_462),
.Y(n_1690)
);

BUFx4f_ASAP7_75t_L g1691 ( 
.A(n_1502),
.Y(n_1691)
);

O2A1O1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1555),
.A2(n_101),
.B(n_97),
.C(n_100),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1609),
.B(n_466),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1577),
.B(n_1565),
.Y(n_1694)
);

INVx2_ASAP7_75t_SL g1695 ( 
.A(n_1557),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1540),
.B(n_102),
.Y(n_1696)
);

O2A1O1Ixp33_ASAP7_75t_L g1697 ( 
.A1(n_1644),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_SL g1698 ( 
.A(n_1581),
.B(n_104),
.Y(n_1698)
);

NOR3xp33_ASAP7_75t_L g1699 ( 
.A(n_1605),
.B(n_106),
.C(n_107),
.Y(n_1699)
);

INVx4_ASAP7_75t_L g1700 ( 
.A(n_1502),
.Y(n_1700)
);

INVx4_ASAP7_75t_L g1701 ( 
.A(n_1502),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_SL g1702 ( 
.A1(n_1585),
.A2(n_109),
.B1(n_106),
.B2(n_107),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1497),
.Y(n_1703)
);

A2O1A1Ixp33_ASAP7_75t_L g1704 ( 
.A1(n_1608),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1551),
.B(n_110),
.Y(n_1705)
);

NOR2xp67_ASAP7_75t_SL g1706 ( 
.A(n_1518),
.B(n_111),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1503),
.Y(n_1707)
);

O2A1O1Ixp5_ASAP7_75t_L g1708 ( 
.A1(n_1526),
.A2(n_1608),
.B(n_1520),
.C(n_1516),
.Y(n_1708)
);

OR2x6_ASAP7_75t_L g1709 ( 
.A(n_1560),
.B(n_467),
.Y(n_1709)
);

A2O1A1Ixp33_ASAP7_75t_L g1710 ( 
.A1(n_1490),
.A2(n_114),
.B(n_112),
.C(n_113),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1545),
.B(n_1552),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1602),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1531),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1618),
.B(n_468),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_SL g1715 ( 
.A1(n_1619),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1562),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1544),
.Y(n_1717)
);

OR2x6_ASAP7_75t_L g1718 ( 
.A(n_1571),
.B(n_470),
.Y(n_1718)
);

AOI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1586),
.A2(n_118),
.B1(n_115),
.B2(n_116),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1522),
.B(n_118),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1517),
.B(n_474),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1523),
.B(n_119),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1573),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1626),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1580),
.A2(n_545),
.B(n_476),
.Y(n_1725)
);

XNOR2xp5_ASAP7_75t_L g1726 ( 
.A(n_1569),
.B(n_475),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1498),
.A2(n_1634),
.B1(n_1532),
.B2(n_1549),
.Y(n_1727)
);

INVxp67_ASAP7_75t_SL g1728 ( 
.A(n_1504),
.Y(n_1728)
);

NAND3xp33_ASAP7_75t_L g1729 ( 
.A(n_1613),
.B(n_120),
.C(n_122),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1524),
.B(n_123),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_R g1731 ( 
.A(n_1487),
.B(n_477),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1536),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1491),
.A2(n_480),
.B(n_478),
.Y(n_1733)
);

BUFx6f_ASAP7_75t_L g1734 ( 
.A(n_1536),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_R g1735 ( 
.A(n_1583),
.B(n_481),
.Y(n_1735)
);

BUFx3_ASAP7_75t_L g1736 ( 
.A(n_1515),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1491),
.A2(n_544),
.B(n_484),
.Y(n_1737)
);

NAND2xp33_ASAP7_75t_SL g1738 ( 
.A(n_1637),
.B(n_124),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1530),
.B(n_124),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1576),
.A2(n_485),
.B(n_482),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1600),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1553),
.A2(n_541),
.B(n_488),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1579),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1599),
.Y(n_1744)
);

OR2x6_ASAP7_75t_L g1745 ( 
.A(n_1632),
.B(n_487),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1615),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_1639),
.Y(n_1747)
);

INVx2_ASAP7_75t_SL g1748 ( 
.A(n_1640),
.Y(n_1748)
);

AOI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1636),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1570),
.B(n_1572),
.Y(n_1750)
);

OAI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1584),
.A2(n_130),
.B(n_131),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1620),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1570),
.B(n_1564),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1582),
.A2(n_492),
.B(n_491),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1607),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1617),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1559),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1612),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1640),
.B(n_493),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1561),
.B(n_1592),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1600),
.B(n_132),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1596),
.B(n_133),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1499),
.Y(n_1763)
);

AO21x1_ASAP7_75t_L g1764 ( 
.A1(n_1597),
.A2(n_134),
.B(n_135),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1629),
.A2(n_138),
.B1(n_135),
.B2(n_136),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1603),
.B(n_499),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1629),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1630),
.Y(n_1768)
);

OAI21x1_ASAP7_75t_L g1769 ( 
.A1(n_1558),
.A2(n_502),
.B(n_500),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1567),
.B(n_136),
.Y(n_1770)
);

BUFx6f_ASAP7_75t_L g1771 ( 
.A(n_1641),
.Y(n_1771)
);

O2A1O1Ixp33_ASAP7_75t_L g1772 ( 
.A1(n_1628),
.A2(n_140),
.B(n_138),
.C(n_139),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1590),
.B(n_504),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1633),
.B(n_139),
.Y(n_1774)
);

BUFx2_ASAP7_75t_L g1775 ( 
.A(n_1550),
.Y(n_1775)
);

OAI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1541),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1638),
.B(n_142),
.Y(n_1777)
);

NOR3xp33_ASAP7_75t_SL g1778 ( 
.A(n_1635),
.B(n_1595),
.C(n_1594),
.Y(n_1778)
);

INVxp33_ASAP7_75t_SL g1779 ( 
.A(n_1631),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1614),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1611),
.B(n_144),
.Y(n_1781)
);

AO31x2_ASAP7_75t_L g1782 ( 
.A1(n_1575),
.A2(n_147),
.A3(n_145),
.B(n_146),
.Y(n_1782)
);

XNOR2xp5_ASAP7_75t_L g1783 ( 
.A(n_1623),
.B(n_1606),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1511),
.A2(n_506),
.B(n_505),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1601),
.B(n_1598),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1506),
.A2(n_539),
.B(n_508),
.Y(n_1786)
);

INVxp67_ASAP7_75t_L g1787 ( 
.A(n_1588),
.Y(n_1787)
);

NOR2xp67_ASAP7_75t_L g1788 ( 
.A(n_1783),
.B(n_1593),
.Y(n_1788)
);

O2A1O1Ixp5_ASAP7_75t_SL g1789 ( 
.A1(n_1698),
.A2(n_1535),
.B(n_1621),
.C(n_1624),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1711),
.B(n_1616),
.Y(n_1790)
);

INVx5_ASAP7_75t_L g1791 ( 
.A(n_1681),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1659),
.B(n_1588),
.Y(n_1792)
);

INVxp67_ASAP7_75t_SL g1793 ( 
.A(n_1666),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1703),
.Y(n_1794)
);

NAND2x1_ASAP7_75t_L g1795 ( 
.A(n_1745),
.B(n_1627),
.Y(n_1795)
);

A2O1A1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1660),
.A2(n_1642),
.B(n_1643),
.C(n_1622),
.Y(n_1796)
);

OAI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1708),
.A2(n_1534),
.B(n_1527),
.Y(n_1797)
);

OAI21x1_ASAP7_75t_L g1798 ( 
.A1(n_1769),
.A2(n_1519),
.B(n_1512),
.Y(n_1798)
);

AOI21x1_ASAP7_75t_L g1799 ( 
.A1(n_1740),
.A2(n_1543),
.B(n_1538),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1707),
.Y(n_1800)
);

OAI21x1_ASAP7_75t_L g1801 ( 
.A1(n_1725),
.A2(n_1563),
.B(n_1578),
.Y(n_1801)
);

INVxp67_ASAP7_75t_SL g1802 ( 
.A(n_1694),
.Y(n_1802)
);

INVx5_ASAP7_75t_L g1803 ( 
.A(n_1681),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1727),
.B(n_1760),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1650),
.B(n_507),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1713),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1648),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1758),
.B(n_147),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1677),
.B(n_509),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1717),
.Y(n_1810)
);

O2A1O1Ixp33_ASAP7_75t_L g1811 ( 
.A1(n_1704),
.A2(n_1568),
.B(n_150),
.C(n_148),
.Y(n_1811)
);

CKINVDCx20_ASAP7_75t_R g1812 ( 
.A(n_1663),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1755),
.B(n_1768),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_SL g1814 ( 
.A(n_1706),
.B(n_149),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1785),
.A2(n_512),
.B(n_511),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1662),
.B(n_149),
.Y(n_1816)
);

INVxp67_ASAP7_75t_L g1817 ( 
.A(n_1683),
.Y(n_1817)
);

OAI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1742),
.A2(n_150),
.B(n_151),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1779),
.A2(n_514),
.B(n_513),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1657),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_1820)
);

BUFx3_ASAP7_75t_L g1821 ( 
.A(n_1716),
.Y(n_1821)
);

OA21x2_ASAP7_75t_L g1822 ( 
.A1(n_1787),
.A2(n_152),
.B(n_153),
.Y(n_1822)
);

O2A1O1Ixp33_ASAP7_75t_SL g1823 ( 
.A1(n_1689),
.A2(n_1654),
.B(n_1656),
.C(n_1710),
.Y(n_1823)
);

BUFx3_ASAP7_75t_L g1824 ( 
.A(n_1716),
.Y(n_1824)
);

O2A1O1Ixp5_ASAP7_75t_SL g1825 ( 
.A1(n_1653),
.A2(n_156),
.B(n_154),
.C(n_155),
.Y(n_1825)
);

A2O1A1Ixp33_ASAP7_75t_L g1826 ( 
.A1(n_1645),
.A2(n_158),
.B(n_154),
.C(n_157),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1753),
.B(n_515),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1723),
.Y(n_1828)
);

AOI221xp5_ASAP7_75t_L g1829 ( 
.A1(n_1699),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.C(n_161),
.Y(n_1829)
);

BUFx3_ASAP7_75t_L g1830 ( 
.A(n_1716),
.Y(n_1830)
);

INVx2_ASAP7_75t_SL g1831 ( 
.A(n_1670),
.Y(n_1831)
);

BUFx3_ASAP7_75t_L g1832 ( 
.A(n_1675),
.Y(n_1832)
);

INVx1_ASAP7_75t_SL g1833 ( 
.A(n_1744),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1728),
.A2(n_517),
.B(n_516),
.Y(n_1834)
);

OAI21xp33_ASAP7_75t_L g1835 ( 
.A1(n_1680),
.A2(n_162),
.B(n_164),
.Y(n_1835)
);

OAI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1751),
.A2(n_164),
.B(n_165),
.Y(n_1836)
);

AND2x4_ASAP7_75t_L g1837 ( 
.A(n_1771),
.B(n_518),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1733),
.A2(n_521),
.B(n_520),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1743),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1732),
.Y(n_1840)
);

A2O1A1Ixp33_ASAP7_75t_L g1841 ( 
.A1(n_1668),
.A2(n_167),
.B(n_165),
.C(n_166),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1649),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1774),
.B(n_169),
.Y(n_1843)
);

NAND3xp33_ASAP7_75t_L g1844 ( 
.A(n_1778),
.B(n_169),
.C(n_170),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1655),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1750),
.B(n_1736),
.Y(n_1846)
);

OAI21x1_ASAP7_75t_L g1847 ( 
.A1(n_1671),
.A2(n_524),
.B(n_523),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1777),
.B(n_170),
.Y(n_1848)
);

AOI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1737),
.A2(n_1784),
.B(n_1786),
.Y(n_1849)
);

INVx5_ASAP7_75t_L g1850 ( 
.A(n_1681),
.Y(n_1850)
);

NAND3x1_ASAP7_75t_L g1851 ( 
.A(n_1749),
.B(n_171),
.C(n_172),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1646),
.B(n_172),
.Y(n_1852)
);

BUFx2_ASAP7_75t_L g1853 ( 
.A(n_1661),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1651),
.B(n_173),
.Y(n_1854)
);

AND2x4_ASAP7_75t_L g1855 ( 
.A(n_1771),
.B(n_526),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1752),
.Y(n_1856)
);

OAI21x1_ASAP7_75t_SL g1857 ( 
.A1(n_1652),
.A2(n_174),
.B(n_175),
.Y(n_1857)
);

OAI21x1_ASAP7_75t_L g1858 ( 
.A1(n_1756),
.A2(n_528),
.B(n_527),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1669),
.B(n_176),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1702),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_L g1861 ( 
.A(n_1773),
.B(n_530),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1745),
.A2(n_532),
.B(n_531),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1714),
.B(n_533),
.Y(n_1863)
);

OAI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1767),
.A2(n_177),
.B(n_178),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1672),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1686),
.B(n_534),
.Y(n_1866)
);

O2A1O1Ixp5_ASAP7_75t_SL g1867 ( 
.A1(n_1781),
.A2(n_181),
.B(n_179),
.C(n_180),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1734),
.Y(n_1868)
);

BUFx2_ASAP7_75t_L g1869 ( 
.A(n_1661),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1685),
.A2(n_180),
.B(n_181),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1782),
.Y(n_1871)
);

INVx3_ASAP7_75t_SL g1872 ( 
.A(n_1664),
.Y(n_1872)
);

AOI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1754),
.A2(n_536),
.B(n_535),
.Y(n_1873)
);

OAI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1712),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_1874)
);

NOR3xp33_ASAP7_75t_L g1875 ( 
.A(n_1692),
.B(n_184),
.C(n_185),
.Y(n_1875)
);

NAND3x1_ASAP7_75t_L g1876 ( 
.A(n_1770),
.B(n_186),
.C(n_187),
.Y(n_1876)
);

AOI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1674),
.A2(n_538),
.B(n_186),
.Y(n_1877)
);

OAI21x1_ASAP7_75t_L g1878 ( 
.A1(n_1658),
.A2(n_187),
.B(n_188),
.Y(n_1878)
);

A2O1A1Ixp33_ASAP7_75t_L g1879 ( 
.A1(n_1690),
.A2(n_191),
.B(n_189),
.C(n_190),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1678),
.A2(n_190),
.B(n_191),
.Y(n_1880)
);

AOI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1688),
.A2(n_192),
.B(n_193),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1802),
.B(n_1673),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1856),
.Y(n_1883)
);

A2O1A1Ixp33_ASAP7_75t_L g1884 ( 
.A1(n_1836),
.A2(n_1697),
.B(n_1693),
.C(n_1729),
.Y(n_1884)
);

BUFx10_ASAP7_75t_L g1885 ( 
.A(n_1837),
.Y(n_1885)
);

INVx1_ASAP7_75t_SL g1886 ( 
.A(n_1833),
.Y(n_1886)
);

OA21x2_ASAP7_75t_L g1887 ( 
.A1(n_1797),
.A2(n_1764),
.B(n_1765),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1840),
.Y(n_1888)
);

AOI21x1_ASAP7_75t_L g1889 ( 
.A1(n_1795),
.A2(n_1665),
.B(n_1761),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1849),
.A2(n_1684),
.B(n_1766),
.Y(n_1890)
);

OAI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1818),
.A2(n_1772),
.B(n_1746),
.Y(n_1891)
);

INVx2_ASAP7_75t_SL g1892 ( 
.A(n_1794),
.Y(n_1892)
);

OAI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1818),
.A2(n_1757),
.B(n_1676),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1792),
.B(n_1782),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1860),
.A2(n_1715),
.B1(n_1719),
.B2(n_1696),
.Y(n_1895)
);

AND2x4_ASAP7_75t_SL g1896 ( 
.A(n_1846),
.B(n_1771),
.Y(n_1896)
);

BUFx2_ASAP7_75t_L g1897 ( 
.A(n_1793),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_SL g1898 ( 
.A1(n_1836),
.A2(n_1682),
.B1(n_1681),
.B2(n_1776),
.Y(n_1898)
);

AND2x4_ASAP7_75t_L g1899 ( 
.A(n_1791),
.B(n_1775),
.Y(n_1899)
);

OAI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1880),
.A2(n_1722),
.B(n_1720),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1800),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_L g1902 ( 
.A1(n_1875),
.A2(n_1738),
.B1(n_1679),
.B2(n_1741),
.Y(n_1902)
);

BUFx2_ASAP7_75t_L g1903 ( 
.A(n_1871),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_SL g1904 ( 
.A1(n_1842),
.A2(n_1763),
.B1(n_1726),
.B2(n_1695),
.Y(n_1904)
);

AO21x2_ASAP7_75t_L g1905 ( 
.A1(n_1797),
.A2(n_1739),
.B(n_1762),
.Y(n_1905)
);

NAND2x1p5_ASAP7_75t_L g1906 ( 
.A(n_1791),
.B(n_1780),
.Y(n_1906)
);

OAI21x1_ASAP7_75t_L g1907 ( 
.A1(n_1798),
.A2(n_1705),
.B(n_1730),
.Y(n_1907)
);

OAI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1881),
.A2(n_1759),
.B(n_1721),
.Y(n_1908)
);

OAI21x1_ASAP7_75t_L g1909 ( 
.A1(n_1801),
.A2(n_1667),
.B(n_1747),
.Y(n_1909)
);

INVx2_ASAP7_75t_SL g1910 ( 
.A(n_1806),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1810),
.B(n_1734),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1828),
.B(n_1734),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1839),
.Y(n_1913)
);

OAI21x1_ASAP7_75t_L g1914 ( 
.A1(n_1799),
.A2(n_1747),
.B(n_1721),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1865),
.Y(n_1915)
);

NAND2xp33_ASAP7_75t_L g1916 ( 
.A(n_1791),
.B(n_1731),
.Y(n_1916)
);

AOI22x1_ASAP7_75t_L g1917 ( 
.A1(n_1864),
.A2(n_1759),
.B1(n_1748),
.B2(n_1647),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1813),
.Y(n_1918)
);

OAI21x1_ASAP7_75t_L g1919 ( 
.A1(n_1847),
.A2(n_1647),
.B(n_1661),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_1812),
.Y(n_1920)
);

NOR2xp67_ASAP7_75t_L g1921 ( 
.A(n_1803),
.B(n_1724),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1807),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1845),
.Y(n_1923)
);

OAI21x1_ASAP7_75t_L g1924 ( 
.A1(n_1789),
.A2(n_1664),
.B(n_1709),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1822),
.Y(n_1925)
);

AND2x4_ASAP7_75t_L g1926 ( 
.A(n_1803),
.B(n_1687),
.Y(n_1926)
);

OAI21x1_ASAP7_75t_L g1927 ( 
.A1(n_1858),
.A2(n_1709),
.B(n_1670),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1803),
.B(n_1850),
.Y(n_1928)
);

AOI22xp33_ASAP7_75t_L g1929 ( 
.A1(n_1835),
.A2(n_1718),
.B1(n_1724),
.B2(n_1735),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1822),
.Y(n_1930)
);

OAI21x1_ASAP7_75t_L g1931 ( 
.A1(n_1878),
.A2(n_1718),
.B(n_1691),
.Y(n_1931)
);

NAND2x1p5_ASAP7_75t_L g1932 ( 
.A(n_1850),
.B(n_1700),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1850),
.B(n_1701),
.Y(n_1933)
);

INVx2_ASAP7_75t_SL g1934 ( 
.A(n_1892),
.Y(n_1934)
);

OAI21x1_ASAP7_75t_SL g1935 ( 
.A1(n_1891),
.A2(n_1870),
.B(n_1864),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1913),
.Y(n_1936)
);

BUFx2_ASAP7_75t_L g1937 ( 
.A(n_1897),
.Y(n_1937)
);

AOI22xp33_ASAP7_75t_L g1938 ( 
.A1(n_1898),
.A2(n_1835),
.B1(n_1804),
.B2(n_1870),
.Y(n_1938)
);

OR2x2_ASAP7_75t_SL g1939 ( 
.A(n_1887),
.B(n_1844),
.Y(n_1939)
);

INVx6_ASAP7_75t_L g1940 ( 
.A(n_1928),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1890),
.A2(n_1838),
.B(n_1796),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1922),
.Y(n_1942)
);

BUFx12f_ASAP7_75t_L g1943 ( 
.A(n_1923),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1901),
.Y(n_1944)
);

BUFx12f_ASAP7_75t_L g1945 ( 
.A(n_1923),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1915),
.Y(n_1946)
);

CKINVDCx11_ASAP7_75t_R g1947 ( 
.A(n_1886),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_SL g1948 ( 
.A1(n_1893),
.A2(n_1814),
.B1(n_1844),
.B2(n_1861),
.Y(n_1948)
);

BUFx8_ASAP7_75t_L g1949 ( 
.A(n_1928),
.Y(n_1949)
);

AOI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1895),
.A2(n_1788),
.B1(n_1860),
.B2(n_1829),
.Y(n_1950)
);

BUFx3_ASAP7_75t_L g1951 ( 
.A(n_1928),
.Y(n_1951)
);

HB1xp67_ASAP7_75t_L g1952 ( 
.A(n_1897),
.Y(n_1952)
);

NAND2x1p5_ASAP7_75t_L g1953 ( 
.A(n_1914),
.B(n_1833),
.Y(n_1953)
);

AOI22xp33_ASAP7_75t_L g1954 ( 
.A1(n_1917),
.A2(n_1788),
.B1(n_1814),
.B2(n_1874),
.Y(n_1954)
);

BUFx8_ASAP7_75t_L g1955 ( 
.A(n_1926),
.Y(n_1955)
);

CKINVDCx6p67_ASAP7_75t_R g1956 ( 
.A(n_1933),
.Y(n_1956)
);

OAI22xp33_ASAP7_75t_L g1957 ( 
.A1(n_1908),
.A2(n_1820),
.B1(n_1862),
.B2(n_1819),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1918),
.B(n_1790),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1892),
.Y(n_1959)
);

NAND2x1p5_ASAP7_75t_L g1960 ( 
.A(n_1914),
.B(n_1853),
.Y(n_1960)
);

HB1xp67_ASAP7_75t_L g1961 ( 
.A(n_1888),
.Y(n_1961)
);

BUFx2_ASAP7_75t_R g1962 ( 
.A(n_1920),
.Y(n_1962)
);

BUFx2_ASAP7_75t_L g1963 ( 
.A(n_1903),
.Y(n_1963)
);

INVx1_ASAP7_75t_SL g1964 ( 
.A(n_1896),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1902),
.A2(n_1877),
.B1(n_1857),
.B2(n_1863),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1936),
.Y(n_1966)
);

AOI22xp33_ASAP7_75t_L g1967 ( 
.A1(n_1935),
.A2(n_1900),
.B1(n_1887),
.B2(n_1905),
.Y(n_1967)
);

AOI22xp33_ASAP7_75t_L g1968 ( 
.A1(n_1935),
.A2(n_1887),
.B1(n_1905),
.B2(n_1929),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1958),
.B(n_1905),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1961),
.B(n_1883),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_SL g1971 ( 
.A1(n_1938),
.A2(n_1884),
.B(n_1879),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1948),
.A2(n_1950),
.B1(n_1957),
.B2(n_1954),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1941),
.A2(n_1894),
.B1(n_1916),
.B2(n_1873),
.Y(n_1973)
);

AOI22xp33_ASAP7_75t_L g1974 ( 
.A1(n_1965),
.A2(n_1894),
.B1(n_1916),
.B2(n_1924),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1952),
.B(n_1903),
.Y(n_1975)
);

AOI22xp33_ASAP7_75t_L g1976 ( 
.A1(n_1947),
.A2(n_1843),
.B1(n_1848),
.B2(n_1816),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1940),
.Y(n_1977)
);

CKINVDCx20_ASAP7_75t_R g1978 ( 
.A(n_1943),
.Y(n_1978)
);

AOI21xp5_ASAP7_75t_L g1979 ( 
.A1(n_1953),
.A2(n_1823),
.B(n_1811),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1939),
.A2(n_1826),
.B1(n_1851),
.B2(n_1841),
.Y(n_1980)
);

AOI222xp33_ASAP7_75t_L g1981 ( 
.A1(n_1939),
.A2(n_1852),
.B1(n_1882),
.B2(n_1817),
.C1(n_1866),
.C2(n_1809),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1951),
.B(n_1910),
.Y(n_1982)
);

AOI22xp33_ASAP7_75t_L g1983 ( 
.A1(n_1943),
.A2(n_1827),
.B1(n_1805),
.B2(n_1808),
.Y(n_1983)
);

AOI22xp33_ASAP7_75t_SL g1984 ( 
.A1(n_1949),
.A2(n_1904),
.B1(n_1924),
.B2(n_1885),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1942),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1949),
.A2(n_1815),
.B1(n_1907),
.B2(n_1834),
.Y(n_1986)
);

INVxp33_ASAP7_75t_SL g1987 ( 
.A(n_1976),
.Y(n_1987)
);

BUFx6f_ASAP7_75t_L g1988 ( 
.A(n_1977),
.Y(n_1988)
);

OR2x4_ASAP7_75t_L g1989 ( 
.A(n_1971),
.B(n_1962),
.Y(n_1989)
);

BUFx3_ASAP7_75t_L g1990 ( 
.A(n_1978),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1966),
.Y(n_1991)
);

AND2x4_ASAP7_75t_L g1992 ( 
.A(n_1977),
.B(n_1951),
.Y(n_1992)
);

BUFx10_ASAP7_75t_L g1993 ( 
.A(n_1979),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_1969),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1985),
.B(n_1963),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1967),
.B(n_1944),
.Y(n_1996)
);

INVx2_ASAP7_75t_SL g1997 ( 
.A(n_1990),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1988),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1992),
.B(n_1951),
.Y(n_1999)
);

AOI221xp5_ASAP7_75t_L g2000 ( 
.A1(n_1987),
.A2(n_1972),
.B1(n_1980),
.B2(n_1967),
.C(n_1968),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1992),
.B(n_1982),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1996),
.B(n_1981),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_2000),
.B(n_1994),
.Y(n_2003)
);

BUFx2_ASAP7_75t_L g2004 ( 
.A(n_1997),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1999),
.B(n_1993),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_2002),
.B(n_1993),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1998),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_2002),
.Y(n_2008)
);

OAI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1999),
.A2(n_1989),
.B1(n_1974),
.B2(n_1968),
.Y(n_2009)
);

OR2x2_ASAP7_75t_L g2010 ( 
.A(n_2001),
.B(n_1996),
.Y(n_2010)
);

BUFx3_ASAP7_75t_L g2011 ( 
.A(n_1997),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1999),
.B(n_1993),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_2004),
.B(n_1993),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_2010),
.B(n_1970),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_2007),
.Y(n_2015)
);

INVx2_ASAP7_75t_SL g2016 ( 
.A(n_2005),
.Y(n_2016)
);

HB1xp67_ASAP7_75t_L g2017 ( 
.A(n_2011),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_2008),
.B(n_1990),
.Y(n_2018)
);

AND2x4_ASAP7_75t_L g2019 ( 
.A(n_2011),
.B(n_1990),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_2006),
.B(n_1976),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_2005),
.B(n_1992),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2007),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_2012),
.B(n_1992),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_2018),
.B(n_2010),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_2019),
.B(n_2017),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_2014),
.B(n_2003),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_2019),
.B(n_2012),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_2015),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_2019),
.B(n_2009),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_2016),
.B(n_1920),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_2022),
.B(n_1991),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2016),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_2025),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2032),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_2027),
.B(n_2029),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_2030),
.Y(n_2036)
);

AOI31xp33_ASAP7_75t_L g2037 ( 
.A1(n_2033),
.A2(n_2030),
.A3(n_2026),
.B(n_2024),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_2035),
.B(n_2036),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_2034),
.B(n_2021),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_2034),
.B(n_2020),
.Y(n_2040)
);

OAI21xp5_ASAP7_75t_SL g2041 ( 
.A1(n_2037),
.A2(n_2013),
.B(n_2028),
.Y(n_2041)
);

O2A1O1Ixp33_ASAP7_75t_L g2042 ( 
.A1(n_2040),
.A2(n_2013),
.B(n_2031),
.C(n_1872),
.Y(n_2042)
);

O2A1O1Ixp33_ASAP7_75t_L g2043 ( 
.A1(n_2038),
.A2(n_2031),
.B(n_2023),
.C(n_2021),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2039),
.Y(n_2044)
);

AOI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_2038),
.A2(n_2023),
.B1(n_1989),
.B2(n_1984),
.Y(n_2045)
);

AOI21xp33_ASAP7_75t_L g2046 ( 
.A1(n_2037),
.A2(n_1945),
.B(n_1943),
.Y(n_2046)
);

AOI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_2045),
.A2(n_1989),
.B1(n_1945),
.B2(n_1988),
.Y(n_2047)
);

AOI22xp5_ASAP7_75t_L g2048 ( 
.A1(n_2044),
.A2(n_1945),
.B1(n_1988),
.B2(n_1876),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_2041),
.B(n_1988),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_2046),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_2043),
.B(n_1988),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2042),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2044),
.B(n_1991),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2044),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2044),
.Y(n_2055)
);

OAI222xp33_ASAP7_75t_L g2056 ( 
.A1(n_2045),
.A2(n_1983),
.B1(n_1973),
.B2(n_1960),
.C1(n_1953),
.C2(n_1986),
.Y(n_2056)
);

AOI21xp5_ASAP7_75t_L g2057 ( 
.A1(n_2049),
.A2(n_1724),
.B(n_1854),
.Y(n_2057)
);

AOI21xp33_ASAP7_75t_SL g2058 ( 
.A1(n_2054),
.A2(n_192),
.B(n_193),
.Y(n_2058)
);

OR2x2_ASAP7_75t_L g2059 ( 
.A(n_2055),
.B(n_1988),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_2051),
.B(n_1995),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_2050),
.B(n_1995),
.Y(n_2061)
);

OAI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_2047),
.A2(n_1921),
.B1(n_1956),
.B2(n_1932),
.Y(n_2062)
);

AOI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_2052),
.A2(n_1983),
.B1(n_1956),
.B2(n_1940),
.Y(n_2063)
);

AOI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_2048),
.A2(n_1940),
.B1(n_1831),
.B2(n_1995),
.Y(n_2064)
);

OAI32xp33_ASAP7_75t_L g2065 ( 
.A1(n_2053),
.A2(n_1960),
.A3(n_1953),
.B1(n_1975),
.B2(n_1859),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_2053),
.Y(n_2066)
);

AOI21xp33_ASAP7_75t_SL g2067 ( 
.A1(n_2056),
.A2(n_194),
.B(n_195),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2054),
.Y(n_2068)
);

AO22x1_ASAP7_75t_L g2069 ( 
.A1(n_2054),
.A2(n_1837),
.B1(n_1855),
.B2(n_1955),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2059),
.Y(n_2070)
);

NOR3x1_ASAP7_75t_L g2071 ( 
.A(n_2061),
.B(n_1869),
.C(n_1937),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_SL g2072 ( 
.A(n_2067),
.B(n_1832),
.Y(n_2072)
);

OAI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_2063),
.A2(n_1940),
.B1(n_1960),
.B2(n_1932),
.Y(n_2073)
);

OAI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_2057),
.A2(n_1825),
.B(n_1867),
.Y(n_2074)
);

OAI21xp33_ASAP7_75t_L g2075 ( 
.A1(n_2064),
.A2(n_1824),
.B(n_1821),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_2058),
.B(n_194),
.Y(n_2076)
);

NOR2xp33_ASAP7_75t_SL g2077 ( 
.A(n_2068),
.B(n_1855),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_2060),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2066),
.B(n_1944),
.Y(n_2079)
);

AOI21xp5_ASAP7_75t_L g2080 ( 
.A1(n_2062),
.A2(n_1907),
.B(n_1926),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2069),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_2065),
.Y(n_2082)
);

NAND3xp33_ASAP7_75t_SL g2083 ( 
.A(n_2067),
.B(n_1932),
.C(n_1964),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_2060),
.B(n_1937),
.Y(n_2084)
);

NAND3xp33_ASAP7_75t_L g2085 ( 
.A(n_2081),
.B(n_195),
.C(n_196),
.Y(n_2085)
);

AOI221x1_ASAP7_75t_L g2086 ( 
.A1(n_2070),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.C(n_199),
.Y(n_2086)
);

AOI221x1_ASAP7_75t_L g2087 ( 
.A1(n_2076),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.C(n_201),
.Y(n_2087)
);

AOI221xp5_ASAP7_75t_L g2088 ( 
.A1(n_2083),
.A2(n_1830),
.B1(n_1930),
.B2(n_1925),
.C(n_204),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_2077),
.B(n_1926),
.Y(n_2089)
);

NOR4xp25_ASAP7_75t_L g2090 ( 
.A(n_2078),
.B(n_203),
.C(n_201),
.D(n_202),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2082),
.B(n_1946),
.Y(n_2091)
);

NOR2xp33_ASAP7_75t_L g2092 ( 
.A(n_2072),
.B(n_204),
.Y(n_2092)
);

NOR2xp67_ASAP7_75t_SL g2093 ( 
.A(n_2084),
.B(n_205),
.Y(n_2093)
);

OAI222xp33_ASAP7_75t_L g2094 ( 
.A1(n_2073),
.A2(n_1963),
.B1(n_1934),
.B2(n_1889),
.C1(n_1906),
.C2(n_1959),
.Y(n_2094)
);

OAI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_2075),
.A2(n_1933),
.B1(n_1934),
.B2(n_1959),
.Y(n_2095)
);

AOI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_2077),
.A2(n_1933),
.B1(n_1949),
.B2(n_1955),
.Y(n_2096)
);

OAI21xp5_ASAP7_75t_L g2097 ( 
.A1(n_2079),
.A2(n_1931),
.B(n_1927),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_2071),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2093),
.Y(n_2099)
);

NAND4xp25_ASAP7_75t_L g2100 ( 
.A(n_2085),
.B(n_2080),
.C(n_2074),
.D(n_207),
.Y(n_2100)
);

A2O1A1Ixp33_ASAP7_75t_L g2101 ( 
.A1(n_2092),
.A2(n_1931),
.B(n_207),
.C(n_205),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2090),
.B(n_206),
.Y(n_2102)
);

NAND3xp33_ASAP7_75t_L g2103 ( 
.A(n_2087),
.B(n_206),
.C(n_208),
.Y(n_2103)
);

NAND3xp33_ASAP7_75t_SL g2104 ( 
.A(n_2098),
.B(n_2088),
.C(n_2091),
.Y(n_2104)
);

OAI221xp5_ASAP7_75t_L g2105 ( 
.A1(n_2096),
.A2(n_2089),
.B1(n_2097),
.B2(n_2095),
.C(n_2086),
.Y(n_2105)
);

NAND3xp33_ASAP7_75t_L g2106 ( 
.A(n_2094),
.B(n_208),
.C(n_210),
.Y(n_2106)
);

NAND3xp33_ASAP7_75t_SL g2107 ( 
.A(n_2090),
.B(n_210),
.C(n_212),
.Y(n_2107)
);

OAI31xp33_ASAP7_75t_L g2108 ( 
.A1(n_2085),
.A2(n_1906),
.A3(n_214),
.B(n_212),
.Y(n_2108)
);

AOI221xp5_ASAP7_75t_L g2109 ( 
.A1(n_2085),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.C(n_216),
.Y(n_2109)
);

AOI211xp5_ASAP7_75t_L g2110 ( 
.A1(n_2085),
.A2(n_218),
.B(n_215),
.C(n_216),
.Y(n_2110)
);

AOI221xp5_ASAP7_75t_L g2111 ( 
.A1(n_2085),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.C(n_221),
.Y(n_2111)
);

NOR2x1_ASAP7_75t_L g2112 ( 
.A(n_2085),
.B(n_219),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2093),
.Y(n_2113)
);

AOI221xp5_ASAP7_75t_L g2114 ( 
.A1(n_2085),
.A2(n_222),
.B1(n_223),
.B2(n_225),
.C(n_226),
.Y(n_2114)
);

AOI222xp33_ASAP7_75t_L g2115 ( 
.A1(n_2089),
.A2(n_222),
.B1(n_223),
.B2(n_225),
.C1(n_226),
.C2(n_227),
.Y(n_2115)
);

INVx1_ASAP7_75t_SL g2116 ( 
.A(n_2098),
.Y(n_2116)
);

NAND3xp33_ASAP7_75t_L g2117 ( 
.A(n_2093),
.B(n_227),
.C(n_228),
.Y(n_2117)
);

NOR2xp33_ASAP7_75t_SL g2118 ( 
.A(n_2093),
.B(n_1955),
.Y(n_2118)
);

OAI21xp5_ASAP7_75t_L g2119 ( 
.A1(n_2085),
.A2(n_1927),
.B(n_1909),
.Y(n_2119)
);

NAND4xp25_ASAP7_75t_L g2120 ( 
.A(n_2118),
.B(n_2116),
.C(n_2108),
.D(n_2103),
.Y(n_2120)
);

AOI211xp5_ASAP7_75t_L g2121 ( 
.A1(n_2107),
.A2(n_229),
.B(n_230),
.C(n_231),
.Y(n_2121)
);

O2A1O1Ixp33_ASAP7_75t_L g2122 ( 
.A1(n_2102),
.A2(n_232),
.B(n_233),
.C(n_234),
.Y(n_2122)
);

A2O1A1O1Ixp25_ASAP7_75t_L g2123 ( 
.A1(n_2105),
.A2(n_232),
.B(n_234),
.C(n_235),
.D(n_236),
.Y(n_2123)
);

HB1xp67_ASAP7_75t_L g2124 ( 
.A(n_2099),
.Y(n_2124)
);

AOI311xp33_ASAP7_75t_L g2125 ( 
.A1(n_2113),
.A2(n_235),
.A3(n_236),
.B(n_237),
.C(n_238),
.Y(n_2125)
);

AOI222xp33_ASAP7_75t_L g2126 ( 
.A1(n_2104),
.A2(n_237),
.B1(n_238),
.B2(n_240),
.C1(n_241),
.C2(n_242),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2115),
.B(n_240),
.Y(n_2127)
);

NOR3xp33_ASAP7_75t_L g2128 ( 
.A(n_2117),
.B(n_241),
.C(n_242),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_2109),
.B(n_2111),
.Y(n_2129)
);

NAND4xp25_ASAP7_75t_SL g2130 ( 
.A(n_2106),
.B(n_243),
.C(n_244),
.D(n_245),
.Y(n_2130)
);

AOI221xp5_ASAP7_75t_L g2131 ( 
.A1(n_2100),
.A2(n_243),
.B1(n_244),
.B2(n_246),
.C(n_247),
.Y(n_2131)
);

A2O1A1Ixp33_ASAP7_75t_L g2132 ( 
.A1(n_2114),
.A2(n_2110),
.B(n_2101),
.C(n_2112),
.Y(n_2132)
);

NOR2x1_ASAP7_75t_L g2133 ( 
.A(n_2119),
.B(n_246),
.Y(n_2133)
);

AOI221x1_ASAP7_75t_L g2134 ( 
.A1(n_2099),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.C(n_250),
.Y(n_2134)
);

AOI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2118),
.A2(n_1949),
.B1(n_1955),
.B2(n_1868),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2099),
.B(n_1896),
.Y(n_2136)
);

AOI221xp5_ASAP7_75t_L g2137 ( 
.A1(n_2105),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.C(n_252),
.Y(n_2137)
);

NAND4xp25_ASAP7_75t_L g2138 ( 
.A(n_2118),
.B(n_252),
.C(n_253),
.D(n_254),
.Y(n_2138)
);

OAI211xp5_ASAP7_75t_SL g2139 ( 
.A1(n_2099),
.A2(n_253),
.B(n_255),
.C(n_256),
.Y(n_2139)
);

OAI31xp33_ASAP7_75t_L g2140 ( 
.A1(n_2103),
.A2(n_1906),
.A3(n_257),
.B(n_258),
.Y(n_2140)
);

OAI21xp33_ASAP7_75t_SL g2141 ( 
.A1(n_2108),
.A2(n_1919),
.B(n_1909),
.Y(n_2141)
);

AOI221xp5_ASAP7_75t_L g2142 ( 
.A1(n_2105),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.C(n_259),
.Y(n_2142)
);

NOR2xp33_ASAP7_75t_R g2143 ( 
.A(n_2107),
.B(n_259),
.Y(n_2143)
);

AOI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_2118),
.A2(n_1899),
.B1(n_1911),
.B2(n_1912),
.Y(n_2144)
);

AOI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_2118),
.A2(n_260),
.B(n_261),
.Y(n_2145)
);

AOI221xp5_ASAP7_75t_SL g2146 ( 
.A1(n_2116),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.C(n_264),
.Y(n_2146)
);

OAI221xp5_ASAP7_75t_L g2147 ( 
.A1(n_2118),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.C(n_267),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2102),
.Y(n_2148)
);

AOI222xp33_ASAP7_75t_L g2149 ( 
.A1(n_2107),
.A2(n_265),
.B1(n_266),
.B2(n_268),
.C1(n_269),
.C2(n_270),
.Y(n_2149)
);

AOI221xp5_ASAP7_75t_L g2150 ( 
.A1(n_2105),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.C(n_271),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_2107),
.B(n_272),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2102),
.Y(n_2152)
);

O2A1O1Ixp33_ASAP7_75t_L g2153 ( 
.A1(n_2107),
.A2(n_272),
.B(n_273),
.C(n_274),
.Y(n_2153)
);

NAND4xp25_ASAP7_75t_L g2154 ( 
.A(n_2121),
.B(n_273),
.C(n_275),
.D(n_276),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2124),
.Y(n_2155)
);

NAND3xp33_ASAP7_75t_L g2156 ( 
.A(n_2123),
.B(n_275),
.C(n_276),
.Y(n_2156)
);

NOR3xp33_ASAP7_75t_L g2157 ( 
.A(n_2120),
.B(n_277),
.C(n_278),
.Y(n_2157)
);

NAND3xp33_ASAP7_75t_L g2158 ( 
.A(n_2126),
.B(n_277),
.C(n_278),
.Y(n_2158)
);

AOI22xp33_ASAP7_75t_L g2159 ( 
.A1(n_2130),
.A2(n_1946),
.B1(n_1912),
.B2(n_1911),
.Y(n_2159)
);

NOR3x1_ASAP7_75t_L g2160 ( 
.A(n_2138),
.B(n_279),
.C(n_280),
.Y(n_2160)
);

NOR3xp33_ASAP7_75t_L g2161 ( 
.A(n_2137),
.B(n_279),
.C(n_280),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2149),
.B(n_281),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2151),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2153),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2127),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2136),
.Y(n_2166)
);

NOR3xp33_ASAP7_75t_L g2167 ( 
.A(n_2142),
.B(n_282),
.C(n_283),
.Y(n_2167)
);

NOR2x1_ASAP7_75t_L g2168 ( 
.A(n_2139),
.B(n_282),
.Y(n_2168)
);

NOR2x1_ASAP7_75t_L g2169 ( 
.A(n_2122),
.B(n_283),
.Y(n_2169)
);

NOR2xp67_ASAP7_75t_L g2170 ( 
.A(n_2147),
.B(n_284),
.Y(n_2170)
);

NAND4xp75_ASAP7_75t_L g2171 ( 
.A(n_2150),
.B(n_284),
.C(n_285),
.D(n_286),
.Y(n_2171)
);

INVx2_ASAP7_75t_SL g2172 ( 
.A(n_2133),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2148),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_2152),
.B(n_285),
.Y(n_2174)
);

NOR2x1_ASAP7_75t_L g2175 ( 
.A(n_2145),
.B(n_286),
.Y(n_2175)
);

NAND4xp75_ASAP7_75t_L g2176 ( 
.A(n_2131),
.B(n_287),
.C(n_288),
.D(n_289),
.Y(n_2176)
);

NOR3x1_ASAP7_75t_L g2177 ( 
.A(n_2129),
.B(n_288),
.C(n_289),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2134),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2135),
.Y(n_2179)
);

NAND4xp75_ASAP7_75t_L g2180 ( 
.A(n_2146),
.B(n_290),
.C(n_291),
.D(n_292),
.Y(n_2180)
);

INVxp67_ASAP7_75t_L g2181 ( 
.A(n_2128),
.Y(n_2181)
);

A2O1A1Ixp33_ASAP7_75t_L g2182 ( 
.A1(n_2155),
.A2(n_2140),
.B(n_2132),
.C(n_2141),
.Y(n_2182)
);

OR2x2_ASAP7_75t_L g2183 ( 
.A(n_2154),
.B(n_2144),
.Y(n_2183)
);

NOR3xp33_ASAP7_75t_L g2184 ( 
.A(n_2157),
.B(n_2143),
.C(n_2125),
.Y(n_2184)
);

NOR3xp33_ASAP7_75t_SL g2185 ( 
.A(n_2158),
.B(n_290),
.C(n_292),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2156),
.Y(n_2186)
);

INVx2_ASAP7_75t_SL g2187 ( 
.A(n_2172),
.Y(n_2187)
);

AO22x2_ASAP7_75t_L g2188 ( 
.A1(n_2178),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_2188)
);

AND2x4_ASAP7_75t_L g2189 ( 
.A(n_2166),
.B(n_294),
.Y(n_2189)
);

AND2x2_ASAP7_75t_SL g2190 ( 
.A(n_2177),
.B(n_296),
.Y(n_2190)
);

NOR2x1_ASAP7_75t_L g2191 ( 
.A(n_2180),
.B(n_296),
.Y(n_2191)
);

OR2x2_ASAP7_75t_L g2192 ( 
.A(n_2162),
.B(n_297),
.Y(n_2192)
);

AND3x1_ASAP7_75t_L g2193 ( 
.A(n_2161),
.B(n_298),
.C(n_299),
.Y(n_2193)
);

NOR4xp75_ASAP7_75t_L g2194 ( 
.A(n_2176),
.B(n_298),
.C(n_299),
.D(n_300),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2174),
.B(n_300),
.Y(n_2195)
);

HB1xp67_ASAP7_75t_L g2196 ( 
.A(n_2168),
.Y(n_2196)
);

NOR3xp33_ASAP7_75t_L g2197 ( 
.A(n_2164),
.B(n_301),
.C(n_302),
.Y(n_2197)
);

NOR3xp33_ASAP7_75t_L g2198 ( 
.A(n_2181),
.B(n_301),
.C(n_303),
.Y(n_2198)
);

NAND3xp33_ASAP7_75t_L g2199 ( 
.A(n_2167),
.B(n_303),
.C(n_304),
.Y(n_2199)
);

NOR3xp33_ASAP7_75t_L g2200 ( 
.A(n_2173),
.B(n_304),
.C(n_305),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2160),
.B(n_306),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2171),
.Y(n_2202)
);

NAND3x1_ASAP7_75t_L g2203 ( 
.A(n_2169),
.B(n_307),
.C(n_308),
.Y(n_2203)
);

NAND3x1_ASAP7_75t_L g2204 ( 
.A(n_2175),
.B(n_307),
.C(n_308),
.Y(n_2204)
);

NAND2x1p5_ASAP7_75t_L g2205 ( 
.A(n_2163),
.B(n_1899),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_2179),
.B(n_310),
.Y(n_2206)
);

OAI21xp33_ASAP7_75t_SL g2207 ( 
.A1(n_2170),
.A2(n_310),
.B(n_311),
.Y(n_2207)
);

AND3x4_ASAP7_75t_L g2208 ( 
.A(n_2165),
.B(n_311),
.C(n_312),
.Y(n_2208)
);

NOR2x1_ASAP7_75t_L g2209 ( 
.A(n_2159),
.B(n_312),
.Y(n_2209)
);

OR2x2_ASAP7_75t_L g2210 ( 
.A(n_2154),
.B(n_313),
.Y(n_2210)
);

NOR2xp33_ASAP7_75t_L g2211 ( 
.A(n_2154),
.B(n_313),
.Y(n_2211)
);

NAND4xp75_ASAP7_75t_L g2212 ( 
.A(n_2177),
.B(n_314),
.C(n_316),
.D(n_317),
.Y(n_2212)
);

OAI22xp5_ASAP7_75t_L g2213 ( 
.A1(n_2156),
.A2(n_1889),
.B1(n_1899),
.B2(n_1910),
.Y(n_2213)
);

AND3x4_ASAP7_75t_L g2214 ( 
.A(n_2168),
.B(n_314),
.C(n_316),
.Y(n_2214)
);

OA21x2_ASAP7_75t_L g2215 ( 
.A1(n_2178),
.A2(n_317),
.B(n_318),
.Y(n_2215)
);

NOR3xp33_ASAP7_75t_L g2216 ( 
.A(n_2155),
.B(n_318),
.C(n_319),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_2154),
.B(n_320),
.Y(n_2217)
);

AOI221xp5_ASAP7_75t_SL g2218 ( 
.A1(n_2182),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.C(n_323),
.Y(n_2218)
);

AOI21xp5_ASAP7_75t_L g2219 ( 
.A1(n_2187),
.A2(n_323),
.B(n_324),
.Y(n_2219)
);

NOR3xp33_ASAP7_75t_L g2220 ( 
.A(n_2186),
.B(n_325),
.C(n_326),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2215),
.Y(n_2221)
);

XNOR2xp5_ASAP7_75t_L g2222 ( 
.A(n_2214),
.B(n_325),
.Y(n_2222)
);

HB1xp67_ASAP7_75t_L g2223 ( 
.A(n_2188),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2208),
.Y(n_2224)
);

OR2x2_ASAP7_75t_L g2225 ( 
.A(n_2210),
.B(n_326),
.Y(n_2225)
);

OR2x2_ASAP7_75t_L g2226 ( 
.A(n_2205),
.B(n_2195),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2189),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_2196),
.Y(n_2228)
);

OAI211xp5_ASAP7_75t_L g2229 ( 
.A1(n_2207),
.A2(n_327),
.B(n_328),
.C(n_329),
.Y(n_2229)
);

AOI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_2184),
.A2(n_1885),
.B1(n_1936),
.B2(n_1942),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2201),
.Y(n_2231)
);

NAND4xp25_ASAP7_75t_L g2232 ( 
.A(n_2191),
.B(n_328),
.C(n_329),
.D(n_330),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_SL g2233 ( 
.A(n_2190),
.B(n_331),
.Y(n_2233)
);

NAND2xp33_ASAP7_75t_SL g2234 ( 
.A(n_2185),
.B(n_332),
.Y(n_2234)
);

AOI21xp5_ASAP7_75t_L g2235 ( 
.A1(n_2211),
.A2(n_332),
.B(n_333),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2206),
.B(n_334),
.Y(n_2236)
);

AND2x4_ASAP7_75t_L g2237 ( 
.A(n_2194),
.B(n_334),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2217),
.B(n_336),
.Y(n_2238)
);

AND2x4_ASAP7_75t_L g2239 ( 
.A(n_2202),
.B(n_336),
.Y(n_2239)
);

NAND4xp25_ASAP7_75t_L g2240 ( 
.A(n_2199),
.B(n_337),
.C(n_338),
.D(n_339),
.Y(n_2240)
);

INVx1_ASAP7_75t_SL g2241 ( 
.A(n_2204),
.Y(n_2241)
);

INVx2_ASAP7_75t_SL g2242 ( 
.A(n_2188),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2216),
.B(n_337),
.Y(n_2243)
);

NAND2x1p5_ASAP7_75t_L g2244 ( 
.A(n_2193),
.B(n_338),
.Y(n_2244)
);

AOI21xp33_ASAP7_75t_L g2245 ( 
.A1(n_2192),
.A2(n_339),
.B(n_342),
.Y(n_2245)
);

NAND3xp33_ASAP7_75t_SL g2246 ( 
.A(n_2197),
.B(n_2198),
.C(n_2200),
.Y(n_2246)
);

NAND2xp33_ASAP7_75t_SL g2247 ( 
.A(n_2237),
.B(n_2183),
.Y(n_2247)
);

NOR2xp33_ASAP7_75t_R g2248 ( 
.A(n_2234),
.B(n_2203),
.Y(n_2248)
);

NOR3xp33_ASAP7_75t_SL g2249 ( 
.A(n_2228),
.B(n_2212),
.C(n_2209),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_R g2250 ( 
.A(n_2222),
.B(n_342),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_R g2251 ( 
.A(n_2221),
.B(n_343),
.Y(n_2251)
);

XNOR2x1_ASAP7_75t_L g2252 ( 
.A(n_2244),
.B(n_2213),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_2237),
.B(n_343),
.Y(n_2253)
);

NAND2xp33_ASAP7_75t_SL g2254 ( 
.A(n_2223),
.B(n_2242),
.Y(n_2254)
);

NAND2xp33_ASAP7_75t_SL g2255 ( 
.A(n_2233),
.B(n_2236),
.Y(n_2255)
);

NOR2xp33_ASAP7_75t_R g2256 ( 
.A(n_2246),
.B(n_344),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2239),
.B(n_344),
.Y(n_2257)
);

NOR2xp33_ASAP7_75t_R g2258 ( 
.A(n_2224),
.B(n_345),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2219),
.B(n_345),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2220),
.B(n_346),
.Y(n_2260)
);

NAND2xp33_ASAP7_75t_SL g2261 ( 
.A(n_2225),
.B(n_346),
.Y(n_2261)
);

NOR2xp33_ASAP7_75t_R g2262 ( 
.A(n_2227),
.B(n_348),
.Y(n_2262)
);

NOR2xp33_ASAP7_75t_R g2263 ( 
.A(n_2231),
.B(n_348),
.Y(n_2263)
);

NOR2xp33_ASAP7_75t_R g2264 ( 
.A(n_2241),
.B(n_2238),
.Y(n_2264)
);

NOR2xp33_ASAP7_75t_R g2265 ( 
.A(n_2243),
.B(n_349),
.Y(n_2265)
);

XNOR2xp5_ASAP7_75t_L g2266 ( 
.A(n_2232),
.B(n_350),
.Y(n_2266)
);

NAND2xp33_ASAP7_75t_SL g2267 ( 
.A(n_2226),
.B(n_351),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_R g2268 ( 
.A(n_2218),
.B(n_351),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2229),
.B(n_2235),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_R g2270 ( 
.A(n_2245),
.B(n_352),
.Y(n_2270)
);

NOR2xp33_ASAP7_75t_R g2271 ( 
.A(n_2240),
.B(n_352),
.Y(n_2271)
);

NAND2xp33_ASAP7_75t_SL g2272 ( 
.A(n_2230),
.B(n_353),
.Y(n_2272)
);

XNOR2xp5_ASAP7_75t_L g2273 ( 
.A(n_2222),
.B(n_353),
.Y(n_2273)
);

NAND3xp33_ASAP7_75t_SL g2274 ( 
.A(n_2241),
.B(n_354),
.C(n_355),
.Y(n_2274)
);

NAND2xp33_ASAP7_75t_SL g2275 ( 
.A(n_2237),
.B(n_354),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2239),
.B(n_355),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2252),
.Y(n_2277)
);

HB1xp67_ASAP7_75t_L g2278 ( 
.A(n_2262),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2273),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2257),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2276),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2266),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2253),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2259),
.Y(n_2284)
);

CKINVDCx20_ASAP7_75t_R g2285 ( 
.A(n_2247),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2274),
.Y(n_2286)
);

INVx1_ASAP7_75t_SL g2287 ( 
.A(n_2263),
.Y(n_2287)
);

AND2x4_ASAP7_75t_L g2288 ( 
.A(n_2249),
.B(n_357),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2260),
.Y(n_2289)
);

BUFx2_ASAP7_75t_L g2290 ( 
.A(n_2251),
.Y(n_2290)
);

HB1xp67_ASAP7_75t_L g2291 ( 
.A(n_2258),
.Y(n_2291)
);

AOI22x1_ASAP7_75t_L g2292 ( 
.A1(n_2267),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2275),
.Y(n_2293)
);

HB1xp67_ASAP7_75t_L g2294 ( 
.A(n_2248),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2269),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2292),
.Y(n_2296)
);

HB1xp67_ASAP7_75t_L g2297 ( 
.A(n_2288),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2288),
.Y(n_2298)
);

AOI22xp5_ASAP7_75t_L g2299 ( 
.A1(n_2285),
.A2(n_2254),
.B1(n_2255),
.B2(n_2261),
.Y(n_2299)
);

AO22x1_ASAP7_75t_L g2300 ( 
.A1(n_2286),
.A2(n_2256),
.B1(n_2250),
.B2(n_2265),
.Y(n_2300)
);

AOI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_2277),
.A2(n_2272),
.B1(n_2271),
.B2(n_2264),
.Y(n_2301)
);

XOR2xp5_ASAP7_75t_L g2302 ( 
.A(n_2294),
.B(n_2270),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2290),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2278),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2293),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2284),
.Y(n_2306)
);

OAI22xp5_ASAP7_75t_SL g2307 ( 
.A1(n_2287),
.A2(n_2268),
.B1(n_360),
.B2(n_361),
.Y(n_2307)
);

AO21x2_ASAP7_75t_L g2308 ( 
.A1(n_2299),
.A2(n_2279),
.B(n_2282),
.Y(n_2308)
);

OR2x2_ASAP7_75t_L g2309 ( 
.A(n_2298),
.B(n_2291),
.Y(n_2309)
);

AO22x2_ASAP7_75t_L g2310 ( 
.A1(n_2296),
.A2(n_2283),
.B1(n_2281),
.B2(n_2280),
.Y(n_2310)
);

HB1xp67_ASAP7_75t_L g2311 ( 
.A(n_2307),
.Y(n_2311)
);

INVx3_ASAP7_75t_L g2312 ( 
.A(n_2305),
.Y(n_2312)
);

AND3x2_ASAP7_75t_L g2313 ( 
.A(n_2297),
.B(n_2295),
.C(n_2289),
.Y(n_2313)
);

OAI22x1_ASAP7_75t_L g2314 ( 
.A1(n_2301),
.A2(n_359),
.B1(n_360),
.B2(n_361),
.Y(n_2314)
);

HB1xp67_ASAP7_75t_L g2315 ( 
.A(n_2302),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2300),
.Y(n_2316)
);

AOI21xp5_ASAP7_75t_L g2317 ( 
.A1(n_2310),
.A2(n_2304),
.B(n_2303),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2312),
.Y(n_2318)
);

NAND5xp2_ASAP7_75t_L g2319 ( 
.A(n_2316),
.B(n_2306),
.C(n_363),
.D(n_364),
.E(n_365),
.Y(n_2319)
);

O2A1O1Ixp33_ASAP7_75t_SL g2320 ( 
.A1(n_2311),
.A2(n_362),
.B(n_363),
.C(n_364),
.Y(n_2320)
);

AOI22xp5_ASAP7_75t_L g2321 ( 
.A1(n_2318),
.A2(n_2308),
.B1(n_2315),
.B2(n_2309),
.Y(n_2321)
);

HB1xp67_ASAP7_75t_L g2322 ( 
.A(n_2317),
.Y(n_2322)
);

OAI22xp5_ASAP7_75t_SL g2323 ( 
.A1(n_2319),
.A2(n_2314),
.B1(n_2313),
.B2(n_369),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2320),
.Y(n_2324)
);

OAI331xp33_ASAP7_75t_L g2325 ( 
.A1(n_2322),
.A2(n_362),
.A3(n_368),
.B1(n_369),
.B2(n_370),
.B3(n_371),
.C1(n_372),
.Y(n_2325)
);

AOI21xp5_ASAP7_75t_L g2326 ( 
.A1(n_2323),
.A2(n_2324),
.B(n_2321),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2322),
.B(n_368),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2327),
.B(n_370),
.Y(n_2328)
);

OAI211xp5_ASAP7_75t_L g2329 ( 
.A1(n_2326),
.A2(n_371),
.B(n_373),
.C(n_374),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2328),
.B(n_2325),
.Y(n_2330)
);

OAI21xp5_ASAP7_75t_L g2331 ( 
.A1(n_2329),
.A2(n_374),
.B(n_375),
.Y(n_2331)
);

O2A1O1Ixp33_ASAP7_75t_L g2332 ( 
.A1(n_2330),
.A2(n_375),
.B(n_377),
.C(n_378),
.Y(n_2332)
);

AOI22xp33_ASAP7_75t_SL g2333 ( 
.A1(n_2332),
.A2(n_2331),
.B1(n_378),
.B2(n_379),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2333),
.B(n_377),
.Y(n_2334)
);

AOI221xp5_ASAP7_75t_L g2335 ( 
.A1(n_2334),
.A2(n_379),
.B1(n_380),
.B2(n_381),
.C(n_382),
.Y(n_2335)
);

AOI211xp5_ASAP7_75t_L g2336 ( 
.A1(n_2335),
.A2(n_380),
.B(n_382),
.C(n_383),
.Y(n_2336)
);


endmodule