module real_jpeg_11364_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_309, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_309;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_3),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_3),
.A2(n_27),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_3),
.B(n_176),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_L g245 ( 
.A1(n_3),
.A2(n_51),
.B1(n_52),
.B2(n_184),
.Y(n_245)
);

O2A1O1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_3),
.A2(n_52),
.B(n_63),
.C(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_3),
.B(n_56),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_3),
.B(n_84),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_3),
.B(n_58),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_3),
.A2(n_36),
.B(n_46),
.C(n_282),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_4),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_4),
.A2(n_33),
.B1(n_36),
.B2(n_133),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_4),
.A2(n_51),
.B1(n_52),
.B2(n_133),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_4),
.A2(n_60),
.B1(n_64),
.B2(n_133),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_6),
.A2(n_33),
.B1(n_36),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_6),
.A2(n_45),
.B1(n_51),
.B2(n_52),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_45),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_6),
.A2(n_45),
.B1(n_60),
.B2(n_64),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_7),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_7),
.A2(n_33),
.B1(n_36),
.B2(n_157),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_7),
.A2(n_51),
.B1(n_52),
.B2(n_157),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_7),
.A2(n_60),
.B1(n_64),
.B2(n_157),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_8),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_8),
.A2(n_33),
.B1(n_36),
.B2(n_91),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_8),
.A2(n_51),
.B1(n_52),
.B2(n_91),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_8),
.A2(n_60),
.B1(n_64),
.B2(n_91),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_12),
.A2(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_12),
.A2(n_30),
.B1(n_51),
.B2(n_52),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_12),
.A2(n_30),
.B1(n_60),
.B2(n_64),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_13),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_13),
.A2(n_33),
.B1(n_36),
.B2(n_173),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_13),
.A2(n_51),
.B1(n_52),
.B2(n_173),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_13),
.A2(n_60),
.B1(n_64),
.B2(n_173),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_14),
.A2(n_33),
.B1(n_36),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_14),
.A2(n_51),
.B1(n_52),
.B2(n_55),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_14),
.A2(n_55),
.B1(n_60),
.B2(n_64),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_15),
.A2(n_51),
.B1(n_52),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_15),
.A2(n_60),
.B1(n_64),
.B2(n_68),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_15),
.A2(n_33),
.B1(n_36),
.B2(n_68),
.Y(n_101)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_17),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_17),
.A2(n_33),
.B1(n_36),
.B2(n_39),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_17),
.A2(n_39),
.B1(n_51),
.B2(n_52),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_17),
.A2(n_39),
.B1(n_60),
.B2(n_64),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_105),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_92),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_22),
.B(n_92),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_70),
.C(n_77),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_23),
.A2(n_70),
.B1(n_71),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_24),
.A2(n_25),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_25),
.B(n_43),
.C(n_57),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_27),
.A2(n_33),
.A3(n_35),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_28),
.B(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_31),
.A2(n_32),
.B1(n_38),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_31),
.A2(n_32),
.B1(n_90),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_31),
.A2(n_32),
.B1(n_132),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_31),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_31),
.A2(n_32),
.B1(n_172),
.B2(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_37),
.Y(n_31)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_32),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_33),
.B(n_184),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_34),
.B(n_36),
.Y(n_182)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_36),
.A2(n_48),
.A3(n_51),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_57),
.B2(n_69),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_53),
.B2(n_56),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_46),
.B1(n_56),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_46),
.A2(n_56),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_46),
.A2(n_56),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_49),
.B(n_52),
.Y(n_225)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_50),
.A2(n_54),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_50),
.A2(n_74),
.B1(n_100),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_50),
.A2(n_100),
.B1(n_130),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_50),
.A2(n_100),
.B1(n_168),
.B2(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_50),
.A2(n_211),
.B(n_281),
.Y(n_280)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_52),
.B1(n_62),
.B2(n_63),
.Y(n_66)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_57),
.A2(n_69),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_65),
.B(n_67),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_65),
.B1(n_67),
.B2(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_65),
.B1(n_76),
.B2(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_58),
.A2(n_65),
.B1(n_88),
.B2(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_58),
.A2(n_65),
.B1(n_151),
.B2(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_58),
.A2(n_65),
.B1(n_189),
.B2(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_58),
.A2(n_65),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_58),
.A2(n_65),
.B1(n_246),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_59),
.A2(n_128),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_59),
.A2(n_152),
.B1(n_219),
.B2(n_284),
.Y(n_283)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_60),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_60),
.B(n_269),
.Y(n_268)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_62),
.A2(n_64),
.B(n_184),
.Y(n_248)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_65),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_72),
.B(n_75),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B(n_89),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_78),
.A2(n_79),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_86),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_81),
.B1(n_89),
.B2(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_80),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_141)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_84),
.B(n_85),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_82),
.A2(n_84),
.B1(n_85),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_82),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_82),
.A2(n_84),
.B1(n_148),
.B2(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_82),
.A2(n_84),
.B1(n_180),
.B2(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_82),
.A2(n_84),
.B1(n_216),
.B2(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_82),
.A2(n_84),
.B1(n_227),
.B2(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_82),
.A2(n_84),
.B1(n_184),
.B2(n_267),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_82),
.A2(n_84),
.B1(n_260),
.B2(n_267),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_83),
.A2(n_124),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_83),
.A2(n_146),
.B1(n_259),
.B2(n_261),
.Y(n_258)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_89),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_102),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_134),
.B(n_307),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_107),
.B(n_110),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.C(n_118),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_129),
.C(n_131),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_120),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_126),
.Y(n_197)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_131),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_160),
.B(n_306),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_158),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_137),
.B(n_158),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_142),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_138),
.B(n_141),
.Y(n_304)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_142),
.B(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_153),
.C(n_155),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_143),
.A2(n_144),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_149),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_155),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_301),
.B(n_305),
.Y(n_160)
);

OAI221xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_204),
.B1(n_299),
.B2(n_300),
.C(n_309),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_195),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_163),
.B(n_195),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_185),
.C(n_186),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_164),
.B(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_177),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_170),
.C(n_177),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_183),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_185),
.B(n_186),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_203),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_197),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_197),
.B(n_202),
.C(n_203),
.Y(n_302)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_295),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_238),
.B(n_294),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_228),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_207),
.B(n_228),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_217),
.C(n_220),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_208),
.B(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_214),
.C(n_215),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_217),
.A2(n_220),
.B1(n_221),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_217),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_224),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_226),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_233),
.B2(n_237),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_229),
.B(n_234),
.C(n_236),
.Y(n_296)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_233),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_288),
.B(n_293),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_276),
.B(n_287),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_256),
.B(n_275),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_249),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_242),
.B(n_249),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_243),
.A2(n_244),
.B1(n_247),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_252),
.C(n_254),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_255),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_264),
.B(n_274),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_262),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_258),
.B(n_262),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_270),
.B(n_273),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_271),
.B(n_272),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_277),
.B(n_278),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_285),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_283),
.C(n_285),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_289),
.B(n_290),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_297),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.Y(n_305)
);


endmodule