module fake_jpeg_23821_n_321 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_6),
.B(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_45),
.Y(n_66)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_48),
.Y(n_53)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_9),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_30),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_24),
.B1(n_18),
.B2(n_34),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_50),
.A2(n_68),
.B1(n_76),
.B2(n_82),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_32),
.C(n_31),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_29),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_56),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_55),
.B(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_20),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_25),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_31),
.B1(n_32),
.B2(n_25),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_60),
.A2(n_61),
.B1(n_71),
.B2(n_79),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_24),
.B1(n_35),
.B2(n_18),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_81),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_31),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_25),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_35),
.B1(n_18),
.B2(n_32),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_30),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_38),
.B1(n_37),
.B2(n_33),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_70),
.A2(n_78),
.B1(n_1),
.B2(n_2),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_40),
.A2(n_30),
.B1(n_33),
.B2(n_37),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_40),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_72),
.Y(n_110)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_42),
.B(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_40),
.A2(n_26),
.B1(n_23),
.B2(n_19),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_26),
.Y(n_77)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_40),
.A2(n_28),
.B1(n_27),
.B2(n_22),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_41),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_28),
.B1(n_27),
.B2(n_25),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_25),
.B1(n_0),
.B2(n_2),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_85),
.B1(n_67),
.B2(n_66),
.Y(n_101)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_89),
.Y(n_127)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_93),
.A2(n_62),
.B(n_60),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_25),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_98),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_0),
.Y(n_98)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_104),
.B1(n_99),
.B2(n_89),
.Y(n_140)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_102),
.B(n_108),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_52),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_111),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_1),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_112),
.Y(n_123)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_109),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_1),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_3),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_55),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_113),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_72),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_4),
.Y(n_118)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_53),
.B(n_4),
.Y(n_119)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_126),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_69),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_125),
.B(n_143),
.C(n_8),
.Y(n_188)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_54),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_142),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_67),
.B1(n_80),
.B2(n_63),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_135),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_134),
.Y(n_172)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_94),
.A2(n_61),
.B1(n_71),
.B2(n_58),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_140),
.B1(n_103),
.B2(n_111),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_86),
.A2(n_79),
.B1(n_84),
.B2(n_60),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_145),
.B1(n_101),
.B2(n_107),
.Y(n_166)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_148),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_60),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_53),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_144),
.B(n_91),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_86),
.A2(n_80),
.B1(n_5),
.B2(n_6),
.Y(n_145)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_153),
.Y(n_187)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_4),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_5),
.C(n_8),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_155),
.B(n_160),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_139),
.B(n_91),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_159),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_152),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_103),
.B1(n_109),
.B2(n_88),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_166),
.B1(n_171),
.B2(n_186),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_117),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_162),
.A2(n_167),
.B(n_8),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_139),
.B(n_105),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_98),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_165),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_88),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_117),
.B(n_88),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_130),
.B(n_95),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_170),
.Y(n_196)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_169),
.B(n_181),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_107),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_120),
.B1(n_116),
.B2(n_96),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_96),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_178),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_137),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_115),
.Y(n_179)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_123),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_183),
.Y(n_191)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_115),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_129),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_97),
.Y(n_185)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_116),
.B1(n_9),
.B2(n_11),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_188),
.A2(n_165),
.B(n_155),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_177),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_192),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_179),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_193),
.B(n_198),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_132),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_204),
.C(n_213),
.Y(n_224)
);

OA21x2_ASAP7_75t_L g197 ( 
.A1(n_162),
.A2(n_133),
.B(n_153),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_197),
.A2(n_209),
.B(n_212),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_173),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_201),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_132),
.B(n_147),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_202),
.A2(n_216),
.B(n_180),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_176),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_206),
.B(n_207),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_175),
.A2(n_129),
.B(n_126),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_211),
.Y(n_223)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_135),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_218),
.Y(n_225)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_205),
.A2(n_200),
.B1(n_161),
.B2(n_156),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_227),
.B1(n_236),
.B2(n_240),
.Y(n_246)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_221),
.B(n_241),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_204),
.B(n_162),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_237),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_197),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_232),
.B1(n_238),
.B2(n_209),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_200),
.A2(n_181),
.B1(n_172),
.B2(n_158),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_167),
.C(n_168),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_229),
.C(n_235),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_157),
.C(n_164),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_241),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_171),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_199),
.A2(n_166),
.B1(n_160),
.B2(n_159),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_169),
.C(n_186),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_122),
.B(n_149),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_199),
.A2(n_215),
.B1(n_197),
.B2(n_190),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_149),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_214),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_197),
.Y(n_243)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_244),
.A2(n_239),
.B1(n_234),
.B2(n_210),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_255),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_235),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_196),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_239),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_196),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_228),
.C(n_229),
.Y(n_267)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_240),
.B(n_212),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_259),
.B(n_236),
.Y(n_276)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_260),
.B(n_261),
.Y(n_264)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_226),
.B(n_191),
.C(n_189),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_262),
.A2(n_278),
.B1(n_263),
.B2(n_274),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_265),
.A2(n_277),
.B(n_203),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_270),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_220),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_217),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_237),
.C(n_189),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_257),
.C(n_247),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_226),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_274),
.B(n_198),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_276),
.B(n_259),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_253),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_246),
.A2(n_190),
.B1(n_231),
.B2(n_218),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_282),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_232),
.B(n_238),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_288),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_245),
.C(n_251),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_284),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_245),
.C(n_254),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_285),
.A2(n_286),
.B1(n_275),
.B2(n_271),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_262),
.A2(n_203),
.B1(n_211),
.B2(n_192),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_287),
.A2(n_288),
.B(n_206),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_270),
.B(n_212),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_249),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g295 ( 
.A(n_290),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_267),
.C(n_264),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_272),
.Y(n_294)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_292),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_296),
.C(n_281),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_268),
.B1(n_266),
.B2(n_278),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_282),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_291),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_11),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_146),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_302),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_304),
.B(n_305),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_283),
.B(n_284),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_306),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_308),
.B1(n_148),
.B2(n_12),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_146),
.Y(n_308)
);

NOR3xp33_ASAP7_75t_SL g312 ( 
.A(n_302),
.B(n_295),
.C(n_12),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_313),
.Y(n_314)
);

AOI31xp67_ASAP7_75t_SL g315 ( 
.A1(n_311),
.A2(n_301),
.A3(n_303),
.B(n_14),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_315),
.A2(n_314),
.B1(n_13),
.B2(n_15),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_309),
.A2(n_310),
.B(n_13),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_11),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_318),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_319),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_16),
.Y(n_321)
);


endmodule